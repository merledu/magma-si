module fancontrol(
  input        clock,
  input        reset,
  output       io_o_reduction_add_0,
  output       io_o_reduction_add_1,
  output       io_o_reduction_add_2,
  output       io_o_reduction_add_3,
  output       io_o_reduction_add_4,
  output       io_o_reduction_add_5,
  output       io_o_reduction_add_6,
  output       io_o_reduction_add_7,
  output       io_o_reduction_add_8,
  output       io_o_reduction_add_9,
  output       io_o_reduction_add_10,
  output       io_o_reduction_add_11,
  output       io_o_reduction_add_12,
  output       io_o_reduction_add_13,
  output       io_o_reduction_add_14,
  output       io_o_reduction_add_15,
  output       io_o_reduction_add_16,
  output       io_o_reduction_add_17,
  output       io_o_reduction_add_18,
  output       io_o_reduction_add_19,
  output       io_o_reduction_add_20,
  output       io_o_reduction_add_21,
  output       io_o_reduction_add_22,
  output       io_o_reduction_add_23,
  output       io_o_reduction_add_24,
  output       io_o_reduction_add_25,
  output       io_o_reduction_add_26,
  output       io_o_reduction_add_27,
  output       io_o_reduction_add_28,
  output       io_o_reduction_add_29,
  output       io_o_reduction_add_30,
  output [2:0] io_o_reduction_cmd_0,
  output [2:0] io_o_reduction_cmd_1,
  output [2:0] io_o_reduction_cmd_2,
  output [2:0] io_o_reduction_cmd_3,
  output [2:0] io_o_reduction_cmd_4,
  output [2:0] io_o_reduction_cmd_5,
  output [2:0] io_o_reduction_cmd_6,
  output [2:0] io_o_reduction_cmd_7,
  output [2:0] io_o_reduction_cmd_8,
  output [2:0] io_o_reduction_cmd_9,
  output [2:0] io_o_reduction_cmd_10,
  output [2:0] io_o_reduction_cmd_11,
  output [2:0] io_o_reduction_cmd_12,
  output [2:0] io_o_reduction_cmd_13,
  output [2:0] io_o_reduction_cmd_14,
  output [2:0] io_o_reduction_cmd_15,
  output [2:0] io_o_reduction_cmd_16,
  output [2:0] io_o_reduction_cmd_17,
  output [2:0] io_o_reduction_cmd_18,
  output [2:0] io_o_reduction_cmd_19,
  output [2:0] io_o_reduction_cmd_20,
  output [2:0] io_o_reduction_cmd_21,
  output [2:0] io_o_reduction_cmd_22,
  output [2:0] io_o_reduction_cmd_23,
  output [2:0] io_o_reduction_cmd_24,
  output [2:0] io_o_reduction_cmd_25,
  output [2:0] io_o_reduction_cmd_26,
  output [2:0] io_o_reduction_cmd_27,
  output [2:0] io_o_reduction_cmd_28,
  output [2:0] io_o_reduction_cmd_29,
  output [2:0] io_o_reduction_cmd_30,
  output [1:0] io_o_reduction_sel_0,
  output [1:0] io_o_reduction_sel_1,
  output [1:0] io_o_reduction_sel_2,
  output [1:0] io_o_reduction_sel_3,
  output [1:0] io_o_reduction_sel_4,
  output [1:0] io_o_reduction_sel_5,
  output [1:0] io_o_reduction_sel_6,
  output [1:0] io_o_reduction_sel_7,
  output [1:0] io_o_reduction_sel_8,
  output [1:0] io_o_reduction_sel_9,
  output [1:0] io_o_reduction_sel_10,
  output [1:0] io_o_reduction_sel_11,
  output [1:0] io_o_reduction_sel_12,
  output [1:0] io_o_reduction_sel_13,
  output [1:0] io_o_reduction_sel_14,
  output [1:0] io_o_reduction_sel_15,
  output [1:0] io_o_reduction_sel_16,
  output [1:0] io_o_reduction_sel_17,
  output [1:0] io_o_reduction_sel_18,
  output [1:0] io_o_reduction_sel_19,
  output       io_o_reduction_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
`endif // RANDOMIZE_REG_INIT
  reg  r_reduction_add_0; // @[FanCtrl.scala 19:34]
  reg  r_reduction_add_1; // @[FanCtrl.scala 19:34]
  reg  r_reduction_add_2; // @[FanCtrl.scala 19:34]
  reg  r_reduction_add_3; // @[FanCtrl.scala 19:34]
  reg  r_reduction_add_4; // @[FanCtrl.scala 19:34]
  reg  r_reduction_add_5; // @[FanCtrl.scala 19:34]
  reg  r_reduction_add_6; // @[FanCtrl.scala 19:34]
  reg  r_reduction_add_7; // @[FanCtrl.scala 19:34]
  reg  r_reduction_add_8; // @[FanCtrl.scala 19:34]
  reg  r_reduction_add_9; // @[FanCtrl.scala 19:34]
  reg  r_reduction_add_10; // @[FanCtrl.scala 19:34]
  reg  r_reduction_add_11; // @[FanCtrl.scala 19:34]
  reg  r_reduction_add_12; // @[FanCtrl.scala 19:34]
  reg  r_reduction_add_13; // @[FanCtrl.scala 19:34]
  reg  r_reduction_add_14; // @[FanCtrl.scala 19:34]
  reg  r_reduction_add_15; // @[FanCtrl.scala 19:34]
  reg  r_reduction_add_16; // @[FanCtrl.scala 19:34]
  reg  r_reduction_add_17; // @[FanCtrl.scala 19:34]
  reg  r_reduction_add_18; // @[FanCtrl.scala 19:34]
  reg  r_reduction_add_19; // @[FanCtrl.scala 19:34]
  reg  r_reduction_add_20; // @[FanCtrl.scala 19:34]
  reg  r_reduction_add_21; // @[FanCtrl.scala 19:34]
  reg  r_reduction_add_22; // @[FanCtrl.scala 19:34]
  reg  r_reduction_add_23; // @[FanCtrl.scala 19:34]
  reg  r_reduction_add_24; // @[FanCtrl.scala 19:34]
  reg  r_reduction_add_25; // @[FanCtrl.scala 19:34]
  reg  r_reduction_add_26; // @[FanCtrl.scala 19:34]
  reg  r_reduction_add_27; // @[FanCtrl.scala 19:34]
  reg  r_reduction_add_28; // @[FanCtrl.scala 19:34]
  reg  r_reduction_add_29; // @[FanCtrl.scala 19:34]
  reg  r_reduction_add_30; // @[FanCtrl.scala 19:34]
  reg [2:0] r_reduction_cmd_0; // @[FanCtrl.scala 20:34]
  reg [2:0] r_reduction_cmd_1; // @[FanCtrl.scala 20:34]
  reg [2:0] r_reduction_cmd_2; // @[FanCtrl.scala 20:34]
  reg [2:0] r_reduction_cmd_3; // @[FanCtrl.scala 20:34]
  reg [2:0] r_reduction_cmd_4; // @[FanCtrl.scala 20:34]
  reg [2:0] r_reduction_cmd_5; // @[FanCtrl.scala 20:34]
  reg [2:0] r_reduction_cmd_6; // @[FanCtrl.scala 20:34]
  reg [2:0] r_reduction_cmd_7; // @[FanCtrl.scala 20:34]
  reg [2:0] r_reduction_cmd_8; // @[FanCtrl.scala 20:34]
  reg [2:0] r_reduction_cmd_9; // @[FanCtrl.scala 20:34]
  reg [2:0] r_reduction_cmd_10; // @[FanCtrl.scala 20:34]
  reg [2:0] r_reduction_cmd_11; // @[FanCtrl.scala 20:34]
  reg [2:0] r_reduction_cmd_12; // @[FanCtrl.scala 20:34]
  reg [2:0] r_reduction_cmd_13; // @[FanCtrl.scala 20:34]
  reg [2:0] r_reduction_cmd_14; // @[FanCtrl.scala 20:34]
  reg [2:0] r_reduction_cmd_15; // @[FanCtrl.scala 20:34]
  reg [2:0] r_reduction_cmd_16; // @[FanCtrl.scala 20:34]
  reg [2:0] r_reduction_cmd_17; // @[FanCtrl.scala 20:34]
  reg [2:0] r_reduction_cmd_18; // @[FanCtrl.scala 20:34]
  reg [2:0] r_reduction_cmd_19; // @[FanCtrl.scala 20:34]
  reg [2:0] r_reduction_cmd_20; // @[FanCtrl.scala 20:34]
  reg [2:0] r_reduction_cmd_21; // @[FanCtrl.scala 20:34]
  reg [2:0] r_reduction_cmd_22; // @[FanCtrl.scala 20:34]
  reg [2:0] r_reduction_cmd_23; // @[FanCtrl.scala 20:34]
  reg [2:0] r_reduction_cmd_24; // @[FanCtrl.scala 20:34]
  reg [2:0] r_reduction_cmd_25; // @[FanCtrl.scala 20:34]
  reg [2:0] r_reduction_cmd_26; // @[FanCtrl.scala 20:34]
  reg [2:0] r_reduction_cmd_27; // @[FanCtrl.scala 20:34]
  reg [2:0] r_reduction_cmd_28; // @[FanCtrl.scala 20:34]
  reg [2:0] r_reduction_cmd_29; // @[FanCtrl.scala 20:34]
  reg [2:0] r_reduction_cmd_30; // @[FanCtrl.scala 20:34]
  reg [1:0] r_reduction_sel_0; // @[FanCtrl.scala 21:34]
  reg [1:0] r_reduction_sel_1; // @[FanCtrl.scala 21:34]
  reg [1:0] r_reduction_sel_2; // @[FanCtrl.scala 21:34]
  reg [1:0] r_reduction_sel_3; // @[FanCtrl.scala 21:34]
  reg [1:0] r_reduction_sel_4; // @[FanCtrl.scala 21:34]
  reg [1:0] r_reduction_sel_5; // @[FanCtrl.scala 21:34]
  reg [1:0] r_reduction_sel_6; // @[FanCtrl.scala 21:34]
  reg [1:0] r_reduction_sel_7; // @[FanCtrl.scala 21:34]
  reg [1:0] r_reduction_sel_8; // @[FanCtrl.scala 21:34]
  reg [1:0] r_reduction_sel_9; // @[FanCtrl.scala 21:34]
  reg [1:0] r_reduction_sel_10; // @[FanCtrl.scala 21:34]
  reg [1:0] r_reduction_sel_11; // @[FanCtrl.scala 21:34]
  reg [1:0] r_reduction_sel_12; // @[FanCtrl.scala 21:34]
  reg [1:0] r_reduction_sel_13; // @[FanCtrl.scala 21:34]
  reg [1:0] r_reduction_sel_14; // @[FanCtrl.scala 21:34]
  reg [1:0] r_reduction_sel_15; // @[FanCtrl.scala 21:34]
  reg [1:0] r_reduction_sel_16; // @[FanCtrl.scala 21:34]
  reg [1:0] r_reduction_sel_17; // @[FanCtrl.scala 21:34]
  reg [1:0] r_reduction_sel_18; // @[FanCtrl.scala 21:34]
  reg [1:0] r_reduction_sel_19; // @[FanCtrl.scala 21:34]
  reg  r_add_lvl_0Reg_0; // @[FanCtrl.scala 23:33]
  reg  r_add_lvl_0Reg_1; // @[FanCtrl.scala 23:33]
  reg  r_add_lvl_0Reg_2; // @[FanCtrl.scala 23:33]
  reg  r_add_lvl_0Reg_3; // @[FanCtrl.scala 23:33]
  reg  r_add_lvl_0Reg_4; // @[FanCtrl.scala 23:33]
  reg  r_add_lvl_0Reg_5; // @[FanCtrl.scala 23:33]
  reg  r_add_lvl_0Reg_6; // @[FanCtrl.scala 23:33]
  reg  r_add_lvl_0Reg_7; // @[FanCtrl.scala 23:33]
  reg  r_add_lvl_0Reg_8; // @[FanCtrl.scala 23:33]
  reg  r_add_lvl_0Reg_9; // @[FanCtrl.scala 23:33]
  reg  r_add_lvl_0Reg_10; // @[FanCtrl.scala 23:33]
  reg  r_add_lvl_0Reg_11; // @[FanCtrl.scala 23:33]
  reg  r_add_lvl_0Reg_12; // @[FanCtrl.scala 23:33]
  reg  r_add_lvl_0Reg_13; // @[FanCtrl.scala 23:33]
  reg  r_add_lvl_0Reg_14; // @[FanCtrl.scala 23:33]
  reg  r_add_lvl_0Reg_15; // @[FanCtrl.scala 23:33]
  reg  r_add_lvl_1Reg_8; // @[FanCtrl.scala 24:33]
  reg  r_add_lvl_1Reg_9; // @[FanCtrl.scala 24:33]
  reg  r_add_lvl_1Reg_10; // @[FanCtrl.scala 24:33]
  reg  r_add_lvl_1Reg_11; // @[FanCtrl.scala 24:33]
  reg  r_add_lvl_1Reg_12; // @[FanCtrl.scala 24:33]
  reg  r_add_lvl_1Reg_13; // @[FanCtrl.scala 24:33]
  reg  r_add_lvl_1Reg_14; // @[FanCtrl.scala 24:33]
  reg  r_add_lvl_1Reg_15; // @[FanCtrl.scala 24:33]
  reg  r_add_lvl_2Reg_8; // @[FanCtrl.scala 25:33]
  reg  r_add_lvl_2Reg_9; // @[FanCtrl.scala 25:33]
  reg  r_add_lvl_2Reg_10; // @[FanCtrl.scala 25:33]
  reg  r_add_lvl_2Reg_11; // @[FanCtrl.scala 25:33]
  reg  r_add_lvl_3Reg_6; // @[FanCtrl.scala 26:33]
  reg  r_add_lvl_3Reg_7; // @[FanCtrl.scala 26:33]
  reg  r_add_lvl_4Reg_4; // @[FanCtrl.scala 27:33]
  reg [2:0] r_cmd_lvl_0Reg_0; // @[FanCtrl.scala 29:33]
  reg [2:0] r_cmd_lvl_0Reg_1; // @[FanCtrl.scala 29:33]
  reg [2:0] r_cmd_lvl_0Reg_2; // @[FanCtrl.scala 29:33]
  reg [2:0] r_cmd_lvl_0Reg_3; // @[FanCtrl.scala 29:33]
  reg [2:0] r_cmd_lvl_0Reg_4; // @[FanCtrl.scala 29:33]
  reg [2:0] r_cmd_lvl_0Reg_5; // @[FanCtrl.scala 29:33]
  reg [2:0] r_cmd_lvl_0Reg_6; // @[FanCtrl.scala 29:33]
  reg [2:0] r_cmd_lvl_0Reg_7; // @[FanCtrl.scala 29:33]
  reg [2:0] r_cmd_lvl_0Reg_8; // @[FanCtrl.scala 29:33]
  reg [2:0] r_cmd_lvl_0Reg_9; // @[FanCtrl.scala 29:33]
  reg [2:0] r_cmd_lvl_0Reg_10; // @[FanCtrl.scala 29:33]
  reg [2:0] r_cmd_lvl_0Reg_11; // @[FanCtrl.scala 29:33]
  reg [2:0] r_cmd_lvl_0Reg_12; // @[FanCtrl.scala 29:33]
  reg [2:0] r_cmd_lvl_0Reg_13; // @[FanCtrl.scala 29:33]
  reg [2:0] r_cmd_lvl_0Reg_14; // @[FanCtrl.scala 29:33]
  reg [2:0] r_cmd_lvl_0Reg_15; // @[FanCtrl.scala 29:33]
  reg [2:0] r_cmd_lvl_1Reg_8; // @[FanCtrl.scala 30:33]
  reg [2:0] r_cmd_lvl_1Reg_9; // @[FanCtrl.scala 30:33]
  reg [2:0] r_cmd_lvl_1Reg_10; // @[FanCtrl.scala 30:33]
  reg [2:0] r_cmd_lvl_1Reg_11; // @[FanCtrl.scala 30:33]
  reg [2:0] r_cmd_lvl_1Reg_12; // @[FanCtrl.scala 30:33]
  reg [2:0] r_cmd_lvl_1Reg_13; // @[FanCtrl.scala 30:33]
  reg [2:0] r_cmd_lvl_1Reg_14; // @[FanCtrl.scala 30:33]
  reg [2:0] r_cmd_lvl_1Reg_15; // @[FanCtrl.scala 30:33]
  reg [2:0] r_cmd_lvl_2Reg_8; // @[FanCtrl.scala 31:33]
  reg [2:0] r_cmd_lvl_2Reg_9; // @[FanCtrl.scala 31:33]
  reg [2:0] r_cmd_lvl_2Reg_10; // @[FanCtrl.scala 31:33]
  reg [2:0] r_cmd_lvl_2Reg_11; // @[FanCtrl.scala 31:33]
  reg [2:0] r_cmd_lvl_3Reg_6; // @[FanCtrl.scala 32:33]
  reg [2:0] r_cmd_lvl_3Reg_7; // @[FanCtrl.scala 32:33]
  reg [2:0] r_cmd_lvl_4Reg_4; // @[FanCtrl.scala 33:33]
  reg [1:0] r_sel_lvl_2Reg_16; // @[FanCtrl.scala 35:33]
  reg [1:0] r_sel_lvl_2Reg_17; // @[FanCtrl.scala 35:33]
  reg [1:0] r_sel_lvl_2Reg_18; // @[FanCtrl.scala 35:33]
  reg [1:0] r_sel_lvl_2Reg_19; // @[FanCtrl.scala 35:33]
  reg [1:0] r_sel_lvl_2Reg_20; // @[FanCtrl.scala 35:33]
  reg [1:0] r_sel_lvl_2Reg_21; // @[FanCtrl.scala 35:33]
  reg [1:0] r_sel_lvl_2Reg_22; // @[FanCtrl.scala 35:33]
  reg [1:0] r_sel_lvl_2Reg_23; // @[FanCtrl.scala 35:33]
  reg [1:0] r_sel_lvl_3Reg_24; // @[FanCtrl.scala 36:33]
  reg [1:0] r_sel_lvl_3Reg_25; // @[FanCtrl.scala 36:33]
  reg [1:0] r_sel_lvl_3Reg_26; // @[FanCtrl.scala 36:33]
  reg [1:0] r_sel_lvl_3Reg_27; // @[FanCtrl.scala 36:33]
  reg [1:0] r_sel_lvl_3Reg_28; // @[FanCtrl.scala 36:33]
  reg [1:0] r_sel_lvl_3Reg_29; // @[FanCtrl.scala 36:33]
  reg [1:0] r_sel_lvl_3Reg_30; // @[FanCtrl.scala 36:33]
  reg [1:0] r_sel_lvl_3Reg_31; // @[FanCtrl.scala 36:33]
  reg [1:0] r_sel_lvl_4Reg_16; // @[FanCtrl.scala 37:33]
  reg [1:0] r_sel_lvl_4Reg_17; // @[FanCtrl.scala 37:33]
  reg [1:0] r_sel_lvl_4Reg_18; // @[FanCtrl.scala 37:33]
  reg [1:0] r_sel_lvl_4Reg_19; // @[FanCtrl.scala 37:33]
  reg [4:0] w_vn_3; // @[FanCtrl.scala 40:23]
  reg [4:0] w_vn_4; // @[FanCtrl.scala 40:23]
  reg [4:0] w_vn_7; // @[FanCtrl.scala 40:23]
  reg [4:0] w_vn_8; // @[FanCtrl.scala 40:23]
  reg [4:0] w_vn_11; // @[FanCtrl.scala 40:23]
  reg [4:0] w_vn_12; // @[FanCtrl.scala 40:23]
  reg [4:0] w_vn_13; // @[FanCtrl.scala 40:23]
  reg [4:0] w_vn_15; // @[FanCtrl.scala 40:23]
  reg [4:0] w_vn_16; // @[FanCtrl.scala 40:23]
  reg [4:0] w_vn_18; // @[FanCtrl.scala 40:23]
  reg [4:0] w_vn_23; // @[FanCtrl.scala 40:23]
  reg [4:0] w_vn_24; // @[FanCtrl.scala 40:23]
  reg  r_valid_0; // @[FanCtrl.scala 41:26]
  reg  r_valid_1; // @[FanCtrl.scala 41:26]
  reg  r_valid_2; // @[FanCtrl.scala 41:26]
  reg  r_valid_3; // @[FanCtrl.scala 41:26]
  wire [2:0] _T_2 = 2'h2 * 1'h0; // @[FanCtrl.scala 48:25]
  wire [3:0] _T_3 = {{1'd0}, _T_2}; // @[FanCtrl.scala 48:31]
  wire [2:0] _T_7 = _T_2 + 3'h1; // @[FanCtrl.scala 48:58]
  wire [4:0] _GEN_3 = 3'h3 == _T_3[2:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_4 = 3'h4 == _T_3[2:0] ? w_vn_4 : _GEN_3; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_5 = 3'h5 == _T_3[2:0] ? 5'h0 : _GEN_4; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_6 = 3'h6 == _T_3[2:0] ? 5'h0 : _GEN_5; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_7 = 3'h7 == _T_3[2:0] ? w_vn_7 : _GEN_6; // @[FanCtrl.scala 48:{39,39}]
  wire [3:0] _GEN_92174 = {{1'd0}, _T_3[2:0]}; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_8 = 4'h8 == _GEN_92174 ? w_vn_8 : _GEN_7; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_9 = 4'h9 == _GEN_92174 ? 5'h0 : _GEN_8; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_10 = 4'ha == _GEN_92174 ? 5'h0 : _GEN_9; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_11 = 4'hb == _GEN_92174 ? w_vn_11 : _GEN_10; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_12 = 4'hc == _GEN_92174 ? w_vn_12 : _GEN_11; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_13 = 4'hd == _GEN_92174 ? w_vn_13 : _GEN_12; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_14 = 4'he == _GEN_92174 ? 5'h0 : _GEN_13; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_15 = 4'hf == _GEN_92174 ? w_vn_15 : _GEN_14; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_92182 = {{2'd0}, _T_3[2:0]}; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_16 = 5'h10 == _GEN_92182 ? w_vn_16 : _GEN_15; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_17 = 5'h11 == _GEN_92182 ? 5'h0 : _GEN_16; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_18 = 5'h12 == _GEN_92182 ? w_vn_18 : _GEN_17; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_19 = 5'h13 == _GEN_92182 ? 5'h0 : _GEN_18; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_20 = 5'h14 == _GEN_92182 ? 5'h0 : _GEN_19; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_21 = 5'h15 == _GEN_92182 ? 5'h0 : _GEN_20; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_22 = 5'h16 == _GEN_92182 ? 5'h0 : _GEN_21; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_23 = 5'h17 == _GEN_92182 ? w_vn_23 : _GEN_22; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_24 = 5'h18 == _GEN_92182 ? w_vn_24 : _GEN_23; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_25 = 5'h19 == _GEN_92182 ? 5'h0 : _GEN_24; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_26 = 5'h1a == _GEN_92182 ? 5'h0 : _GEN_25; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_27 = 5'h1b == _GEN_92182 ? 5'h0 : _GEN_26; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_28 = 5'h1c == _GEN_92182 ? 5'h0 : _GEN_27; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_29 = 5'h1d == _GEN_92182 ? 5'h0 : _GEN_28; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_30 = 5'h1e == _GEN_92182 ? 5'h0 : _GEN_29; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_31 = 5'h1f == _GEN_92182 ? 5'h0 : _GEN_30; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_35 = 3'h3 == _T_7 ? w_vn_3 : 5'h0; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_36 = 3'h4 == _T_7 ? w_vn_4 : _GEN_35; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_37 = 3'h5 == _T_7 ? 5'h0 : _GEN_36; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_38 = 3'h6 == _T_7 ? 5'h0 : _GEN_37; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_39 = 3'h7 == _T_7 ? w_vn_7 : _GEN_38; // @[FanCtrl.scala 48:{39,39}]
  wire [3:0] _GEN_92198 = {{1'd0}, _T_7}; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_40 = 4'h8 == _GEN_92198 ? w_vn_8 : _GEN_39; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_41 = 4'h9 == _GEN_92198 ? 5'h0 : _GEN_40; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_42 = 4'ha == _GEN_92198 ? 5'h0 : _GEN_41; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_43 = 4'hb == _GEN_92198 ? w_vn_11 : _GEN_42; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_44 = 4'hc == _GEN_92198 ? w_vn_12 : _GEN_43; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_45 = 4'hd == _GEN_92198 ? w_vn_13 : _GEN_44; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_46 = 4'he == _GEN_92198 ? 5'h0 : _GEN_45; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_47 = 4'hf == _GEN_92198 ? w_vn_15 : _GEN_46; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_92206 = {{2'd0}, _T_7}; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_48 = 5'h10 == _GEN_92206 ? w_vn_16 : _GEN_47; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_49 = 5'h11 == _GEN_92206 ? 5'h0 : _GEN_48; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_50 = 5'h12 == _GEN_92206 ? w_vn_18 : _GEN_49; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_51 = 5'h13 == _GEN_92206 ? 5'h0 : _GEN_50; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_52 = 5'h14 == _GEN_92206 ? 5'h0 : _GEN_51; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_53 = 5'h15 == _GEN_92206 ? 5'h0 : _GEN_52; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_54 = 5'h16 == _GEN_92206 ? 5'h0 : _GEN_53; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_55 = 5'h17 == _GEN_92206 ? w_vn_23 : _GEN_54; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_56 = 5'h18 == _GEN_92206 ? w_vn_24 : _GEN_55; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_57 = 5'h19 == _GEN_92206 ? 5'h0 : _GEN_56; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_58 = 5'h1a == _GEN_92206 ? 5'h0 : _GEN_57; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_59 = 5'h1b == _GEN_92206 ? 5'h0 : _GEN_58; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_60 = 5'h1c == _GEN_92206 ? 5'h0 : _GEN_59; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_61 = 5'h1d == _GEN_92206 ? 5'h0 : _GEN_60; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_62 = 5'h1e == _GEN_92206 ? 5'h0 : _GEN_61; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_63 = 5'h1f == _GEN_92206 ? 5'h0 : _GEN_62; // @[FanCtrl.scala 48:{39,39}]
  wire  _T_8 = _GEN_31 == _GEN_63; // @[FanCtrl.scala 48:39]
  wire [2:0] _T_18 = _T_2 + 3'h2; // @[FanCtrl.scala 55:32]
  wire [4:0] _GEN_192 = 3'h3 == _T_18 ? w_vn_3 : 5'h0; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_193 = 3'h4 == _T_18 ? w_vn_4 : _GEN_192; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_194 = 3'h5 == _T_18 ? 5'h0 : _GEN_193; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_195 = 3'h6 == _T_18 ? 5'h0 : _GEN_194; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_196 = 3'h7 == _T_18 ? w_vn_7 : _GEN_195; // @[FanCtrl.scala 54:{41,41}]
  wire [3:0] _GEN_92246 = {{1'd0}, _T_18}; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_197 = 4'h8 == _GEN_92246 ? w_vn_8 : _GEN_196; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_198 = 4'h9 == _GEN_92246 ? 5'h0 : _GEN_197; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_199 = 4'ha == _GEN_92246 ? 5'h0 : _GEN_198; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_200 = 4'hb == _GEN_92246 ? w_vn_11 : _GEN_199; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_201 = 4'hc == _GEN_92246 ? w_vn_12 : _GEN_200; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_202 = 4'hd == _GEN_92246 ? w_vn_13 : _GEN_201; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_203 = 4'he == _GEN_92246 ? 5'h0 : _GEN_202; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_204 = 4'hf == _GEN_92246 ? w_vn_15 : _GEN_203; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_92254 = {{2'd0}, _T_18}; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_205 = 5'h10 == _GEN_92254 ? w_vn_16 : _GEN_204; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_206 = 5'h11 == _GEN_92254 ? 5'h0 : _GEN_205; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_207 = 5'h12 == _GEN_92254 ? w_vn_18 : _GEN_206; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_208 = 5'h13 == _GEN_92254 ? 5'h0 : _GEN_207; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_209 = 5'h14 == _GEN_92254 ? 5'h0 : _GEN_208; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_210 = 5'h15 == _GEN_92254 ? 5'h0 : _GEN_209; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_211 = 5'h16 == _GEN_92254 ? 5'h0 : _GEN_210; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_212 = 5'h17 == _GEN_92254 ? w_vn_23 : _GEN_211; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_213 = 5'h18 == _GEN_92254 ? w_vn_24 : _GEN_212; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_214 = 5'h19 == _GEN_92254 ? 5'h0 : _GEN_213; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_215 = 5'h1a == _GEN_92254 ? 5'h0 : _GEN_214; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_216 = 5'h1b == _GEN_92254 ? 5'h0 : _GEN_215; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_217 = 5'h1c == _GEN_92254 ? 5'h0 : _GEN_216; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_218 = 5'h1d == _GEN_92254 ? 5'h0 : _GEN_217; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_219 = 5'h1e == _GEN_92254 ? 5'h0 : _GEN_218; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_220 = 5'h1f == _GEN_92254 ? 5'h0 : _GEN_219; // @[FanCtrl.scala 54:{41,41}]
  wire  _T_19 = _GEN_63 != _GEN_220; // @[FanCtrl.scala 54:41]
  wire  _T_26 = _GEN_31 != _GEN_63; // @[FanCtrl.scala 56:41]
  wire  _T_27 = _T_19 & _T_26; // @[FanCtrl.scala 55:41]
  wire  _T_34 = _GEN_63 == _GEN_220; // @[FanCtrl.scala 61:48]
  wire  _T_42 = _T_34 & _T_26; // @[FanCtrl.scala 62:46]
  wire [1:0] _GEN_413 = _T_42 ? 2'h3 : 2'h0; // @[FanCtrl.scala 64:48 66:40 69:38]
  wire [2:0] _GEN_414 = _T_27 ? 3'h5 : {{1'd0}, _GEN_413}; // @[FanCtrl.scala 57:42 59:37]
  wire  _GEN_446 = r_valid_1 & _T_8; // @[FanCtrl.scala 47:34]
  wire [2:0] _GEN_477 = r_valid_1 ? _GEN_414 : 3'h0; // @[FanCtrl.scala 47:34 74:33]
  wire [2:0] _T_179 = 2'h2 * 1'h1; // @[FanCtrl.scala 48:25]
  wire [3:0] _T_180 = {{1'd0}, _T_179}; // @[FanCtrl.scala 48:31]
  wire [2:0] _T_184 = _T_179 + 3'h1; // @[FanCtrl.scala 48:58]
  wire [4:0] _GEN_1884 = 3'h3 == _T_180[2:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_1885 = 3'h4 == _T_180[2:0] ? w_vn_4 : _GEN_1884; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_1886 = 3'h5 == _T_180[2:0] ? 5'h0 : _GEN_1885; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_1887 = 3'h6 == _T_180[2:0] ? 5'h0 : _GEN_1886; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_1888 = 3'h7 == _T_180[2:0] ? w_vn_7 : _GEN_1887; // @[FanCtrl.scala 48:{39,39}]
  wire [3:0] _GEN_93134 = {{1'd0}, _T_180[2:0]}; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_1889 = 4'h8 == _GEN_93134 ? w_vn_8 : _GEN_1888; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_1890 = 4'h9 == _GEN_93134 ? 5'h0 : _GEN_1889; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_1891 = 4'ha == _GEN_93134 ? 5'h0 : _GEN_1890; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_1892 = 4'hb == _GEN_93134 ? w_vn_11 : _GEN_1891; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_1893 = 4'hc == _GEN_93134 ? w_vn_12 : _GEN_1892; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_1894 = 4'hd == _GEN_93134 ? w_vn_13 : _GEN_1893; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_1895 = 4'he == _GEN_93134 ? 5'h0 : _GEN_1894; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_1896 = 4'hf == _GEN_93134 ? w_vn_15 : _GEN_1895; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_93142 = {{2'd0}, _T_180[2:0]}; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_1897 = 5'h10 == _GEN_93142 ? w_vn_16 : _GEN_1896; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_1898 = 5'h11 == _GEN_93142 ? 5'h0 : _GEN_1897; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_1899 = 5'h12 == _GEN_93142 ? w_vn_18 : _GEN_1898; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_1900 = 5'h13 == _GEN_93142 ? 5'h0 : _GEN_1899; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_1901 = 5'h14 == _GEN_93142 ? 5'h0 : _GEN_1900; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_1902 = 5'h15 == _GEN_93142 ? 5'h0 : _GEN_1901; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_1903 = 5'h16 == _GEN_93142 ? 5'h0 : _GEN_1902; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_1904 = 5'h17 == _GEN_93142 ? w_vn_23 : _GEN_1903; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_1905 = 5'h18 == _GEN_93142 ? w_vn_24 : _GEN_1904; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_1906 = 5'h19 == _GEN_93142 ? 5'h0 : _GEN_1905; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_1907 = 5'h1a == _GEN_93142 ? 5'h0 : _GEN_1906; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_1908 = 5'h1b == _GEN_93142 ? 5'h0 : _GEN_1907; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_1909 = 5'h1c == _GEN_93142 ? 5'h0 : _GEN_1908; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_1910 = 5'h1d == _GEN_93142 ? 5'h0 : _GEN_1909; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_1911 = 5'h1e == _GEN_93142 ? 5'h0 : _GEN_1910; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_1912 = 5'h1f == _GEN_93142 ? 5'h0 : _GEN_1911; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_1916 = 3'h3 == _T_184 ? w_vn_3 : 5'h0; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_1917 = 3'h4 == _T_184 ? w_vn_4 : _GEN_1916; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_1918 = 3'h5 == _T_184 ? 5'h0 : _GEN_1917; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_1919 = 3'h6 == _T_184 ? 5'h0 : _GEN_1918; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_1920 = 3'h7 == _T_184 ? w_vn_7 : _GEN_1919; // @[FanCtrl.scala 48:{39,39}]
  wire [3:0] _GEN_93158 = {{1'd0}, _T_184}; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_1921 = 4'h8 == _GEN_93158 ? w_vn_8 : _GEN_1920; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_1922 = 4'h9 == _GEN_93158 ? 5'h0 : _GEN_1921; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_1923 = 4'ha == _GEN_93158 ? 5'h0 : _GEN_1922; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_1924 = 4'hb == _GEN_93158 ? w_vn_11 : _GEN_1923; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_1925 = 4'hc == _GEN_93158 ? w_vn_12 : _GEN_1924; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_1926 = 4'hd == _GEN_93158 ? w_vn_13 : _GEN_1925; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_1927 = 4'he == _GEN_93158 ? 5'h0 : _GEN_1926; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_1928 = 4'hf == _GEN_93158 ? w_vn_15 : _GEN_1927; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_93166 = {{2'd0}, _T_184}; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_1929 = 5'h10 == _GEN_93166 ? w_vn_16 : _GEN_1928; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_1930 = 5'h11 == _GEN_93166 ? 5'h0 : _GEN_1929; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_1931 = 5'h12 == _GEN_93166 ? w_vn_18 : _GEN_1930; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_1932 = 5'h13 == _GEN_93166 ? 5'h0 : _GEN_1931; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_1933 = 5'h14 == _GEN_93166 ? 5'h0 : _GEN_1932; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_1934 = 5'h15 == _GEN_93166 ? 5'h0 : _GEN_1933; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_1935 = 5'h16 == _GEN_93166 ? 5'h0 : _GEN_1934; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_1936 = 5'h17 == _GEN_93166 ? w_vn_23 : _GEN_1935; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_1937 = 5'h18 == _GEN_93166 ? w_vn_24 : _GEN_1936; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_1938 = 5'h19 == _GEN_93166 ? 5'h0 : _GEN_1937; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_1939 = 5'h1a == _GEN_93166 ? 5'h0 : _GEN_1938; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_1940 = 5'h1b == _GEN_93166 ? 5'h0 : _GEN_1939; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_1941 = 5'h1c == _GEN_93166 ? 5'h0 : _GEN_1940; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_1942 = 5'h1d == _GEN_93166 ? 5'h0 : _GEN_1941; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_1943 = 5'h1e == _GEN_93166 ? 5'h0 : _GEN_1942; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_1944 = 5'h1f == _GEN_93166 ? 5'h0 : _GEN_1943; // @[FanCtrl.scala 48:{39,39}]
  wire  _T_185 = _GEN_1912 == _GEN_1944; // @[FanCtrl.scala 48:39]
  wire [2:0] _T_195 = _T_179 + 3'h2; // @[FanCtrl.scala 55:32]
  wire [4:0] _GEN_2073 = 3'h3 == _T_195 ? w_vn_3 : 5'h0; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_2074 = 3'h4 == _T_195 ? w_vn_4 : _GEN_2073; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_2075 = 3'h5 == _T_195 ? 5'h0 : _GEN_2074; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_2076 = 3'h6 == _T_195 ? 5'h0 : _GEN_2075; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_2077 = 3'h7 == _T_195 ? w_vn_7 : _GEN_2076; // @[FanCtrl.scala 54:{41,41}]
  wire [3:0] _GEN_93206 = {{1'd0}, _T_195}; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_2078 = 4'h8 == _GEN_93206 ? w_vn_8 : _GEN_2077; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_2079 = 4'h9 == _GEN_93206 ? 5'h0 : _GEN_2078; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_2080 = 4'ha == _GEN_93206 ? 5'h0 : _GEN_2079; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_2081 = 4'hb == _GEN_93206 ? w_vn_11 : _GEN_2080; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_2082 = 4'hc == _GEN_93206 ? w_vn_12 : _GEN_2081; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_2083 = 4'hd == _GEN_93206 ? w_vn_13 : _GEN_2082; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_2084 = 4'he == _GEN_93206 ? 5'h0 : _GEN_2083; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_2085 = 4'hf == _GEN_93206 ? w_vn_15 : _GEN_2084; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_93214 = {{2'd0}, _T_195}; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_2086 = 5'h10 == _GEN_93214 ? w_vn_16 : _GEN_2085; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_2087 = 5'h11 == _GEN_93214 ? 5'h0 : _GEN_2086; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_2088 = 5'h12 == _GEN_93214 ? w_vn_18 : _GEN_2087; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_2089 = 5'h13 == _GEN_93214 ? 5'h0 : _GEN_2088; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_2090 = 5'h14 == _GEN_93214 ? 5'h0 : _GEN_2089; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_2091 = 5'h15 == _GEN_93214 ? 5'h0 : _GEN_2090; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_2092 = 5'h16 == _GEN_93214 ? 5'h0 : _GEN_2091; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_2093 = 5'h17 == _GEN_93214 ? w_vn_23 : _GEN_2092; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_2094 = 5'h18 == _GEN_93214 ? w_vn_24 : _GEN_2093; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_2095 = 5'h19 == _GEN_93214 ? 5'h0 : _GEN_2094; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_2096 = 5'h1a == _GEN_93214 ? 5'h0 : _GEN_2095; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_2097 = 5'h1b == _GEN_93214 ? 5'h0 : _GEN_2096; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_2098 = 5'h1c == _GEN_93214 ? 5'h0 : _GEN_2097; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_2099 = 5'h1d == _GEN_93214 ? 5'h0 : _GEN_2098; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_2100 = 5'h1e == _GEN_93214 ? 5'h0 : _GEN_2099; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_2101 = 5'h1f == _GEN_93214 ? 5'h0 : _GEN_2100; // @[FanCtrl.scala 54:{41,41}]
  wire  _T_196 = _GEN_1944 != _GEN_2101; // @[FanCtrl.scala 54:41]
  wire  _T_203 = _GEN_1912 != _GEN_1944; // @[FanCtrl.scala 56:41]
  wire  _T_211 = _GEN_1944 == _GEN_2101; // @[FanCtrl.scala 61:48]
  wire  _GEN_2328 = r_valid_1 & _T_185; // @[FanCtrl.scala 47:34]
  wire [2:0] _T_242 = _T_179 - 3'h1; // @[FanCtrl.scala 94:58]
  wire [4:0] _GEN_2582 = 3'h3 == _T_242 ? w_vn_3 : 5'h0; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_2583 = 3'h4 == _T_242 ? w_vn_4 : _GEN_2582; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_2584 = 3'h5 == _T_242 ? 5'h0 : _GEN_2583; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_2585 = 3'h6 == _T_242 ? 5'h0 : _GEN_2584; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_2586 = 3'h7 == _T_242 ? w_vn_7 : _GEN_2585; // @[FanCtrl.scala 94:{39,39}]
  wire [3:0] _GEN_93446 = {{1'd0}, _T_242}; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_2587 = 4'h8 == _GEN_93446 ? w_vn_8 : _GEN_2586; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_2588 = 4'h9 == _GEN_93446 ? 5'h0 : _GEN_2587; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_2589 = 4'ha == _GEN_93446 ? 5'h0 : _GEN_2588; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_2590 = 4'hb == _GEN_93446 ? w_vn_11 : _GEN_2589; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_2591 = 4'hc == _GEN_93446 ? w_vn_12 : _GEN_2590; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_2592 = 4'hd == _GEN_93446 ? w_vn_13 : _GEN_2591; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_2593 = 4'he == _GEN_93446 ? 5'h0 : _GEN_2592; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_2594 = 4'hf == _GEN_93446 ? w_vn_15 : _GEN_2593; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_93454 = {{2'd0}, _T_242}; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_2595 = 5'h10 == _GEN_93454 ? w_vn_16 : _GEN_2594; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_2596 = 5'h11 == _GEN_93454 ? 5'h0 : _GEN_2595; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_2597 = 5'h12 == _GEN_93454 ? w_vn_18 : _GEN_2596; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_2598 = 5'h13 == _GEN_93454 ? 5'h0 : _GEN_2597; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_2599 = 5'h14 == _GEN_93454 ? 5'h0 : _GEN_2598; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_2600 = 5'h15 == _GEN_93454 ? 5'h0 : _GEN_2599; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_2601 = 5'h16 == _GEN_93454 ? 5'h0 : _GEN_2600; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_2602 = 5'h17 == _GEN_93454 ? w_vn_23 : _GEN_2601; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_2603 = 5'h18 == _GEN_93454 ? w_vn_24 : _GEN_2602; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_2604 = 5'h19 == _GEN_93454 ? 5'h0 : _GEN_2603; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_2605 = 5'h1a == _GEN_93454 ? 5'h0 : _GEN_2604; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_2606 = 5'h1b == _GEN_93454 ? 5'h0 : _GEN_2605; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_2607 = 5'h1c == _GEN_93454 ? 5'h0 : _GEN_2606; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_2608 = 5'h1d == _GEN_93454 ? 5'h0 : _GEN_2607; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_2609 = 5'h1e == _GEN_93454 ? 5'h0 : _GEN_2608; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_2610 = 5'h1f == _GEN_93454 ? 5'h0 : _GEN_2609; // @[FanCtrl.scala 94:{39,39}]
  wire  _T_243 = _GEN_1912 != _GEN_2610; // @[FanCtrl.scala 94:39]
  wire  _T_258 = _GEN_1912 == _GEN_2610; // @[FanCtrl.scala 99:46]
  wire  _T_297 = _T_243 & _T_196; // @[FanCtrl.scala 125:65]
  wire  _T_305 = _T_297 & _T_203; // @[FanCtrl.scala 126:65]
  wire  _T_320 = _T_258 & _T_196; // @[FanCtrl.scala 131:70]
  wire  _T_328 = _T_320 & _T_203; // @[FanCtrl.scala 132:72]
  wire  _T_343 = _T_243 & _T_211; // @[FanCtrl.scala 137:72]
  wire  _T_351 = _T_343 & _T_203; // @[FanCtrl.scala 138:71]
  wire [1:0] _GEN_3632 = _T_351 ? 2'h3 : 2'h1; // @[FanCtrl.scala 139:73 141:34 144:35]
  wire [2:0] _GEN_3633 = _T_328 ? 3'h4 : {{1'd0}, _GEN_3632}; // @[FanCtrl.scala 133:73 135:35]
  wire [2:0] _GEN_3634 = _T_305 ? 3'h5 : _GEN_3633; // @[FanCtrl.scala 127:66 129:35]
  wire [2:0] _GEN_3697 = r_valid_1 ? _GEN_3634 : 3'h0; // @[FanCtrl.scala 117:32 148:33]
  wire [3:0] _T_356 = 2'h2 * 2'h2; // @[FanCtrl.scala 48:25]
  wire [4:0] _T_357 = {{1'd0}, _T_356}; // @[FanCtrl.scala 48:31]
  wire [3:0] _T_361 = _T_356 + 4'h1; // @[FanCtrl.scala 48:58]
  wire [4:0] _GEN_3766 = 4'h3 == _T_357[3:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_3767 = 4'h4 == _T_357[3:0] ? w_vn_4 : _GEN_3766; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_3768 = 4'h5 == _T_357[3:0] ? 5'h0 : _GEN_3767; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_3769 = 4'h6 == _T_357[3:0] ? 5'h0 : _GEN_3768; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_3770 = 4'h7 == _T_357[3:0] ? w_vn_7 : _GEN_3769; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_3771 = 4'h8 == _T_357[3:0] ? w_vn_8 : _GEN_3770; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_3772 = 4'h9 == _T_357[3:0] ? 5'h0 : _GEN_3771; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_3773 = 4'ha == _T_357[3:0] ? 5'h0 : _GEN_3772; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_3774 = 4'hb == _T_357[3:0] ? w_vn_11 : _GEN_3773; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_3775 = 4'hc == _T_357[3:0] ? w_vn_12 : _GEN_3774; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_3776 = 4'hd == _T_357[3:0] ? w_vn_13 : _GEN_3775; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_3777 = 4'he == _T_357[3:0] ? 5'h0 : _GEN_3776; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_3778 = 4'hf == _T_357[3:0] ? w_vn_15 : _GEN_3777; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_94094 = {{1'd0}, _T_357[3:0]}; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_3779 = 5'h10 == _GEN_94094 ? w_vn_16 : _GEN_3778; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_3780 = 5'h11 == _GEN_94094 ? 5'h0 : _GEN_3779; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_3781 = 5'h12 == _GEN_94094 ? w_vn_18 : _GEN_3780; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_3782 = 5'h13 == _GEN_94094 ? 5'h0 : _GEN_3781; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_3783 = 5'h14 == _GEN_94094 ? 5'h0 : _GEN_3782; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_3784 = 5'h15 == _GEN_94094 ? 5'h0 : _GEN_3783; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_3785 = 5'h16 == _GEN_94094 ? 5'h0 : _GEN_3784; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_3786 = 5'h17 == _GEN_94094 ? w_vn_23 : _GEN_3785; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_3787 = 5'h18 == _GEN_94094 ? w_vn_24 : _GEN_3786; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_3788 = 5'h19 == _GEN_94094 ? 5'h0 : _GEN_3787; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_3789 = 5'h1a == _GEN_94094 ? 5'h0 : _GEN_3788; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_3790 = 5'h1b == _GEN_94094 ? 5'h0 : _GEN_3789; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_3791 = 5'h1c == _GEN_94094 ? 5'h0 : _GEN_3790; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_3792 = 5'h1d == _GEN_94094 ? 5'h0 : _GEN_3791; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_3793 = 5'h1e == _GEN_94094 ? 5'h0 : _GEN_3792; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_3794 = 5'h1f == _GEN_94094 ? 5'h0 : _GEN_3793; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_3798 = 4'h3 == _T_361 ? w_vn_3 : 5'h0; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_3799 = 4'h4 == _T_361 ? w_vn_4 : _GEN_3798; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_3800 = 4'h5 == _T_361 ? 5'h0 : _GEN_3799; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_3801 = 4'h6 == _T_361 ? 5'h0 : _GEN_3800; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_3802 = 4'h7 == _T_361 ? w_vn_7 : _GEN_3801; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_3803 = 4'h8 == _T_361 ? w_vn_8 : _GEN_3802; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_3804 = 4'h9 == _T_361 ? 5'h0 : _GEN_3803; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_3805 = 4'ha == _T_361 ? 5'h0 : _GEN_3804; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_3806 = 4'hb == _T_361 ? w_vn_11 : _GEN_3805; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_3807 = 4'hc == _T_361 ? w_vn_12 : _GEN_3806; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_3808 = 4'hd == _T_361 ? w_vn_13 : _GEN_3807; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_3809 = 4'he == _T_361 ? 5'h0 : _GEN_3808; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_3810 = 4'hf == _T_361 ? w_vn_15 : _GEN_3809; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_94110 = {{1'd0}, _T_361}; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_3811 = 5'h10 == _GEN_94110 ? w_vn_16 : _GEN_3810; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_3812 = 5'h11 == _GEN_94110 ? 5'h0 : _GEN_3811; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_3813 = 5'h12 == _GEN_94110 ? w_vn_18 : _GEN_3812; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_3814 = 5'h13 == _GEN_94110 ? 5'h0 : _GEN_3813; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_3815 = 5'h14 == _GEN_94110 ? 5'h0 : _GEN_3814; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_3816 = 5'h15 == _GEN_94110 ? 5'h0 : _GEN_3815; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_3817 = 5'h16 == _GEN_94110 ? 5'h0 : _GEN_3816; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_3818 = 5'h17 == _GEN_94110 ? w_vn_23 : _GEN_3817; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_3819 = 5'h18 == _GEN_94110 ? w_vn_24 : _GEN_3818; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_3820 = 5'h19 == _GEN_94110 ? 5'h0 : _GEN_3819; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_3821 = 5'h1a == _GEN_94110 ? 5'h0 : _GEN_3820; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_3822 = 5'h1b == _GEN_94110 ? 5'h0 : _GEN_3821; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_3823 = 5'h1c == _GEN_94110 ? 5'h0 : _GEN_3822; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_3824 = 5'h1d == _GEN_94110 ? 5'h0 : _GEN_3823; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_3825 = 5'h1e == _GEN_94110 ? 5'h0 : _GEN_3824; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_3826 = 5'h1f == _GEN_94110 ? 5'h0 : _GEN_3825; // @[FanCtrl.scala 48:{39,39}]
  wire  _T_362 = _GEN_3794 == _GEN_3826; // @[FanCtrl.scala 48:39]
  wire [3:0] _T_372 = _T_356 + 4'h2; // @[FanCtrl.scala 55:32]
  wire [4:0] _GEN_3955 = 4'h3 == _T_372 ? w_vn_3 : 5'h0; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_3956 = 4'h4 == _T_372 ? w_vn_4 : _GEN_3955; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_3957 = 4'h5 == _T_372 ? 5'h0 : _GEN_3956; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_3958 = 4'h6 == _T_372 ? 5'h0 : _GEN_3957; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_3959 = 4'h7 == _T_372 ? w_vn_7 : _GEN_3958; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_3960 = 4'h8 == _T_372 ? w_vn_8 : _GEN_3959; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_3961 = 4'h9 == _T_372 ? 5'h0 : _GEN_3960; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_3962 = 4'ha == _T_372 ? 5'h0 : _GEN_3961; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_3963 = 4'hb == _T_372 ? w_vn_11 : _GEN_3962; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_3964 = 4'hc == _T_372 ? w_vn_12 : _GEN_3963; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_3965 = 4'hd == _T_372 ? w_vn_13 : _GEN_3964; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_3966 = 4'he == _T_372 ? 5'h0 : _GEN_3965; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_3967 = 4'hf == _T_372 ? w_vn_15 : _GEN_3966; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_94142 = {{1'd0}, _T_372}; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_3968 = 5'h10 == _GEN_94142 ? w_vn_16 : _GEN_3967; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_3969 = 5'h11 == _GEN_94142 ? 5'h0 : _GEN_3968; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_3970 = 5'h12 == _GEN_94142 ? w_vn_18 : _GEN_3969; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_3971 = 5'h13 == _GEN_94142 ? 5'h0 : _GEN_3970; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_3972 = 5'h14 == _GEN_94142 ? 5'h0 : _GEN_3971; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_3973 = 5'h15 == _GEN_94142 ? 5'h0 : _GEN_3972; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_3974 = 5'h16 == _GEN_94142 ? 5'h0 : _GEN_3973; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_3975 = 5'h17 == _GEN_94142 ? w_vn_23 : _GEN_3974; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_3976 = 5'h18 == _GEN_94142 ? w_vn_24 : _GEN_3975; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_3977 = 5'h19 == _GEN_94142 ? 5'h0 : _GEN_3976; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_3978 = 5'h1a == _GEN_94142 ? 5'h0 : _GEN_3977; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_3979 = 5'h1b == _GEN_94142 ? 5'h0 : _GEN_3978; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_3980 = 5'h1c == _GEN_94142 ? 5'h0 : _GEN_3979; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_3981 = 5'h1d == _GEN_94142 ? 5'h0 : _GEN_3980; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_3982 = 5'h1e == _GEN_94142 ? 5'h0 : _GEN_3981; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_3983 = 5'h1f == _GEN_94142 ? 5'h0 : _GEN_3982; // @[FanCtrl.scala 54:{41,41}]
  wire  _T_373 = _GEN_3826 != _GEN_3983; // @[FanCtrl.scala 54:41]
  wire  _T_380 = _GEN_3794 != _GEN_3826; // @[FanCtrl.scala 56:41]
  wire  _T_388 = _GEN_3826 == _GEN_3983; // @[FanCtrl.scala 61:48]
  wire  _GEN_4211 = r_valid_1 & _T_362; // @[FanCtrl.scala 47:34]
  wire [3:0] _T_419 = _T_356 - 4'h1; // @[FanCtrl.scala 94:58]
  wire [4:0] _GEN_4464 = 4'h3 == _T_419 ? w_vn_3 : 5'h0; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_4465 = 4'h4 == _T_419 ? w_vn_4 : _GEN_4464; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_4466 = 4'h5 == _T_419 ? 5'h0 : _GEN_4465; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_4467 = 4'h6 == _T_419 ? 5'h0 : _GEN_4466; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_4468 = 4'h7 == _T_419 ? w_vn_7 : _GEN_4467; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_4469 = 4'h8 == _T_419 ? w_vn_8 : _GEN_4468; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_4470 = 4'h9 == _T_419 ? 5'h0 : _GEN_4469; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_4471 = 4'ha == _T_419 ? 5'h0 : _GEN_4470; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_4472 = 4'hb == _T_419 ? w_vn_11 : _GEN_4471; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_4473 = 4'hc == _T_419 ? w_vn_12 : _GEN_4472; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_4474 = 4'hd == _T_419 ? w_vn_13 : _GEN_4473; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_4475 = 4'he == _T_419 ? 5'h0 : _GEN_4474; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_4476 = 4'hf == _T_419 ? w_vn_15 : _GEN_4475; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_94302 = {{1'd0}, _T_419}; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_4477 = 5'h10 == _GEN_94302 ? w_vn_16 : _GEN_4476; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_4478 = 5'h11 == _GEN_94302 ? 5'h0 : _GEN_4477; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_4479 = 5'h12 == _GEN_94302 ? w_vn_18 : _GEN_4478; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_4480 = 5'h13 == _GEN_94302 ? 5'h0 : _GEN_4479; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_4481 = 5'h14 == _GEN_94302 ? 5'h0 : _GEN_4480; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_4482 = 5'h15 == _GEN_94302 ? 5'h0 : _GEN_4481; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_4483 = 5'h16 == _GEN_94302 ? 5'h0 : _GEN_4482; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_4484 = 5'h17 == _GEN_94302 ? w_vn_23 : _GEN_4483; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_4485 = 5'h18 == _GEN_94302 ? w_vn_24 : _GEN_4484; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_4486 = 5'h19 == _GEN_94302 ? 5'h0 : _GEN_4485; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_4487 = 5'h1a == _GEN_94302 ? 5'h0 : _GEN_4486; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_4488 = 5'h1b == _GEN_94302 ? 5'h0 : _GEN_4487; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_4489 = 5'h1c == _GEN_94302 ? 5'h0 : _GEN_4488; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_4490 = 5'h1d == _GEN_94302 ? 5'h0 : _GEN_4489; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_4491 = 5'h1e == _GEN_94302 ? 5'h0 : _GEN_4490; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_4492 = 5'h1f == _GEN_94302 ? 5'h0 : _GEN_4491; // @[FanCtrl.scala 94:{39,39}]
  wire  _T_420 = _GEN_3794 != _GEN_4492; // @[FanCtrl.scala 94:39]
  wire  _T_435 = _GEN_3794 == _GEN_4492; // @[FanCtrl.scala 99:46]
  wire  _T_474 = _T_420 & _T_373; // @[FanCtrl.scala 125:65]
  wire  _T_482 = _T_474 & _T_380; // @[FanCtrl.scala 126:65]
  wire  _T_497 = _T_435 & _T_373; // @[FanCtrl.scala 131:70]
  wire  _T_505 = _T_497 & _T_380; // @[FanCtrl.scala 132:72]
  wire  _T_520 = _T_420 & _T_388; // @[FanCtrl.scala 137:72]
  wire  _T_528 = _T_520 & _T_380; // @[FanCtrl.scala 138:71]
  wire [1:0] _GEN_5514 = _T_528 ? 2'h3 : 2'h1; // @[FanCtrl.scala 139:73 141:34 144:35]
  wire [2:0] _GEN_5515 = _T_505 ? 3'h4 : {{1'd0}, _GEN_5514}; // @[FanCtrl.scala 133:73 135:35]
  wire [2:0] _GEN_5516 = _T_482 ? 3'h5 : _GEN_5515; // @[FanCtrl.scala 127:66 129:35]
  wire [2:0] _GEN_5579 = r_valid_1 ? _GEN_5516 : 3'h0; // @[FanCtrl.scala 117:32 148:33]
  wire [3:0] _T_533 = 2'h2 * 2'h3; // @[FanCtrl.scala 48:25]
  wire [4:0] _T_534 = {{1'd0}, _T_533}; // @[FanCtrl.scala 48:31]
  wire [3:0] _T_538 = _T_533 + 4'h1; // @[FanCtrl.scala 48:58]
  wire [4:0] _GEN_5648 = 4'h3 == _T_534[3:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_5649 = 4'h4 == _T_534[3:0] ? w_vn_4 : _GEN_5648; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_5650 = 4'h5 == _T_534[3:0] ? 5'h0 : _GEN_5649; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_5651 = 4'h6 == _T_534[3:0] ? 5'h0 : _GEN_5650; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_5652 = 4'h7 == _T_534[3:0] ? w_vn_7 : _GEN_5651; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_5653 = 4'h8 == _T_534[3:0] ? w_vn_8 : _GEN_5652; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_5654 = 4'h9 == _T_534[3:0] ? 5'h0 : _GEN_5653; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_5655 = 4'ha == _T_534[3:0] ? 5'h0 : _GEN_5654; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_5656 = 4'hb == _T_534[3:0] ? w_vn_11 : _GEN_5655; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_5657 = 4'hc == _T_534[3:0] ? w_vn_12 : _GEN_5656; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_5658 = 4'hd == _T_534[3:0] ? w_vn_13 : _GEN_5657; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_5659 = 4'he == _T_534[3:0] ? 5'h0 : _GEN_5658; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_5660 = 4'hf == _T_534[3:0] ? w_vn_15 : _GEN_5659; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_94734 = {{1'd0}, _T_534[3:0]}; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_5661 = 5'h10 == _GEN_94734 ? w_vn_16 : _GEN_5660; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_5662 = 5'h11 == _GEN_94734 ? 5'h0 : _GEN_5661; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_5663 = 5'h12 == _GEN_94734 ? w_vn_18 : _GEN_5662; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_5664 = 5'h13 == _GEN_94734 ? 5'h0 : _GEN_5663; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_5665 = 5'h14 == _GEN_94734 ? 5'h0 : _GEN_5664; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_5666 = 5'h15 == _GEN_94734 ? 5'h0 : _GEN_5665; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_5667 = 5'h16 == _GEN_94734 ? 5'h0 : _GEN_5666; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_5668 = 5'h17 == _GEN_94734 ? w_vn_23 : _GEN_5667; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_5669 = 5'h18 == _GEN_94734 ? w_vn_24 : _GEN_5668; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_5670 = 5'h19 == _GEN_94734 ? 5'h0 : _GEN_5669; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_5671 = 5'h1a == _GEN_94734 ? 5'h0 : _GEN_5670; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_5672 = 5'h1b == _GEN_94734 ? 5'h0 : _GEN_5671; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_5673 = 5'h1c == _GEN_94734 ? 5'h0 : _GEN_5672; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_5674 = 5'h1d == _GEN_94734 ? 5'h0 : _GEN_5673; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_5675 = 5'h1e == _GEN_94734 ? 5'h0 : _GEN_5674; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_5676 = 5'h1f == _GEN_94734 ? 5'h0 : _GEN_5675; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_5680 = 4'h3 == _T_538 ? w_vn_3 : 5'h0; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_5681 = 4'h4 == _T_538 ? w_vn_4 : _GEN_5680; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_5682 = 4'h5 == _T_538 ? 5'h0 : _GEN_5681; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_5683 = 4'h6 == _T_538 ? 5'h0 : _GEN_5682; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_5684 = 4'h7 == _T_538 ? w_vn_7 : _GEN_5683; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_5685 = 4'h8 == _T_538 ? w_vn_8 : _GEN_5684; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_5686 = 4'h9 == _T_538 ? 5'h0 : _GEN_5685; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_5687 = 4'ha == _T_538 ? 5'h0 : _GEN_5686; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_5688 = 4'hb == _T_538 ? w_vn_11 : _GEN_5687; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_5689 = 4'hc == _T_538 ? w_vn_12 : _GEN_5688; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_5690 = 4'hd == _T_538 ? w_vn_13 : _GEN_5689; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_5691 = 4'he == _T_538 ? 5'h0 : _GEN_5690; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_5692 = 4'hf == _T_538 ? w_vn_15 : _GEN_5691; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_94750 = {{1'd0}, _T_538}; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_5693 = 5'h10 == _GEN_94750 ? w_vn_16 : _GEN_5692; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_5694 = 5'h11 == _GEN_94750 ? 5'h0 : _GEN_5693; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_5695 = 5'h12 == _GEN_94750 ? w_vn_18 : _GEN_5694; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_5696 = 5'h13 == _GEN_94750 ? 5'h0 : _GEN_5695; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_5697 = 5'h14 == _GEN_94750 ? 5'h0 : _GEN_5696; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_5698 = 5'h15 == _GEN_94750 ? 5'h0 : _GEN_5697; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_5699 = 5'h16 == _GEN_94750 ? 5'h0 : _GEN_5698; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_5700 = 5'h17 == _GEN_94750 ? w_vn_23 : _GEN_5699; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_5701 = 5'h18 == _GEN_94750 ? w_vn_24 : _GEN_5700; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_5702 = 5'h19 == _GEN_94750 ? 5'h0 : _GEN_5701; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_5703 = 5'h1a == _GEN_94750 ? 5'h0 : _GEN_5702; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_5704 = 5'h1b == _GEN_94750 ? 5'h0 : _GEN_5703; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_5705 = 5'h1c == _GEN_94750 ? 5'h0 : _GEN_5704; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_5706 = 5'h1d == _GEN_94750 ? 5'h0 : _GEN_5705; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_5707 = 5'h1e == _GEN_94750 ? 5'h0 : _GEN_5706; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_5708 = 5'h1f == _GEN_94750 ? 5'h0 : _GEN_5707; // @[FanCtrl.scala 48:{39,39}]
  wire  _T_539 = _GEN_5676 == _GEN_5708; // @[FanCtrl.scala 48:39]
  wire [3:0] _T_549 = _T_533 + 4'h2; // @[FanCtrl.scala 55:32]
  wire [4:0] _GEN_5837 = 4'h3 == _T_549 ? w_vn_3 : 5'h0; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_5838 = 4'h4 == _T_549 ? w_vn_4 : _GEN_5837; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_5839 = 4'h5 == _T_549 ? 5'h0 : _GEN_5838; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_5840 = 4'h6 == _T_549 ? 5'h0 : _GEN_5839; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_5841 = 4'h7 == _T_549 ? w_vn_7 : _GEN_5840; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_5842 = 4'h8 == _T_549 ? w_vn_8 : _GEN_5841; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_5843 = 4'h9 == _T_549 ? 5'h0 : _GEN_5842; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_5844 = 4'ha == _T_549 ? 5'h0 : _GEN_5843; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_5845 = 4'hb == _T_549 ? w_vn_11 : _GEN_5844; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_5846 = 4'hc == _T_549 ? w_vn_12 : _GEN_5845; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_5847 = 4'hd == _T_549 ? w_vn_13 : _GEN_5846; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_5848 = 4'he == _T_549 ? 5'h0 : _GEN_5847; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_5849 = 4'hf == _T_549 ? w_vn_15 : _GEN_5848; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_94782 = {{1'd0}, _T_549}; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_5850 = 5'h10 == _GEN_94782 ? w_vn_16 : _GEN_5849; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_5851 = 5'h11 == _GEN_94782 ? 5'h0 : _GEN_5850; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_5852 = 5'h12 == _GEN_94782 ? w_vn_18 : _GEN_5851; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_5853 = 5'h13 == _GEN_94782 ? 5'h0 : _GEN_5852; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_5854 = 5'h14 == _GEN_94782 ? 5'h0 : _GEN_5853; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_5855 = 5'h15 == _GEN_94782 ? 5'h0 : _GEN_5854; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_5856 = 5'h16 == _GEN_94782 ? 5'h0 : _GEN_5855; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_5857 = 5'h17 == _GEN_94782 ? w_vn_23 : _GEN_5856; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_5858 = 5'h18 == _GEN_94782 ? w_vn_24 : _GEN_5857; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_5859 = 5'h19 == _GEN_94782 ? 5'h0 : _GEN_5858; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_5860 = 5'h1a == _GEN_94782 ? 5'h0 : _GEN_5859; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_5861 = 5'h1b == _GEN_94782 ? 5'h0 : _GEN_5860; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_5862 = 5'h1c == _GEN_94782 ? 5'h0 : _GEN_5861; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_5863 = 5'h1d == _GEN_94782 ? 5'h0 : _GEN_5862; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_5864 = 5'h1e == _GEN_94782 ? 5'h0 : _GEN_5863; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_5865 = 5'h1f == _GEN_94782 ? 5'h0 : _GEN_5864; // @[FanCtrl.scala 54:{41,41}]
  wire  _T_550 = _GEN_5708 != _GEN_5865; // @[FanCtrl.scala 54:41]
  wire  _T_557 = _GEN_5676 != _GEN_5708; // @[FanCtrl.scala 56:41]
  wire  _T_565 = _GEN_5708 == _GEN_5865; // @[FanCtrl.scala 61:48]
  wire  _GEN_6094 = r_valid_1 & _T_539; // @[FanCtrl.scala 47:34]
  wire [3:0] _T_596 = _T_533 - 4'h1; // @[FanCtrl.scala 94:58]
  wire [4:0] _GEN_6346 = 4'h3 == _T_596 ? w_vn_3 : 5'h0; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_6347 = 4'h4 == _T_596 ? w_vn_4 : _GEN_6346; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_6348 = 4'h5 == _T_596 ? 5'h0 : _GEN_6347; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_6349 = 4'h6 == _T_596 ? 5'h0 : _GEN_6348; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_6350 = 4'h7 == _T_596 ? w_vn_7 : _GEN_6349; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_6351 = 4'h8 == _T_596 ? w_vn_8 : _GEN_6350; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_6352 = 4'h9 == _T_596 ? 5'h0 : _GEN_6351; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_6353 = 4'ha == _T_596 ? 5'h0 : _GEN_6352; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_6354 = 4'hb == _T_596 ? w_vn_11 : _GEN_6353; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_6355 = 4'hc == _T_596 ? w_vn_12 : _GEN_6354; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_6356 = 4'hd == _T_596 ? w_vn_13 : _GEN_6355; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_6357 = 4'he == _T_596 ? 5'h0 : _GEN_6356; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_6358 = 4'hf == _T_596 ? w_vn_15 : _GEN_6357; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_94942 = {{1'd0}, _T_596}; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_6359 = 5'h10 == _GEN_94942 ? w_vn_16 : _GEN_6358; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_6360 = 5'h11 == _GEN_94942 ? 5'h0 : _GEN_6359; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_6361 = 5'h12 == _GEN_94942 ? w_vn_18 : _GEN_6360; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_6362 = 5'h13 == _GEN_94942 ? 5'h0 : _GEN_6361; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_6363 = 5'h14 == _GEN_94942 ? 5'h0 : _GEN_6362; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_6364 = 5'h15 == _GEN_94942 ? 5'h0 : _GEN_6363; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_6365 = 5'h16 == _GEN_94942 ? 5'h0 : _GEN_6364; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_6366 = 5'h17 == _GEN_94942 ? w_vn_23 : _GEN_6365; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_6367 = 5'h18 == _GEN_94942 ? w_vn_24 : _GEN_6366; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_6368 = 5'h19 == _GEN_94942 ? 5'h0 : _GEN_6367; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_6369 = 5'h1a == _GEN_94942 ? 5'h0 : _GEN_6368; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_6370 = 5'h1b == _GEN_94942 ? 5'h0 : _GEN_6369; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_6371 = 5'h1c == _GEN_94942 ? 5'h0 : _GEN_6370; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_6372 = 5'h1d == _GEN_94942 ? 5'h0 : _GEN_6371; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_6373 = 5'h1e == _GEN_94942 ? 5'h0 : _GEN_6372; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_6374 = 5'h1f == _GEN_94942 ? 5'h0 : _GEN_6373; // @[FanCtrl.scala 94:{39,39}]
  wire  _T_597 = _GEN_5676 != _GEN_6374; // @[FanCtrl.scala 94:39]
  wire  _T_612 = _GEN_5676 == _GEN_6374; // @[FanCtrl.scala 99:46]
  wire  _T_651 = _T_597 & _T_550; // @[FanCtrl.scala 125:65]
  wire  _T_659 = _T_651 & _T_557; // @[FanCtrl.scala 126:65]
  wire  _T_674 = _T_612 & _T_550; // @[FanCtrl.scala 131:70]
  wire  _T_682 = _T_674 & _T_557; // @[FanCtrl.scala 132:72]
  wire  _T_697 = _T_597 & _T_565; // @[FanCtrl.scala 137:72]
  wire  _T_705 = _T_697 & _T_557; // @[FanCtrl.scala 138:71]
  wire [1:0] _GEN_7396 = _T_705 ? 2'h3 : 2'h1; // @[FanCtrl.scala 139:73 141:34 144:35]
  wire [2:0] _GEN_7397 = _T_682 ? 3'h4 : {{1'd0}, _GEN_7396}; // @[FanCtrl.scala 133:73 135:35]
  wire [2:0] _GEN_7398 = _T_659 ? 3'h5 : _GEN_7397; // @[FanCtrl.scala 127:66 129:35]
  wire [2:0] _GEN_7461 = r_valid_1 ? _GEN_7398 : 3'h0; // @[FanCtrl.scala 117:32 148:33]
  wire [4:0] _T_710 = 2'h2 * 3'h4; // @[FanCtrl.scala 48:25]
  wire [5:0] _T_711 = {{1'd0}, _T_710}; // @[FanCtrl.scala 48:31]
  wire [4:0] _T_715 = _T_710 + 5'h1; // @[FanCtrl.scala 48:58]
  wire [4:0] _GEN_7530 = 5'h3 == _T_711[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_7531 = 5'h4 == _T_711[4:0] ? w_vn_4 : _GEN_7530; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_7532 = 5'h5 == _T_711[4:0] ? 5'h0 : _GEN_7531; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_7533 = 5'h6 == _T_711[4:0] ? 5'h0 : _GEN_7532; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_7534 = 5'h7 == _T_711[4:0] ? w_vn_7 : _GEN_7533; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_7535 = 5'h8 == _T_711[4:0] ? w_vn_8 : _GEN_7534; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_7536 = 5'h9 == _T_711[4:0] ? 5'h0 : _GEN_7535; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_7537 = 5'ha == _T_711[4:0] ? 5'h0 : _GEN_7536; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_7538 = 5'hb == _T_711[4:0] ? w_vn_11 : _GEN_7537; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_7539 = 5'hc == _T_711[4:0] ? w_vn_12 : _GEN_7538; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_7540 = 5'hd == _T_711[4:0] ? w_vn_13 : _GEN_7539; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_7541 = 5'he == _T_711[4:0] ? 5'h0 : _GEN_7540; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_7542 = 5'hf == _T_711[4:0] ? w_vn_15 : _GEN_7541; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_7543 = 5'h10 == _T_711[4:0] ? w_vn_16 : _GEN_7542; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_7544 = 5'h11 == _T_711[4:0] ? 5'h0 : _GEN_7543; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_7545 = 5'h12 == _T_711[4:0] ? w_vn_18 : _GEN_7544; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_7546 = 5'h13 == _T_711[4:0] ? 5'h0 : _GEN_7545; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_7547 = 5'h14 == _T_711[4:0] ? 5'h0 : _GEN_7546; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_7548 = 5'h15 == _T_711[4:0] ? 5'h0 : _GEN_7547; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_7549 = 5'h16 == _T_711[4:0] ? 5'h0 : _GEN_7548; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_7550 = 5'h17 == _T_711[4:0] ? w_vn_23 : _GEN_7549; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_7551 = 5'h18 == _T_711[4:0] ? w_vn_24 : _GEN_7550; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_7552 = 5'h19 == _T_711[4:0] ? 5'h0 : _GEN_7551; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_7553 = 5'h1a == _T_711[4:0] ? 5'h0 : _GEN_7552; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_7554 = 5'h1b == _T_711[4:0] ? 5'h0 : _GEN_7553; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_7555 = 5'h1c == _T_711[4:0] ? 5'h0 : _GEN_7554; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_7556 = 5'h1d == _T_711[4:0] ? 5'h0 : _GEN_7555; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_7557 = 5'h1e == _T_711[4:0] ? 5'h0 : _GEN_7556; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_7558 = 5'h1f == _T_711[4:0] ? 5'h0 : _GEN_7557; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_7562 = 5'h3 == _T_715 ? w_vn_3 : 5'h0; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_7563 = 5'h4 == _T_715 ? w_vn_4 : _GEN_7562; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_7564 = 5'h5 == _T_715 ? 5'h0 : _GEN_7563; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_7565 = 5'h6 == _T_715 ? 5'h0 : _GEN_7564; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_7566 = 5'h7 == _T_715 ? w_vn_7 : _GEN_7565; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_7567 = 5'h8 == _T_715 ? w_vn_8 : _GEN_7566; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_7568 = 5'h9 == _T_715 ? 5'h0 : _GEN_7567; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_7569 = 5'ha == _T_715 ? 5'h0 : _GEN_7568; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_7570 = 5'hb == _T_715 ? w_vn_11 : _GEN_7569; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_7571 = 5'hc == _T_715 ? w_vn_12 : _GEN_7570; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_7572 = 5'hd == _T_715 ? w_vn_13 : _GEN_7571; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_7573 = 5'he == _T_715 ? 5'h0 : _GEN_7572; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_7574 = 5'hf == _T_715 ? w_vn_15 : _GEN_7573; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_7575 = 5'h10 == _T_715 ? w_vn_16 : _GEN_7574; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_7576 = 5'h11 == _T_715 ? 5'h0 : _GEN_7575; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_7577 = 5'h12 == _T_715 ? w_vn_18 : _GEN_7576; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_7578 = 5'h13 == _T_715 ? 5'h0 : _GEN_7577; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_7579 = 5'h14 == _T_715 ? 5'h0 : _GEN_7578; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_7580 = 5'h15 == _T_715 ? 5'h0 : _GEN_7579; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_7581 = 5'h16 == _T_715 ? 5'h0 : _GEN_7580; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_7582 = 5'h17 == _T_715 ? w_vn_23 : _GEN_7581; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_7583 = 5'h18 == _T_715 ? w_vn_24 : _GEN_7582; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_7584 = 5'h19 == _T_715 ? 5'h0 : _GEN_7583; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_7585 = 5'h1a == _T_715 ? 5'h0 : _GEN_7584; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_7586 = 5'h1b == _T_715 ? 5'h0 : _GEN_7585; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_7587 = 5'h1c == _T_715 ? 5'h0 : _GEN_7586; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_7588 = 5'h1d == _T_715 ? 5'h0 : _GEN_7587; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_7589 = 5'h1e == _T_715 ? 5'h0 : _GEN_7588; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_7590 = 5'h1f == _T_715 ? 5'h0 : _GEN_7589; // @[FanCtrl.scala 48:{39,39}]
  wire  _T_716 = _GEN_7558 == _GEN_7590; // @[FanCtrl.scala 48:39]
  wire [4:0] _T_726 = _T_710 + 5'h2; // @[FanCtrl.scala 55:32]
  wire [4:0] _GEN_7719 = 5'h3 == _T_726 ? w_vn_3 : 5'h0; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_7720 = 5'h4 == _T_726 ? w_vn_4 : _GEN_7719; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_7721 = 5'h5 == _T_726 ? 5'h0 : _GEN_7720; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_7722 = 5'h6 == _T_726 ? 5'h0 : _GEN_7721; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_7723 = 5'h7 == _T_726 ? w_vn_7 : _GEN_7722; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_7724 = 5'h8 == _T_726 ? w_vn_8 : _GEN_7723; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_7725 = 5'h9 == _T_726 ? 5'h0 : _GEN_7724; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_7726 = 5'ha == _T_726 ? 5'h0 : _GEN_7725; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_7727 = 5'hb == _T_726 ? w_vn_11 : _GEN_7726; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_7728 = 5'hc == _T_726 ? w_vn_12 : _GEN_7727; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_7729 = 5'hd == _T_726 ? w_vn_13 : _GEN_7728; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_7730 = 5'he == _T_726 ? 5'h0 : _GEN_7729; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_7731 = 5'hf == _T_726 ? w_vn_15 : _GEN_7730; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_7732 = 5'h10 == _T_726 ? w_vn_16 : _GEN_7731; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_7733 = 5'h11 == _T_726 ? 5'h0 : _GEN_7732; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_7734 = 5'h12 == _T_726 ? w_vn_18 : _GEN_7733; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_7735 = 5'h13 == _T_726 ? 5'h0 : _GEN_7734; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_7736 = 5'h14 == _T_726 ? 5'h0 : _GEN_7735; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_7737 = 5'h15 == _T_726 ? 5'h0 : _GEN_7736; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_7738 = 5'h16 == _T_726 ? 5'h0 : _GEN_7737; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_7739 = 5'h17 == _T_726 ? w_vn_23 : _GEN_7738; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_7740 = 5'h18 == _T_726 ? w_vn_24 : _GEN_7739; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_7741 = 5'h19 == _T_726 ? 5'h0 : _GEN_7740; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_7742 = 5'h1a == _T_726 ? 5'h0 : _GEN_7741; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_7743 = 5'h1b == _T_726 ? 5'h0 : _GEN_7742; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_7744 = 5'h1c == _T_726 ? 5'h0 : _GEN_7743; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_7745 = 5'h1d == _T_726 ? 5'h0 : _GEN_7744; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_7746 = 5'h1e == _T_726 ? 5'h0 : _GEN_7745; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_7747 = 5'h1f == _T_726 ? 5'h0 : _GEN_7746; // @[FanCtrl.scala 54:{41,41}]
  wire  _T_727 = _GEN_7590 != _GEN_7747; // @[FanCtrl.scala 54:41]
  wire  _T_734 = _GEN_7558 != _GEN_7590; // @[FanCtrl.scala 56:41]
  wire  _T_742 = _GEN_7590 == _GEN_7747; // @[FanCtrl.scala 61:48]
  wire  _GEN_7977 = r_valid_1 & _T_716; // @[FanCtrl.scala 47:34]
  wire [4:0] _T_773 = _T_710 - 5'h1; // @[FanCtrl.scala 94:58]
  wire [4:0] _GEN_8228 = 5'h3 == _T_773 ? w_vn_3 : 5'h0; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_8229 = 5'h4 == _T_773 ? w_vn_4 : _GEN_8228; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_8230 = 5'h5 == _T_773 ? 5'h0 : _GEN_8229; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_8231 = 5'h6 == _T_773 ? 5'h0 : _GEN_8230; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_8232 = 5'h7 == _T_773 ? w_vn_7 : _GEN_8231; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_8233 = 5'h8 == _T_773 ? w_vn_8 : _GEN_8232; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_8234 = 5'h9 == _T_773 ? 5'h0 : _GEN_8233; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_8235 = 5'ha == _T_773 ? 5'h0 : _GEN_8234; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_8236 = 5'hb == _T_773 ? w_vn_11 : _GEN_8235; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_8237 = 5'hc == _T_773 ? w_vn_12 : _GEN_8236; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_8238 = 5'hd == _T_773 ? w_vn_13 : _GEN_8237; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_8239 = 5'he == _T_773 ? 5'h0 : _GEN_8238; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_8240 = 5'hf == _T_773 ? w_vn_15 : _GEN_8239; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_8241 = 5'h10 == _T_773 ? w_vn_16 : _GEN_8240; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_8242 = 5'h11 == _T_773 ? 5'h0 : _GEN_8241; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_8243 = 5'h12 == _T_773 ? w_vn_18 : _GEN_8242; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_8244 = 5'h13 == _T_773 ? 5'h0 : _GEN_8243; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_8245 = 5'h14 == _T_773 ? 5'h0 : _GEN_8244; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_8246 = 5'h15 == _T_773 ? 5'h0 : _GEN_8245; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_8247 = 5'h16 == _T_773 ? 5'h0 : _GEN_8246; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_8248 = 5'h17 == _T_773 ? w_vn_23 : _GEN_8247; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_8249 = 5'h18 == _T_773 ? w_vn_24 : _GEN_8248; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_8250 = 5'h19 == _T_773 ? 5'h0 : _GEN_8249; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_8251 = 5'h1a == _T_773 ? 5'h0 : _GEN_8250; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_8252 = 5'h1b == _T_773 ? 5'h0 : _GEN_8251; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_8253 = 5'h1c == _T_773 ? 5'h0 : _GEN_8252; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_8254 = 5'h1d == _T_773 ? 5'h0 : _GEN_8253; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_8255 = 5'h1e == _T_773 ? 5'h0 : _GEN_8254; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_8256 = 5'h1f == _T_773 ? 5'h0 : _GEN_8255; // @[FanCtrl.scala 94:{39,39}]
  wire  _T_774 = _GEN_7558 != _GEN_8256; // @[FanCtrl.scala 94:39]
  wire  _T_789 = _GEN_7558 == _GEN_8256; // @[FanCtrl.scala 99:46]
  wire  _T_828 = _T_774 & _T_727; // @[FanCtrl.scala 125:65]
  wire  _T_836 = _T_828 & _T_734; // @[FanCtrl.scala 126:65]
  wire  _T_851 = _T_789 & _T_727; // @[FanCtrl.scala 131:70]
  wire  _T_859 = _T_851 & _T_734; // @[FanCtrl.scala 132:72]
  wire  _T_874 = _T_774 & _T_742; // @[FanCtrl.scala 137:72]
  wire  _T_882 = _T_874 & _T_734; // @[FanCtrl.scala 138:71]
  wire [1:0] _GEN_9278 = _T_882 ? 2'h3 : 2'h1; // @[FanCtrl.scala 139:73 141:34 144:35]
  wire [2:0] _GEN_9279 = _T_859 ? 3'h4 : {{1'd0}, _GEN_9278}; // @[FanCtrl.scala 133:73 135:35]
  wire [2:0] _GEN_9280 = _T_836 ? 3'h5 : _GEN_9279; // @[FanCtrl.scala 127:66 129:35]
  wire [2:0] _GEN_9343 = r_valid_1 ? _GEN_9280 : 3'h0; // @[FanCtrl.scala 117:32 148:33]
  wire [4:0] _T_887 = 2'h2 * 3'h5; // @[FanCtrl.scala 48:25]
  wire [5:0] _T_888 = {{1'd0}, _T_887}; // @[FanCtrl.scala 48:31]
  wire [4:0] _T_892 = _T_887 + 5'h1; // @[FanCtrl.scala 48:58]
  wire [4:0] _GEN_9412 = 5'h3 == _T_888[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_9413 = 5'h4 == _T_888[4:0] ? w_vn_4 : _GEN_9412; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_9414 = 5'h5 == _T_888[4:0] ? 5'h0 : _GEN_9413; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_9415 = 5'h6 == _T_888[4:0] ? 5'h0 : _GEN_9414; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_9416 = 5'h7 == _T_888[4:0] ? w_vn_7 : _GEN_9415; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_9417 = 5'h8 == _T_888[4:0] ? w_vn_8 : _GEN_9416; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_9418 = 5'h9 == _T_888[4:0] ? 5'h0 : _GEN_9417; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_9419 = 5'ha == _T_888[4:0] ? 5'h0 : _GEN_9418; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_9420 = 5'hb == _T_888[4:0] ? w_vn_11 : _GEN_9419; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_9421 = 5'hc == _T_888[4:0] ? w_vn_12 : _GEN_9420; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_9422 = 5'hd == _T_888[4:0] ? w_vn_13 : _GEN_9421; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_9423 = 5'he == _T_888[4:0] ? 5'h0 : _GEN_9422; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_9424 = 5'hf == _T_888[4:0] ? w_vn_15 : _GEN_9423; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_9425 = 5'h10 == _T_888[4:0] ? w_vn_16 : _GEN_9424; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_9426 = 5'h11 == _T_888[4:0] ? 5'h0 : _GEN_9425; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_9427 = 5'h12 == _T_888[4:0] ? w_vn_18 : _GEN_9426; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_9428 = 5'h13 == _T_888[4:0] ? 5'h0 : _GEN_9427; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_9429 = 5'h14 == _T_888[4:0] ? 5'h0 : _GEN_9428; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_9430 = 5'h15 == _T_888[4:0] ? 5'h0 : _GEN_9429; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_9431 = 5'h16 == _T_888[4:0] ? 5'h0 : _GEN_9430; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_9432 = 5'h17 == _T_888[4:0] ? w_vn_23 : _GEN_9431; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_9433 = 5'h18 == _T_888[4:0] ? w_vn_24 : _GEN_9432; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_9434 = 5'h19 == _T_888[4:0] ? 5'h0 : _GEN_9433; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_9435 = 5'h1a == _T_888[4:0] ? 5'h0 : _GEN_9434; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_9436 = 5'h1b == _T_888[4:0] ? 5'h0 : _GEN_9435; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_9437 = 5'h1c == _T_888[4:0] ? 5'h0 : _GEN_9436; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_9438 = 5'h1d == _T_888[4:0] ? 5'h0 : _GEN_9437; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_9439 = 5'h1e == _T_888[4:0] ? 5'h0 : _GEN_9438; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_9440 = 5'h1f == _T_888[4:0] ? 5'h0 : _GEN_9439; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_9444 = 5'h3 == _T_892 ? w_vn_3 : 5'h0; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_9445 = 5'h4 == _T_892 ? w_vn_4 : _GEN_9444; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_9446 = 5'h5 == _T_892 ? 5'h0 : _GEN_9445; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_9447 = 5'h6 == _T_892 ? 5'h0 : _GEN_9446; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_9448 = 5'h7 == _T_892 ? w_vn_7 : _GEN_9447; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_9449 = 5'h8 == _T_892 ? w_vn_8 : _GEN_9448; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_9450 = 5'h9 == _T_892 ? 5'h0 : _GEN_9449; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_9451 = 5'ha == _T_892 ? 5'h0 : _GEN_9450; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_9452 = 5'hb == _T_892 ? w_vn_11 : _GEN_9451; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_9453 = 5'hc == _T_892 ? w_vn_12 : _GEN_9452; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_9454 = 5'hd == _T_892 ? w_vn_13 : _GEN_9453; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_9455 = 5'he == _T_892 ? 5'h0 : _GEN_9454; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_9456 = 5'hf == _T_892 ? w_vn_15 : _GEN_9455; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_9457 = 5'h10 == _T_892 ? w_vn_16 : _GEN_9456; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_9458 = 5'h11 == _T_892 ? 5'h0 : _GEN_9457; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_9459 = 5'h12 == _T_892 ? w_vn_18 : _GEN_9458; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_9460 = 5'h13 == _T_892 ? 5'h0 : _GEN_9459; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_9461 = 5'h14 == _T_892 ? 5'h0 : _GEN_9460; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_9462 = 5'h15 == _T_892 ? 5'h0 : _GEN_9461; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_9463 = 5'h16 == _T_892 ? 5'h0 : _GEN_9462; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_9464 = 5'h17 == _T_892 ? w_vn_23 : _GEN_9463; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_9465 = 5'h18 == _T_892 ? w_vn_24 : _GEN_9464; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_9466 = 5'h19 == _T_892 ? 5'h0 : _GEN_9465; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_9467 = 5'h1a == _T_892 ? 5'h0 : _GEN_9466; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_9468 = 5'h1b == _T_892 ? 5'h0 : _GEN_9467; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_9469 = 5'h1c == _T_892 ? 5'h0 : _GEN_9468; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_9470 = 5'h1d == _T_892 ? 5'h0 : _GEN_9469; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_9471 = 5'h1e == _T_892 ? 5'h0 : _GEN_9470; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_9472 = 5'h1f == _T_892 ? 5'h0 : _GEN_9471; // @[FanCtrl.scala 48:{39,39}]
  wire  _T_893 = _GEN_9440 == _GEN_9472; // @[FanCtrl.scala 48:39]
  wire [4:0] _T_903 = _T_887 + 5'h2; // @[FanCtrl.scala 55:32]
  wire [4:0] _GEN_9601 = 5'h3 == _T_903 ? w_vn_3 : 5'h0; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_9602 = 5'h4 == _T_903 ? w_vn_4 : _GEN_9601; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_9603 = 5'h5 == _T_903 ? 5'h0 : _GEN_9602; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_9604 = 5'h6 == _T_903 ? 5'h0 : _GEN_9603; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_9605 = 5'h7 == _T_903 ? w_vn_7 : _GEN_9604; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_9606 = 5'h8 == _T_903 ? w_vn_8 : _GEN_9605; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_9607 = 5'h9 == _T_903 ? 5'h0 : _GEN_9606; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_9608 = 5'ha == _T_903 ? 5'h0 : _GEN_9607; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_9609 = 5'hb == _T_903 ? w_vn_11 : _GEN_9608; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_9610 = 5'hc == _T_903 ? w_vn_12 : _GEN_9609; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_9611 = 5'hd == _T_903 ? w_vn_13 : _GEN_9610; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_9612 = 5'he == _T_903 ? 5'h0 : _GEN_9611; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_9613 = 5'hf == _T_903 ? w_vn_15 : _GEN_9612; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_9614 = 5'h10 == _T_903 ? w_vn_16 : _GEN_9613; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_9615 = 5'h11 == _T_903 ? 5'h0 : _GEN_9614; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_9616 = 5'h12 == _T_903 ? w_vn_18 : _GEN_9615; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_9617 = 5'h13 == _T_903 ? 5'h0 : _GEN_9616; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_9618 = 5'h14 == _T_903 ? 5'h0 : _GEN_9617; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_9619 = 5'h15 == _T_903 ? 5'h0 : _GEN_9618; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_9620 = 5'h16 == _T_903 ? 5'h0 : _GEN_9619; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_9621 = 5'h17 == _T_903 ? w_vn_23 : _GEN_9620; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_9622 = 5'h18 == _T_903 ? w_vn_24 : _GEN_9621; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_9623 = 5'h19 == _T_903 ? 5'h0 : _GEN_9622; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_9624 = 5'h1a == _T_903 ? 5'h0 : _GEN_9623; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_9625 = 5'h1b == _T_903 ? 5'h0 : _GEN_9624; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_9626 = 5'h1c == _T_903 ? 5'h0 : _GEN_9625; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_9627 = 5'h1d == _T_903 ? 5'h0 : _GEN_9626; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_9628 = 5'h1e == _T_903 ? 5'h0 : _GEN_9627; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_9629 = 5'h1f == _T_903 ? 5'h0 : _GEN_9628; // @[FanCtrl.scala 54:{41,41}]
  wire  _T_904 = _GEN_9472 != _GEN_9629; // @[FanCtrl.scala 54:41]
  wire  _T_911 = _GEN_9440 != _GEN_9472; // @[FanCtrl.scala 56:41]
  wire  _T_919 = _GEN_9472 == _GEN_9629; // @[FanCtrl.scala 61:48]
  wire  _GEN_9860 = r_valid_1 & _T_893; // @[FanCtrl.scala 47:34]
  wire [4:0] _T_950 = _T_887 - 5'h1; // @[FanCtrl.scala 94:58]
  wire [4:0] _GEN_10110 = 5'h3 == _T_950 ? w_vn_3 : 5'h0; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_10111 = 5'h4 == _T_950 ? w_vn_4 : _GEN_10110; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_10112 = 5'h5 == _T_950 ? 5'h0 : _GEN_10111; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_10113 = 5'h6 == _T_950 ? 5'h0 : _GEN_10112; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_10114 = 5'h7 == _T_950 ? w_vn_7 : _GEN_10113; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_10115 = 5'h8 == _T_950 ? w_vn_8 : _GEN_10114; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_10116 = 5'h9 == _T_950 ? 5'h0 : _GEN_10115; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_10117 = 5'ha == _T_950 ? 5'h0 : _GEN_10116; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_10118 = 5'hb == _T_950 ? w_vn_11 : _GEN_10117; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_10119 = 5'hc == _T_950 ? w_vn_12 : _GEN_10118; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_10120 = 5'hd == _T_950 ? w_vn_13 : _GEN_10119; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_10121 = 5'he == _T_950 ? 5'h0 : _GEN_10120; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_10122 = 5'hf == _T_950 ? w_vn_15 : _GEN_10121; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_10123 = 5'h10 == _T_950 ? w_vn_16 : _GEN_10122; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_10124 = 5'h11 == _T_950 ? 5'h0 : _GEN_10123; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_10125 = 5'h12 == _T_950 ? w_vn_18 : _GEN_10124; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_10126 = 5'h13 == _T_950 ? 5'h0 : _GEN_10125; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_10127 = 5'h14 == _T_950 ? 5'h0 : _GEN_10126; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_10128 = 5'h15 == _T_950 ? 5'h0 : _GEN_10127; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_10129 = 5'h16 == _T_950 ? 5'h0 : _GEN_10128; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_10130 = 5'h17 == _T_950 ? w_vn_23 : _GEN_10129; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_10131 = 5'h18 == _T_950 ? w_vn_24 : _GEN_10130; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_10132 = 5'h19 == _T_950 ? 5'h0 : _GEN_10131; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_10133 = 5'h1a == _T_950 ? 5'h0 : _GEN_10132; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_10134 = 5'h1b == _T_950 ? 5'h0 : _GEN_10133; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_10135 = 5'h1c == _T_950 ? 5'h0 : _GEN_10134; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_10136 = 5'h1d == _T_950 ? 5'h0 : _GEN_10135; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_10137 = 5'h1e == _T_950 ? 5'h0 : _GEN_10136; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_10138 = 5'h1f == _T_950 ? 5'h0 : _GEN_10137; // @[FanCtrl.scala 94:{39,39}]
  wire  _T_951 = _GEN_9440 != _GEN_10138; // @[FanCtrl.scala 94:39]
  wire  _T_966 = _GEN_9440 == _GEN_10138; // @[FanCtrl.scala 99:46]
  wire  _T_1005 = _T_951 & _T_904; // @[FanCtrl.scala 125:65]
  wire  _T_1013 = _T_1005 & _T_911; // @[FanCtrl.scala 126:65]
  wire  _T_1028 = _T_966 & _T_904; // @[FanCtrl.scala 131:70]
  wire  _T_1036 = _T_1028 & _T_911; // @[FanCtrl.scala 132:72]
  wire  _T_1051 = _T_951 & _T_919; // @[FanCtrl.scala 137:72]
  wire  _T_1059 = _T_1051 & _T_911; // @[FanCtrl.scala 138:71]
  wire [1:0] _GEN_11160 = _T_1059 ? 2'h3 : 2'h1; // @[FanCtrl.scala 139:73 141:34 144:35]
  wire [2:0] _GEN_11161 = _T_1036 ? 3'h4 : {{1'd0}, _GEN_11160}; // @[FanCtrl.scala 133:73 135:35]
  wire [2:0] _GEN_11162 = _T_1013 ? 3'h5 : _GEN_11161; // @[FanCtrl.scala 127:66 129:35]
  wire [2:0] _GEN_11225 = r_valid_1 ? _GEN_11162 : 3'h0; // @[FanCtrl.scala 117:32 148:33]
  wire [4:0] _T_1064 = 2'h2 * 3'h6; // @[FanCtrl.scala 48:25]
  wire [5:0] _T_1065 = {{1'd0}, _T_1064}; // @[FanCtrl.scala 48:31]
  wire [4:0] _T_1069 = _T_1064 + 5'h1; // @[FanCtrl.scala 48:58]
  wire [4:0] _GEN_11294 = 5'h3 == _T_1065[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_11295 = 5'h4 == _T_1065[4:0] ? w_vn_4 : _GEN_11294; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_11296 = 5'h5 == _T_1065[4:0] ? 5'h0 : _GEN_11295; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_11297 = 5'h6 == _T_1065[4:0] ? 5'h0 : _GEN_11296; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_11298 = 5'h7 == _T_1065[4:0] ? w_vn_7 : _GEN_11297; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_11299 = 5'h8 == _T_1065[4:0] ? w_vn_8 : _GEN_11298; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_11300 = 5'h9 == _T_1065[4:0] ? 5'h0 : _GEN_11299; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_11301 = 5'ha == _T_1065[4:0] ? 5'h0 : _GEN_11300; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_11302 = 5'hb == _T_1065[4:0] ? w_vn_11 : _GEN_11301; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_11303 = 5'hc == _T_1065[4:0] ? w_vn_12 : _GEN_11302; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_11304 = 5'hd == _T_1065[4:0] ? w_vn_13 : _GEN_11303; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_11305 = 5'he == _T_1065[4:0] ? 5'h0 : _GEN_11304; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_11306 = 5'hf == _T_1065[4:0] ? w_vn_15 : _GEN_11305; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_11307 = 5'h10 == _T_1065[4:0] ? w_vn_16 : _GEN_11306; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_11308 = 5'h11 == _T_1065[4:0] ? 5'h0 : _GEN_11307; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_11309 = 5'h12 == _T_1065[4:0] ? w_vn_18 : _GEN_11308; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_11310 = 5'h13 == _T_1065[4:0] ? 5'h0 : _GEN_11309; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_11311 = 5'h14 == _T_1065[4:0] ? 5'h0 : _GEN_11310; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_11312 = 5'h15 == _T_1065[4:0] ? 5'h0 : _GEN_11311; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_11313 = 5'h16 == _T_1065[4:0] ? 5'h0 : _GEN_11312; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_11314 = 5'h17 == _T_1065[4:0] ? w_vn_23 : _GEN_11313; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_11315 = 5'h18 == _T_1065[4:0] ? w_vn_24 : _GEN_11314; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_11316 = 5'h19 == _T_1065[4:0] ? 5'h0 : _GEN_11315; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_11317 = 5'h1a == _T_1065[4:0] ? 5'h0 : _GEN_11316; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_11318 = 5'h1b == _T_1065[4:0] ? 5'h0 : _GEN_11317; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_11319 = 5'h1c == _T_1065[4:0] ? 5'h0 : _GEN_11318; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_11320 = 5'h1d == _T_1065[4:0] ? 5'h0 : _GEN_11319; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_11321 = 5'h1e == _T_1065[4:0] ? 5'h0 : _GEN_11320; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_11322 = 5'h1f == _T_1065[4:0] ? 5'h0 : _GEN_11321; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_11326 = 5'h3 == _T_1069 ? w_vn_3 : 5'h0; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_11327 = 5'h4 == _T_1069 ? w_vn_4 : _GEN_11326; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_11328 = 5'h5 == _T_1069 ? 5'h0 : _GEN_11327; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_11329 = 5'h6 == _T_1069 ? 5'h0 : _GEN_11328; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_11330 = 5'h7 == _T_1069 ? w_vn_7 : _GEN_11329; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_11331 = 5'h8 == _T_1069 ? w_vn_8 : _GEN_11330; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_11332 = 5'h9 == _T_1069 ? 5'h0 : _GEN_11331; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_11333 = 5'ha == _T_1069 ? 5'h0 : _GEN_11332; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_11334 = 5'hb == _T_1069 ? w_vn_11 : _GEN_11333; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_11335 = 5'hc == _T_1069 ? w_vn_12 : _GEN_11334; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_11336 = 5'hd == _T_1069 ? w_vn_13 : _GEN_11335; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_11337 = 5'he == _T_1069 ? 5'h0 : _GEN_11336; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_11338 = 5'hf == _T_1069 ? w_vn_15 : _GEN_11337; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_11339 = 5'h10 == _T_1069 ? w_vn_16 : _GEN_11338; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_11340 = 5'h11 == _T_1069 ? 5'h0 : _GEN_11339; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_11341 = 5'h12 == _T_1069 ? w_vn_18 : _GEN_11340; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_11342 = 5'h13 == _T_1069 ? 5'h0 : _GEN_11341; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_11343 = 5'h14 == _T_1069 ? 5'h0 : _GEN_11342; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_11344 = 5'h15 == _T_1069 ? 5'h0 : _GEN_11343; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_11345 = 5'h16 == _T_1069 ? 5'h0 : _GEN_11344; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_11346 = 5'h17 == _T_1069 ? w_vn_23 : _GEN_11345; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_11347 = 5'h18 == _T_1069 ? w_vn_24 : _GEN_11346; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_11348 = 5'h19 == _T_1069 ? 5'h0 : _GEN_11347; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_11349 = 5'h1a == _T_1069 ? 5'h0 : _GEN_11348; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_11350 = 5'h1b == _T_1069 ? 5'h0 : _GEN_11349; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_11351 = 5'h1c == _T_1069 ? 5'h0 : _GEN_11350; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_11352 = 5'h1d == _T_1069 ? 5'h0 : _GEN_11351; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_11353 = 5'h1e == _T_1069 ? 5'h0 : _GEN_11352; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_11354 = 5'h1f == _T_1069 ? 5'h0 : _GEN_11353; // @[FanCtrl.scala 48:{39,39}]
  wire  _T_1070 = _GEN_11322 == _GEN_11354; // @[FanCtrl.scala 48:39]
  wire [4:0] _T_1080 = _T_1064 + 5'h2; // @[FanCtrl.scala 55:32]
  wire [4:0] _GEN_11483 = 5'h3 == _T_1080 ? w_vn_3 : 5'h0; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_11484 = 5'h4 == _T_1080 ? w_vn_4 : _GEN_11483; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_11485 = 5'h5 == _T_1080 ? 5'h0 : _GEN_11484; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_11486 = 5'h6 == _T_1080 ? 5'h0 : _GEN_11485; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_11487 = 5'h7 == _T_1080 ? w_vn_7 : _GEN_11486; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_11488 = 5'h8 == _T_1080 ? w_vn_8 : _GEN_11487; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_11489 = 5'h9 == _T_1080 ? 5'h0 : _GEN_11488; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_11490 = 5'ha == _T_1080 ? 5'h0 : _GEN_11489; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_11491 = 5'hb == _T_1080 ? w_vn_11 : _GEN_11490; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_11492 = 5'hc == _T_1080 ? w_vn_12 : _GEN_11491; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_11493 = 5'hd == _T_1080 ? w_vn_13 : _GEN_11492; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_11494 = 5'he == _T_1080 ? 5'h0 : _GEN_11493; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_11495 = 5'hf == _T_1080 ? w_vn_15 : _GEN_11494; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_11496 = 5'h10 == _T_1080 ? w_vn_16 : _GEN_11495; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_11497 = 5'h11 == _T_1080 ? 5'h0 : _GEN_11496; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_11498 = 5'h12 == _T_1080 ? w_vn_18 : _GEN_11497; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_11499 = 5'h13 == _T_1080 ? 5'h0 : _GEN_11498; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_11500 = 5'h14 == _T_1080 ? 5'h0 : _GEN_11499; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_11501 = 5'h15 == _T_1080 ? 5'h0 : _GEN_11500; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_11502 = 5'h16 == _T_1080 ? 5'h0 : _GEN_11501; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_11503 = 5'h17 == _T_1080 ? w_vn_23 : _GEN_11502; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_11504 = 5'h18 == _T_1080 ? w_vn_24 : _GEN_11503; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_11505 = 5'h19 == _T_1080 ? 5'h0 : _GEN_11504; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_11506 = 5'h1a == _T_1080 ? 5'h0 : _GEN_11505; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_11507 = 5'h1b == _T_1080 ? 5'h0 : _GEN_11506; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_11508 = 5'h1c == _T_1080 ? 5'h0 : _GEN_11507; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_11509 = 5'h1d == _T_1080 ? 5'h0 : _GEN_11508; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_11510 = 5'h1e == _T_1080 ? 5'h0 : _GEN_11509; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_11511 = 5'h1f == _T_1080 ? 5'h0 : _GEN_11510; // @[FanCtrl.scala 54:{41,41}]
  wire  _T_1081 = _GEN_11354 != _GEN_11511; // @[FanCtrl.scala 54:41]
  wire  _T_1088 = _GEN_11322 != _GEN_11354; // @[FanCtrl.scala 56:41]
  wire  _T_1096 = _GEN_11354 == _GEN_11511; // @[FanCtrl.scala 61:48]
  wire  _GEN_11743 = r_valid_1 & _T_1070; // @[FanCtrl.scala 47:34]
  wire [4:0] _T_1127 = _T_1064 - 5'h1; // @[FanCtrl.scala 94:58]
  wire [4:0] _GEN_11992 = 5'h3 == _T_1127 ? w_vn_3 : 5'h0; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_11993 = 5'h4 == _T_1127 ? w_vn_4 : _GEN_11992; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_11994 = 5'h5 == _T_1127 ? 5'h0 : _GEN_11993; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_11995 = 5'h6 == _T_1127 ? 5'h0 : _GEN_11994; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_11996 = 5'h7 == _T_1127 ? w_vn_7 : _GEN_11995; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_11997 = 5'h8 == _T_1127 ? w_vn_8 : _GEN_11996; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_11998 = 5'h9 == _T_1127 ? 5'h0 : _GEN_11997; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_11999 = 5'ha == _T_1127 ? 5'h0 : _GEN_11998; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_12000 = 5'hb == _T_1127 ? w_vn_11 : _GEN_11999; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_12001 = 5'hc == _T_1127 ? w_vn_12 : _GEN_12000; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_12002 = 5'hd == _T_1127 ? w_vn_13 : _GEN_12001; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_12003 = 5'he == _T_1127 ? 5'h0 : _GEN_12002; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_12004 = 5'hf == _T_1127 ? w_vn_15 : _GEN_12003; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_12005 = 5'h10 == _T_1127 ? w_vn_16 : _GEN_12004; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_12006 = 5'h11 == _T_1127 ? 5'h0 : _GEN_12005; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_12007 = 5'h12 == _T_1127 ? w_vn_18 : _GEN_12006; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_12008 = 5'h13 == _T_1127 ? 5'h0 : _GEN_12007; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_12009 = 5'h14 == _T_1127 ? 5'h0 : _GEN_12008; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_12010 = 5'h15 == _T_1127 ? 5'h0 : _GEN_12009; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_12011 = 5'h16 == _T_1127 ? 5'h0 : _GEN_12010; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_12012 = 5'h17 == _T_1127 ? w_vn_23 : _GEN_12011; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_12013 = 5'h18 == _T_1127 ? w_vn_24 : _GEN_12012; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_12014 = 5'h19 == _T_1127 ? 5'h0 : _GEN_12013; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_12015 = 5'h1a == _T_1127 ? 5'h0 : _GEN_12014; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_12016 = 5'h1b == _T_1127 ? 5'h0 : _GEN_12015; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_12017 = 5'h1c == _T_1127 ? 5'h0 : _GEN_12016; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_12018 = 5'h1d == _T_1127 ? 5'h0 : _GEN_12017; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_12019 = 5'h1e == _T_1127 ? 5'h0 : _GEN_12018; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_12020 = 5'h1f == _T_1127 ? 5'h0 : _GEN_12019; // @[FanCtrl.scala 94:{39,39}]
  wire  _T_1128 = _GEN_11322 != _GEN_12020; // @[FanCtrl.scala 94:39]
  wire  _T_1143 = _GEN_11322 == _GEN_12020; // @[FanCtrl.scala 99:46]
  wire  _T_1182 = _T_1128 & _T_1081; // @[FanCtrl.scala 125:65]
  wire  _T_1190 = _T_1182 & _T_1088; // @[FanCtrl.scala 126:65]
  wire  _T_1205 = _T_1143 & _T_1081; // @[FanCtrl.scala 131:70]
  wire  _T_1213 = _T_1205 & _T_1088; // @[FanCtrl.scala 132:72]
  wire  _T_1228 = _T_1128 & _T_1096; // @[FanCtrl.scala 137:72]
  wire  _T_1236 = _T_1228 & _T_1088; // @[FanCtrl.scala 138:71]
  wire [1:0] _GEN_13042 = _T_1236 ? 2'h3 : 2'h1; // @[FanCtrl.scala 139:73 141:34 144:35]
  wire [2:0] _GEN_13043 = _T_1213 ? 3'h4 : {{1'd0}, _GEN_13042}; // @[FanCtrl.scala 133:73 135:35]
  wire [2:0] _GEN_13044 = _T_1190 ? 3'h5 : _GEN_13043; // @[FanCtrl.scala 127:66 129:35]
  wire [2:0] _GEN_13107 = r_valid_1 ? _GEN_13044 : 3'h0; // @[FanCtrl.scala 117:32 148:33]
  wire [4:0] _T_1241 = 2'h2 * 3'h7; // @[FanCtrl.scala 48:25]
  wire [5:0] _T_1242 = {{1'd0}, _T_1241}; // @[FanCtrl.scala 48:31]
  wire [4:0] _T_1246 = _T_1241 + 5'h1; // @[FanCtrl.scala 48:58]
  wire [4:0] _GEN_13176 = 5'h3 == _T_1242[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_13177 = 5'h4 == _T_1242[4:0] ? w_vn_4 : _GEN_13176; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_13178 = 5'h5 == _T_1242[4:0] ? 5'h0 : _GEN_13177; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_13179 = 5'h6 == _T_1242[4:0] ? 5'h0 : _GEN_13178; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_13180 = 5'h7 == _T_1242[4:0] ? w_vn_7 : _GEN_13179; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_13181 = 5'h8 == _T_1242[4:0] ? w_vn_8 : _GEN_13180; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_13182 = 5'h9 == _T_1242[4:0] ? 5'h0 : _GEN_13181; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_13183 = 5'ha == _T_1242[4:0] ? 5'h0 : _GEN_13182; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_13184 = 5'hb == _T_1242[4:0] ? w_vn_11 : _GEN_13183; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_13185 = 5'hc == _T_1242[4:0] ? w_vn_12 : _GEN_13184; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_13186 = 5'hd == _T_1242[4:0] ? w_vn_13 : _GEN_13185; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_13187 = 5'he == _T_1242[4:0] ? 5'h0 : _GEN_13186; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_13188 = 5'hf == _T_1242[4:0] ? w_vn_15 : _GEN_13187; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_13189 = 5'h10 == _T_1242[4:0] ? w_vn_16 : _GEN_13188; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_13190 = 5'h11 == _T_1242[4:0] ? 5'h0 : _GEN_13189; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_13191 = 5'h12 == _T_1242[4:0] ? w_vn_18 : _GEN_13190; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_13192 = 5'h13 == _T_1242[4:0] ? 5'h0 : _GEN_13191; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_13193 = 5'h14 == _T_1242[4:0] ? 5'h0 : _GEN_13192; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_13194 = 5'h15 == _T_1242[4:0] ? 5'h0 : _GEN_13193; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_13195 = 5'h16 == _T_1242[4:0] ? 5'h0 : _GEN_13194; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_13196 = 5'h17 == _T_1242[4:0] ? w_vn_23 : _GEN_13195; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_13197 = 5'h18 == _T_1242[4:0] ? w_vn_24 : _GEN_13196; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_13198 = 5'h19 == _T_1242[4:0] ? 5'h0 : _GEN_13197; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_13199 = 5'h1a == _T_1242[4:0] ? 5'h0 : _GEN_13198; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_13200 = 5'h1b == _T_1242[4:0] ? 5'h0 : _GEN_13199; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_13201 = 5'h1c == _T_1242[4:0] ? 5'h0 : _GEN_13200; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_13202 = 5'h1d == _T_1242[4:0] ? 5'h0 : _GEN_13201; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_13203 = 5'h1e == _T_1242[4:0] ? 5'h0 : _GEN_13202; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_13204 = 5'h1f == _T_1242[4:0] ? 5'h0 : _GEN_13203; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_13208 = 5'h3 == _T_1246 ? w_vn_3 : 5'h0; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_13209 = 5'h4 == _T_1246 ? w_vn_4 : _GEN_13208; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_13210 = 5'h5 == _T_1246 ? 5'h0 : _GEN_13209; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_13211 = 5'h6 == _T_1246 ? 5'h0 : _GEN_13210; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_13212 = 5'h7 == _T_1246 ? w_vn_7 : _GEN_13211; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_13213 = 5'h8 == _T_1246 ? w_vn_8 : _GEN_13212; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_13214 = 5'h9 == _T_1246 ? 5'h0 : _GEN_13213; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_13215 = 5'ha == _T_1246 ? 5'h0 : _GEN_13214; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_13216 = 5'hb == _T_1246 ? w_vn_11 : _GEN_13215; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_13217 = 5'hc == _T_1246 ? w_vn_12 : _GEN_13216; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_13218 = 5'hd == _T_1246 ? w_vn_13 : _GEN_13217; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_13219 = 5'he == _T_1246 ? 5'h0 : _GEN_13218; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_13220 = 5'hf == _T_1246 ? w_vn_15 : _GEN_13219; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_13221 = 5'h10 == _T_1246 ? w_vn_16 : _GEN_13220; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_13222 = 5'h11 == _T_1246 ? 5'h0 : _GEN_13221; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_13223 = 5'h12 == _T_1246 ? w_vn_18 : _GEN_13222; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_13224 = 5'h13 == _T_1246 ? 5'h0 : _GEN_13223; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_13225 = 5'h14 == _T_1246 ? 5'h0 : _GEN_13224; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_13226 = 5'h15 == _T_1246 ? 5'h0 : _GEN_13225; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_13227 = 5'h16 == _T_1246 ? 5'h0 : _GEN_13226; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_13228 = 5'h17 == _T_1246 ? w_vn_23 : _GEN_13227; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_13229 = 5'h18 == _T_1246 ? w_vn_24 : _GEN_13228; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_13230 = 5'h19 == _T_1246 ? 5'h0 : _GEN_13229; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_13231 = 5'h1a == _T_1246 ? 5'h0 : _GEN_13230; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_13232 = 5'h1b == _T_1246 ? 5'h0 : _GEN_13231; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_13233 = 5'h1c == _T_1246 ? 5'h0 : _GEN_13232; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_13234 = 5'h1d == _T_1246 ? 5'h0 : _GEN_13233; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_13235 = 5'h1e == _T_1246 ? 5'h0 : _GEN_13234; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_13236 = 5'h1f == _T_1246 ? 5'h0 : _GEN_13235; // @[FanCtrl.scala 48:{39,39}]
  wire  _T_1247 = _GEN_13204 == _GEN_13236; // @[FanCtrl.scala 48:39]
  wire [4:0] _T_1257 = _T_1241 + 5'h2; // @[FanCtrl.scala 55:32]
  wire [4:0] _GEN_13365 = 5'h3 == _T_1257 ? w_vn_3 : 5'h0; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_13366 = 5'h4 == _T_1257 ? w_vn_4 : _GEN_13365; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_13367 = 5'h5 == _T_1257 ? 5'h0 : _GEN_13366; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_13368 = 5'h6 == _T_1257 ? 5'h0 : _GEN_13367; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_13369 = 5'h7 == _T_1257 ? w_vn_7 : _GEN_13368; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_13370 = 5'h8 == _T_1257 ? w_vn_8 : _GEN_13369; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_13371 = 5'h9 == _T_1257 ? 5'h0 : _GEN_13370; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_13372 = 5'ha == _T_1257 ? 5'h0 : _GEN_13371; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_13373 = 5'hb == _T_1257 ? w_vn_11 : _GEN_13372; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_13374 = 5'hc == _T_1257 ? w_vn_12 : _GEN_13373; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_13375 = 5'hd == _T_1257 ? w_vn_13 : _GEN_13374; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_13376 = 5'he == _T_1257 ? 5'h0 : _GEN_13375; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_13377 = 5'hf == _T_1257 ? w_vn_15 : _GEN_13376; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_13378 = 5'h10 == _T_1257 ? w_vn_16 : _GEN_13377; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_13379 = 5'h11 == _T_1257 ? 5'h0 : _GEN_13378; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_13380 = 5'h12 == _T_1257 ? w_vn_18 : _GEN_13379; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_13381 = 5'h13 == _T_1257 ? 5'h0 : _GEN_13380; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_13382 = 5'h14 == _T_1257 ? 5'h0 : _GEN_13381; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_13383 = 5'h15 == _T_1257 ? 5'h0 : _GEN_13382; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_13384 = 5'h16 == _T_1257 ? 5'h0 : _GEN_13383; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_13385 = 5'h17 == _T_1257 ? w_vn_23 : _GEN_13384; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_13386 = 5'h18 == _T_1257 ? w_vn_24 : _GEN_13385; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_13387 = 5'h19 == _T_1257 ? 5'h0 : _GEN_13386; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_13388 = 5'h1a == _T_1257 ? 5'h0 : _GEN_13387; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_13389 = 5'h1b == _T_1257 ? 5'h0 : _GEN_13388; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_13390 = 5'h1c == _T_1257 ? 5'h0 : _GEN_13389; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_13391 = 5'h1d == _T_1257 ? 5'h0 : _GEN_13390; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_13392 = 5'h1e == _T_1257 ? 5'h0 : _GEN_13391; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_13393 = 5'h1f == _T_1257 ? 5'h0 : _GEN_13392; // @[FanCtrl.scala 54:{41,41}]
  wire  _T_1258 = _GEN_13236 != _GEN_13393; // @[FanCtrl.scala 54:41]
  wire  _T_1265 = _GEN_13204 != _GEN_13236; // @[FanCtrl.scala 56:41]
  wire  _T_1273 = _GEN_13236 == _GEN_13393; // @[FanCtrl.scala 61:48]
  wire  _GEN_13626 = r_valid_1 & _T_1247; // @[FanCtrl.scala 47:34]
  wire [4:0] _T_1304 = _T_1241 - 5'h1; // @[FanCtrl.scala 94:58]
  wire [4:0] _GEN_13874 = 5'h3 == _T_1304 ? w_vn_3 : 5'h0; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_13875 = 5'h4 == _T_1304 ? w_vn_4 : _GEN_13874; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_13876 = 5'h5 == _T_1304 ? 5'h0 : _GEN_13875; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_13877 = 5'h6 == _T_1304 ? 5'h0 : _GEN_13876; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_13878 = 5'h7 == _T_1304 ? w_vn_7 : _GEN_13877; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_13879 = 5'h8 == _T_1304 ? w_vn_8 : _GEN_13878; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_13880 = 5'h9 == _T_1304 ? 5'h0 : _GEN_13879; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_13881 = 5'ha == _T_1304 ? 5'h0 : _GEN_13880; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_13882 = 5'hb == _T_1304 ? w_vn_11 : _GEN_13881; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_13883 = 5'hc == _T_1304 ? w_vn_12 : _GEN_13882; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_13884 = 5'hd == _T_1304 ? w_vn_13 : _GEN_13883; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_13885 = 5'he == _T_1304 ? 5'h0 : _GEN_13884; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_13886 = 5'hf == _T_1304 ? w_vn_15 : _GEN_13885; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_13887 = 5'h10 == _T_1304 ? w_vn_16 : _GEN_13886; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_13888 = 5'h11 == _T_1304 ? 5'h0 : _GEN_13887; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_13889 = 5'h12 == _T_1304 ? w_vn_18 : _GEN_13888; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_13890 = 5'h13 == _T_1304 ? 5'h0 : _GEN_13889; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_13891 = 5'h14 == _T_1304 ? 5'h0 : _GEN_13890; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_13892 = 5'h15 == _T_1304 ? 5'h0 : _GEN_13891; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_13893 = 5'h16 == _T_1304 ? 5'h0 : _GEN_13892; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_13894 = 5'h17 == _T_1304 ? w_vn_23 : _GEN_13893; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_13895 = 5'h18 == _T_1304 ? w_vn_24 : _GEN_13894; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_13896 = 5'h19 == _T_1304 ? 5'h0 : _GEN_13895; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_13897 = 5'h1a == _T_1304 ? 5'h0 : _GEN_13896; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_13898 = 5'h1b == _T_1304 ? 5'h0 : _GEN_13897; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_13899 = 5'h1c == _T_1304 ? 5'h0 : _GEN_13898; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_13900 = 5'h1d == _T_1304 ? 5'h0 : _GEN_13899; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_13901 = 5'h1e == _T_1304 ? 5'h0 : _GEN_13900; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_13902 = 5'h1f == _T_1304 ? 5'h0 : _GEN_13901; // @[FanCtrl.scala 94:{39,39}]
  wire  _T_1305 = _GEN_13204 != _GEN_13902; // @[FanCtrl.scala 94:39]
  wire  _T_1320 = _GEN_13204 == _GEN_13902; // @[FanCtrl.scala 99:46]
  wire  _T_1359 = _T_1305 & _T_1258; // @[FanCtrl.scala 125:65]
  wire  _T_1367 = _T_1359 & _T_1265; // @[FanCtrl.scala 126:65]
  wire  _T_1382 = _T_1320 & _T_1258; // @[FanCtrl.scala 131:70]
  wire  _T_1390 = _T_1382 & _T_1265; // @[FanCtrl.scala 132:72]
  wire  _T_1405 = _T_1305 & _T_1273; // @[FanCtrl.scala 137:72]
  wire  _T_1413 = _T_1405 & _T_1265; // @[FanCtrl.scala 138:71]
  wire [1:0] _GEN_14924 = _T_1413 ? 2'h3 : 2'h1; // @[FanCtrl.scala 139:73 141:34 144:35]
  wire [2:0] _GEN_14925 = _T_1390 ? 3'h4 : {{1'd0}, _GEN_14924}; // @[FanCtrl.scala 133:73 135:35]
  wire [2:0] _GEN_14926 = _T_1367 ? 3'h5 : _GEN_14925; // @[FanCtrl.scala 127:66 129:35]
  wire [2:0] _GEN_14989 = r_valid_1 ? _GEN_14926 : 3'h0; // @[FanCtrl.scala 117:32 148:33]
  wire [5:0] _T_1418 = 2'h2 * 4'h8; // @[FanCtrl.scala 48:25]
  wire [6:0] _T_1419 = {{1'd0}, _T_1418}; // @[FanCtrl.scala 48:31]
  wire [5:0] _T_1424 = _T_1418 + 6'h1; // @[FanCtrl.scala 48:58]
  wire [4:0] _GEN_15058 = 5'h3 == _T_1419[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_15059 = 5'h4 == _T_1419[4:0] ? w_vn_4 : _GEN_15058; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_15060 = 5'h5 == _T_1419[4:0] ? 5'h0 : _GEN_15059; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_15061 = 5'h6 == _T_1419[4:0] ? 5'h0 : _GEN_15060; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_15062 = 5'h7 == _T_1419[4:0] ? w_vn_7 : _GEN_15061; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_15063 = 5'h8 == _T_1419[4:0] ? w_vn_8 : _GEN_15062; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_15064 = 5'h9 == _T_1419[4:0] ? 5'h0 : _GEN_15063; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_15065 = 5'ha == _T_1419[4:0] ? 5'h0 : _GEN_15064; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_15066 = 5'hb == _T_1419[4:0] ? w_vn_11 : _GEN_15065; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_15067 = 5'hc == _T_1419[4:0] ? w_vn_12 : _GEN_15066; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_15068 = 5'hd == _T_1419[4:0] ? w_vn_13 : _GEN_15067; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_15069 = 5'he == _T_1419[4:0] ? 5'h0 : _GEN_15068; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_15070 = 5'hf == _T_1419[4:0] ? w_vn_15 : _GEN_15069; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_15071 = 5'h10 == _T_1419[4:0] ? w_vn_16 : _GEN_15070; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_15072 = 5'h11 == _T_1419[4:0] ? 5'h0 : _GEN_15071; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_15073 = 5'h12 == _T_1419[4:0] ? w_vn_18 : _GEN_15072; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_15074 = 5'h13 == _T_1419[4:0] ? 5'h0 : _GEN_15073; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_15075 = 5'h14 == _T_1419[4:0] ? 5'h0 : _GEN_15074; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_15076 = 5'h15 == _T_1419[4:0] ? 5'h0 : _GEN_15075; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_15077 = 5'h16 == _T_1419[4:0] ? 5'h0 : _GEN_15076; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_15078 = 5'h17 == _T_1419[4:0] ? w_vn_23 : _GEN_15077; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_15079 = 5'h18 == _T_1419[4:0] ? w_vn_24 : _GEN_15078; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_15080 = 5'h19 == _T_1419[4:0] ? 5'h0 : _GEN_15079; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_15081 = 5'h1a == _T_1419[4:0] ? 5'h0 : _GEN_15080; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_15082 = 5'h1b == _T_1419[4:0] ? 5'h0 : _GEN_15081; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_15083 = 5'h1c == _T_1419[4:0] ? 5'h0 : _GEN_15082; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_15084 = 5'h1d == _T_1419[4:0] ? 5'h0 : _GEN_15083; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_15085 = 5'h1e == _T_1419[4:0] ? 5'h0 : _GEN_15084; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_15086 = 5'h1f == _T_1419[4:0] ? 5'h0 : _GEN_15085; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_15090 = 5'h3 == _T_1424[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_15091 = 5'h4 == _T_1424[4:0] ? w_vn_4 : _GEN_15090; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_15092 = 5'h5 == _T_1424[4:0] ? 5'h0 : _GEN_15091; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_15093 = 5'h6 == _T_1424[4:0] ? 5'h0 : _GEN_15092; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_15094 = 5'h7 == _T_1424[4:0] ? w_vn_7 : _GEN_15093; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_15095 = 5'h8 == _T_1424[4:0] ? w_vn_8 : _GEN_15094; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_15096 = 5'h9 == _T_1424[4:0] ? 5'h0 : _GEN_15095; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_15097 = 5'ha == _T_1424[4:0] ? 5'h0 : _GEN_15096; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_15098 = 5'hb == _T_1424[4:0] ? w_vn_11 : _GEN_15097; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_15099 = 5'hc == _T_1424[4:0] ? w_vn_12 : _GEN_15098; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_15100 = 5'hd == _T_1424[4:0] ? w_vn_13 : _GEN_15099; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_15101 = 5'he == _T_1424[4:0] ? 5'h0 : _GEN_15100; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_15102 = 5'hf == _T_1424[4:0] ? w_vn_15 : _GEN_15101; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_15103 = 5'h10 == _T_1424[4:0] ? w_vn_16 : _GEN_15102; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_15104 = 5'h11 == _T_1424[4:0] ? 5'h0 : _GEN_15103; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_15105 = 5'h12 == _T_1424[4:0] ? w_vn_18 : _GEN_15104; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_15106 = 5'h13 == _T_1424[4:0] ? 5'h0 : _GEN_15105; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_15107 = 5'h14 == _T_1424[4:0] ? 5'h0 : _GEN_15106; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_15108 = 5'h15 == _T_1424[4:0] ? 5'h0 : _GEN_15107; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_15109 = 5'h16 == _T_1424[4:0] ? 5'h0 : _GEN_15108; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_15110 = 5'h17 == _T_1424[4:0] ? w_vn_23 : _GEN_15109; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_15111 = 5'h18 == _T_1424[4:0] ? w_vn_24 : _GEN_15110; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_15112 = 5'h19 == _T_1424[4:0] ? 5'h0 : _GEN_15111; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_15113 = 5'h1a == _T_1424[4:0] ? 5'h0 : _GEN_15112; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_15114 = 5'h1b == _T_1424[4:0] ? 5'h0 : _GEN_15113; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_15115 = 5'h1c == _T_1424[4:0] ? 5'h0 : _GEN_15114; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_15116 = 5'h1d == _T_1424[4:0] ? 5'h0 : _GEN_15115; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_15117 = 5'h1e == _T_1424[4:0] ? 5'h0 : _GEN_15116; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_15118 = 5'h1f == _T_1424[4:0] ? 5'h0 : _GEN_15117; // @[FanCtrl.scala 48:{39,39}]
  wire  _T_1426 = _GEN_15086 == _GEN_15118; // @[FanCtrl.scala 48:39]
  wire [5:0] _T_1437 = _T_1418 + 6'h2; // @[FanCtrl.scala 55:32]
  wire [4:0] _GEN_15247 = 5'h3 == _T_1437[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_15248 = 5'h4 == _T_1437[4:0] ? w_vn_4 : _GEN_15247; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_15249 = 5'h5 == _T_1437[4:0] ? 5'h0 : _GEN_15248; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_15250 = 5'h6 == _T_1437[4:0] ? 5'h0 : _GEN_15249; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_15251 = 5'h7 == _T_1437[4:0] ? w_vn_7 : _GEN_15250; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_15252 = 5'h8 == _T_1437[4:0] ? w_vn_8 : _GEN_15251; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_15253 = 5'h9 == _T_1437[4:0] ? 5'h0 : _GEN_15252; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_15254 = 5'ha == _T_1437[4:0] ? 5'h0 : _GEN_15253; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_15255 = 5'hb == _T_1437[4:0] ? w_vn_11 : _GEN_15254; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_15256 = 5'hc == _T_1437[4:0] ? w_vn_12 : _GEN_15255; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_15257 = 5'hd == _T_1437[4:0] ? w_vn_13 : _GEN_15256; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_15258 = 5'he == _T_1437[4:0] ? 5'h0 : _GEN_15257; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_15259 = 5'hf == _T_1437[4:0] ? w_vn_15 : _GEN_15258; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_15260 = 5'h10 == _T_1437[4:0] ? w_vn_16 : _GEN_15259; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_15261 = 5'h11 == _T_1437[4:0] ? 5'h0 : _GEN_15260; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_15262 = 5'h12 == _T_1437[4:0] ? w_vn_18 : _GEN_15261; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_15263 = 5'h13 == _T_1437[4:0] ? 5'h0 : _GEN_15262; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_15264 = 5'h14 == _T_1437[4:0] ? 5'h0 : _GEN_15263; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_15265 = 5'h15 == _T_1437[4:0] ? 5'h0 : _GEN_15264; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_15266 = 5'h16 == _T_1437[4:0] ? 5'h0 : _GEN_15265; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_15267 = 5'h17 == _T_1437[4:0] ? w_vn_23 : _GEN_15266; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_15268 = 5'h18 == _T_1437[4:0] ? w_vn_24 : _GEN_15267; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_15269 = 5'h19 == _T_1437[4:0] ? 5'h0 : _GEN_15268; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_15270 = 5'h1a == _T_1437[4:0] ? 5'h0 : _GEN_15269; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_15271 = 5'h1b == _T_1437[4:0] ? 5'h0 : _GEN_15270; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_15272 = 5'h1c == _T_1437[4:0] ? 5'h0 : _GEN_15271; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_15273 = 5'h1d == _T_1437[4:0] ? 5'h0 : _GEN_15272; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_15274 = 5'h1e == _T_1437[4:0] ? 5'h0 : _GEN_15273; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_15275 = 5'h1f == _T_1437[4:0] ? 5'h0 : _GEN_15274; // @[FanCtrl.scala 54:{41,41}]
  wire  _T_1439 = _GEN_15118 != _GEN_15275; // @[FanCtrl.scala 54:41]
  wire  _T_1448 = _GEN_15086 != _GEN_15118; // @[FanCtrl.scala 56:41]
  wire  _T_1458 = _GEN_15118 == _GEN_15275; // @[FanCtrl.scala 61:48]
  wire  _GEN_15509 = r_valid_1 & _T_1426; // @[FanCtrl.scala 47:34]
  wire [5:0] _T_1494 = _T_1418 - 6'h1; // @[FanCtrl.scala 94:58]
  wire [4:0] _GEN_15756 = 5'h3 == _T_1494[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_15757 = 5'h4 == _T_1494[4:0] ? w_vn_4 : _GEN_15756; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_15758 = 5'h5 == _T_1494[4:0] ? 5'h0 : _GEN_15757; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_15759 = 5'h6 == _T_1494[4:0] ? 5'h0 : _GEN_15758; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_15760 = 5'h7 == _T_1494[4:0] ? w_vn_7 : _GEN_15759; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_15761 = 5'h8 == _T_1494[4:0] ? w_vn_8 : _GEN_15760; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_15762 = 5'h9 == _T_1494[4:0] ? 5'h0 : _GEN_15761; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_15763 = 5'ha == _T_1494[4:0] ? 5'h0 : _GEN_15762; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_15764 = 5'hb == _T_1494[4:0] ? w_vn_11 : _GEN_15763; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_15765 = 5'hc == _T_1494[4:0] ? w_vn_12 : _GEN_15764; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_15766 = 5'hd == _T_1494[4:0] ? w_vn_13 : _GEN_15765; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_15767 = 5'he == _T_1494[4:0] ? 5'h0 : _GEN_15766; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_15768 = 5'hf == _T_1494[4:0] ? w_vn_15 : _GEN_15767; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_15769 = 5'h10 == _T_1494[4:0] ? w_vn_16 : _GEN_15768; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_15770 = 5'h11 == _T_1494[4:0] ? 5'h0 : _GEN_15769; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_15771 = 5'h12 == _T_1494[4:0] ? w_vn_18 : _GEN_15770; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_15772 = 5'h13 == _T_1494[4:0] ? 5'h0 : _GEN_15771; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_15773 = 5'h14 == _T_1494[4:0] ? 5'h0 : _GEN_15772; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_15774 = 5'h15 == _T_1494[4:0] ? 5'h0 : _GEN_15773; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_15775 = 5'h16 == _T_1494[4:0] ? 5'h0 : _GEN_15774; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_15776 = 5'h17 == _T_1494[4:0] ? w_vn_23 : _GEN_15775; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_15777 = 5'h18 == _T_1494[4:0] ? w_vn_24 : _GEN_15776; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_15778 = 5'h19 == _T_1494[4:0] ? 5'h0 : _GEN_15777; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_15779 = 5'h1a == _T_1494[4:0] ? 5'h0 : _GEN_15778; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_15780 = 5'h1b == _T_1494[4:0] ? 5'h0 : _GEN_15779; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_15781 = 5'h1c == _T_1494[4:0] ? 5'h0 : _GEN_15780; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_15782 = 5'h1d == _T_1494[4:0] ? 5'h0 : _GEN_15781; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_15783 = 5'h1e == _T_1494[4:0] ? 5'h0 : _GEN_15782; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_15784 = 5'h1f == _T_1494[4:0] ? 5'h0 : _GEN_15783; // @[FanCtrl.scala 94:{39,39}]
  wire  _T_1496 = _GEN_15086 != _GEN_15784; // @[FanCtrl.scala 94:39]
  wire  _T_1515 = _GEN_15086 == _GEN_15784; // @[FanCtrl.scala 99:46]
  wire  _T_1562 = _T_1496 & _T_1439; // @[FanCtrl.scala 125:65]
  wire  _T_1572 = _T_1562 & _T_1448; // @[FanCtrl.scala 126:65]
  wire  _T_1591 = _T_1515 & _T_1439; // @[FanCtrl.scala 131:70]
  wire  _T_1601 = _T_1591 & _T_1448; // @[FanCtrl.scala 132:72]
  wire  _T_1620 = _T_1496 & _T_1458; // @[FanCtrl.scala 137:72]
  wire  _T_1630 = _T_1620 & _T_1448; // @[FanCtrl.scala 138:71]
  wire [1:0] _GEN_16806 = _T_1630 ? 2'h3 : 2'h1; // @[FanCtrl.scala 139:73 141:34 144:35]
  wire [2:0] _GEN_16807 = _T_1601 ? 3'h4 : {{1'd0}, _GEN_16806}; // @[FanCtrl.scala 133:73 135:35]
  wire [2:0] _GEN_16808 = _T_1572 ? 3'h5 : _GEN_16807; // @[FanCtrl.scala 127:66 129:35]
  wire [2:0] _GEN_16871 = r_valid_1 ? _GEN_16808 : 3'h0; // @[FanCtrl.scala 117:32 148:33]
  wire [5:0] _T_1635 = 2'h2 * 4'h9; // @[FanCtrl.scala 48:25]
  wire [6:0] _T_1636 = {{1'd0}, _T_1635}; // @[FanCtrl.scala 48:31]
  wire [5:0] _T_1641 = _T_1635 + 6'h1; // @[FanCtrl.scala 48:58]
  wire [4:0] _GEN_16940 = 5'h3 == _T_1636[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_16941 = 5'h4 == _T_1636[4:0] ? w_vn_4 : _GEN_16940; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_16942 = 5'h5 == _T_1636[4:0] ? 5'h0 : _GEN_16941; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_16943 = 5'h6 == _T_1636[4:0] ? 5'h0 : _GEN_16942; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_16944 = 5'h7 == _T_1636[4:0] ? w_vn_7 : _GEN_16943; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_16945 = 5'h8 == _T_1636[4:0] ? w_vn_8 : _GEN_16944; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_16946 = 5'h9 == _T_1636[4:0] ? 5'h0 : _GEN_16945; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_16947 = 5'ha == _T_1636[4:0] ? 5'h0 : _GEN_16946; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_16948 = 5'hb == _T_1636[4:0] ? w_vn_11 : _GEN_16947; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_16949 = 5'hc == _T_1636[4:0] ? w_vn_12 : _GEN_16948; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_16950 = 5'hd == _T_1636[4:0] ? w_vn_13 : _GEN_16949; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_16951 = 5'he == _T_1636[4:0] ? 5'h0 : _GEN_16950; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_16952 = 5'hf == _T_1636[4:0] ? w_vn_15 : _GEN_16951; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_16953 = 5'h10 == _T_1636[4:0] ? w_vn_16 : _GEN_16952; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_16954 = 5'h11 == _T_1636[4:0] ? 5'h0 : _GEN_16953; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_16955 = 5'h12 == _T_1636[4:0] ? w_vn_18 : _GEN_16954; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_16956 = 5'h13 == _T_1636[4:0] ? 5'h0 : _GEN_16955; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_16957 = 5'h14 == _T_1636[4:0] ? 5'h0 : _GEN_16956; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_16958 = 5'h15 == _T_1636[4:0] ? 5'h0 : _GEN_16957; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_16959 = 5'h16 == _T_1636[4:0] ? 5'h0 : _GEN_16958; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_16960 = 5'h17 == _T_1636[4:0] ? w_vn_23 : _GEN_16959; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_16961 = 5'h18 == _T_1636[4:0] ? w_vn_24 : _GEN_16960; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_16962 = 5'h19 == _T_1636[4:0] ? 5'h0 : _GEN_16961; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_16963 = 5'h1a == _T_1636[4:0] ? 5'h0 : _GEN_16962; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_16964 = 5'h1b == _T_1636[4:0] ? 5'h0 : _GEN_16963; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_16965 = 5'h1c == _T_1636[4:0] ? 5'h0 : _GEN_16964; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_16966 = 5'h1d == _T_1636[4:0] ? 5'h0 : _GEN_16965; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_16967 = 5'h1e == _T_1636[4:0] ? 5'h0 : _GEN_16966; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_16968 = 5'h1f == _T_1636[4:0] ? 5'h0 : _GEN_16967; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_16972 = 5'h3 == _T_1641[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_16973 = 5'h4 == _T_1641[4:0] ? w_vn_4 : _GEN_16972; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_16974 = 5'h5 == _T_1641[4:0] ? 5'h0 : _GEN_16973; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_16975 = 5'h6 == _T_1641[4:0] ? 5'h0 : _GEN_16974; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_16976 = 5'h7 == _T_1641[4:0] ? w_vn_7 : _GEN_16975; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_16977 = 5'h8 == _T_1641[4:0] ? w_vn_8 : _GEN_16976; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_16978 = 5'h9 == _T_1641[4:0] ? 5'h0 : _GEN_16977; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_16979 = 5'ha == _T_1641[4:0] ? 5'h0 : _GEN_16978; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_16980 = 5'hb == _T_1641[4:0] ? w_vn_11 : _GEN_16979; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_16981 = 5'hc == _T_1641[4:0] ? w_vn_12 : _GEN_16980; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_16982 = 5'hd == _T_1641[4:0] ? w_vn_13 : _GEN_16981; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_16983 = 5'he == _T_1641[4:0] ? 5'h0 : _GEN_16982; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_16984 = 5'hf == _T_1641[4:0] ? w_vn_15 : _GEN_16983; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_16985 = 5'h10 == _T_1641[4:0] ? w_vn_16 : _GEN_16984; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_16986 = 5'h11 == _T_1641[4:0] ? 5'h0 : _GEN_16985; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_16987 = 5'h12 == _T_1641[4:0] ? w_vn_18 : _GEN_16986; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_16988 = 5'h13 == _T_1641[4:0] ? 5'h0 : _GEN_16987; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_16989 = 5'h14 == _T_1641[4:0] ? 5'h0 : _GEN_16988; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_16990 = 5'h15 == _T_1641[4:0] ? 5'h0 : _GEN_16989; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_16991 = 5'h16 == _T_1641[4:0] ? 5'h0 : _GEN_16990; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_16992 = 5'h17 == _T_1641[4:0] ? w_vn_23 : _GEN_16991; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_16993 = 5'h18 == _T_1641[4:0] ? w_vn_24 : _GEN_16992; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_16994 = 5'h19 == _T_1641[4:0] ? 5'h0 : _GEN_16993; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_16995 = 5'h1a == _T_1641[4:0] ? 5'h0 : _GEN_16994; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_16996 = 5'h1b == _T_1641[4:0] ? 5'h0 : _GEN_16995; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_16997 = 5'h1c == _T_1641[4:0] ? 5'h0 : _GEN_16996; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_16998 = 5'h1d == _T_1641[4:0] ? 5'h0 : _GEN_16997; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_16999 = 5'h1e == _T_1641[4:0] ? 5'h0 : _GEN_16998; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_17000 = 5'h1f == _T_1641[4:0] ? 5'h0 : _GEN_16999; // @[FanCtrl.scala 48:{39,39}]
  wire  _T_1643 = _GEN_16968 == _GEN_17000; // @[FanCtrl.scala 48:39]
  wire [5:0] _T_1654 = _T_1635 + 6'h2; // @[FanCtrl.scala 55:32]
  wire [4:0] _GEN_17129 = 5'h3 == _T_1654[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_17130 = 5'h4 == _T_1654[4:0] ? w_vn_4 : _GEN_17129; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_17131 = 5'h5 == _T_1654[4:0] ? 5'h0 : _GEN_17130; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_17132 = 5'h6 == _T_1654[4:0] ? 5'h0 : _GEN_17131; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_17133 = 5'h7 == _T_1654[4:0] ? w_vn_7 : _GEN_17132; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_17134 = 5'h8 == _T_1654[4:0] ? w_vn_8 : _GEN_17133; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_17135 = 5'h9 == _T_1654[4:0] ? 5'h0 : _GEN_17134; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_17136 = 5'ha == _T_1654[4:0] ? 5'h0 : _GEN_17135; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_17137 = 5'hb == _T_1654[4:0] ? w_vn_11 : _GEN_17136; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_17138 = 5'hc == _T_1654[4:0] ? w_vn_12 : _GEN_17137; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_17139 = 5'hd == _T_1654[4:0] ? w_vn_13 : _GEN_17138; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_17140 = 5'he == _T_1654[4:0] ? 5'h0 : _GEN_17139; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_17141 = 5'hf == _T_1654[4:0] ? w_vn_15 : _GEN_17140; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_17142 = 5'h10 == _T_1654[4:0] ? w_vn_16 : _GEN_17141; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_17143 = 5'h11 == _T_1654[4:0] ? 5'h0 : _GEN_17142; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_17144 = 5'h12 == _T_1654[4:0] ? w_vn_18 : _GEN_17143; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_17145 = 5'h13 == _T_1654[4:0] ? 5'h0 : _GEN_17144; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_17146 = 5'h14 == _T_1654[4:0] ? 5'h0 : _GEN_17145; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_17147 = 5'h15 == _T_1654[4:0] ? 5'h0 : _GEN_17146; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_17148 = 5'h16 == _T_1654[4:0] ? 5'h0 : _GEN_17147; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_17149 = 5'h17 == _T_1654[4:0] ? w_vn_23 : _GEN_17148; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_17150 = 5'h18 == _T_1654[4:0] ? w_vn_24 : _GEN_17149; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_17151 = 5'h19 == _T_1654[4:0] ? 5'h0 : _GEN_17150; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_17152 = 5'h1a == _T_1654[4:0] ? 5'h0 : _GEN_17151; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_17153 = 5'h1b == _T_1654[4:0] ? 5'h0 : _GEN_17152; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_17154 = 5'h1c == _T_1654[4:0] ? 5'h0 : _GEN_17153; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_17155 = 5'h1d == _T_1654[4:0] ? 5'h0 : _GEN_17154; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_17156 = 5'h1e == _T_1654[4:0] ? 5'h0 : _GEN_17155; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_17157 = 5'h1f == _T_1654[4:0] ? 5'h0 : _GEN_17156; // @[FanCtrl.scala 54:{41,41}]
  wire  _T_1656 = _GEN_17000 != _GEN_17157; // @[FanCtrl.scala 54:41]
  wire  _T_1665 = _GEN_16968 != _GEN_17000; // @[FanCtrl.scala 56:41]
  wire  _T_1675 = _GEN_17000 == _GEN_17157; // @[FanCtrl.scala 61:48]
  wire  _GEN_17392 = r_valid_1 & _T_1643; // @[FanCtrl.scala 47:34]
  wire [5:0] _T_1711 = _T_1635 - 6'h1; // @[FanCtrl.scala 94:58]
  wire [4:0] _GEN_17638 = 5'h3 == _T_1711[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_17639 = 5'h4 == _T_1711[4:0] ? w_vn_4 : _GEN_17638; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_17640 = 5'h5 == _T_1711[4:0] ? 5'h0 : _GEN_17639; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_17641 = 5'h6 == _T_1711[4:0] ? 5'h0 : _GEN_17640; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_17642 = 5'h7 == _T_1711[4:0] ? w_vn_7 : _GEN_17641; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_17643 = 5'h8 == _T_1711[4:0] ? w_vn_8 : _GEN_17642; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_17644 = 5'h9 == _T_1711[4:0] ? 5'h0 : _GEN_17643; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_17645 = 5'ha == _T_1711[4:0] ? 5'h0 : _GEN_17644; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_17646 = 5'hb == _T_1711[4:0] ? w_vn_11 : _GEN_17645; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_17647 = 5'hc == _T_1711[4:0] ? w_vn_12 : _GEN_17646; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_17648 = 5'hd == _T_1711[4:0] ? w_vn_13 : _GEN_17647; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_17649 = 5'he == _T_1711[4:0] ? 5'h0 : _GEN_17648; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_17650 = 5'hf == _T_1711[4:0] ? w_vn_15 : _GEN_17649; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_17651 = 5'h10 == _T_1711[4:0] ? w_vn_16 : _GEN_17650; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_17652 = 5'h11 == _T_1711[4:0] ? 5'h0 : _GEN_17651; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_17653 = 5'h12 == _T_1711[4:0] ? w_vn_18 : _GEN_17652; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_17654 = 5'h13 == _T_1711[4:0] ? 5'h0 : _GEN_17653; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_17655 = 5'h14 == _T_1711[4:0] ? 5'h0 : _GEN_17654; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_17656 = 5'h15 == _T_1711[4:0] ? 5'h0 : _GEN_17655; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_17657 = 5'h16 == _T_1711[4:0] ? 5'h0 : _GEN_17656; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_17658 = 5'h17 == _T_1711[4:0] ? w_vn_23 : _GEN_17657; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_17659 = 5'h18 == _T_1711[4:0] ? w_vn_24 : _GEN_17658; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_17660 = 5'h19 == _T_1711[4:0] ? 5'h0 : _GEN_17659; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_17661 = 5'h1a == _T_1711[4:0] ? 5'h0 : _GEN_17660; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_17662 = 5'h1b == _T_1711[4:0] ? 5'h0 : _GEN_17661; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_17663 = 5'h1c == _T_1711[4:0] ? 5'h0 : _GEN_17662; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_17664 = 5'h1d == _T_1711[4:0] ? 5'h0 : _GEN_17663; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_17665 = 5'h1e == _T_1711[4:0] ? 5'h0 : _GEN_17664; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_17666 = 5'h1f == _T_1711[4:0] ? 5'h0 : _GEN_17665; // @[FanCtrl.scala 94:{39,39}]
  wire  _T_1713 = _GEN_16968 != _GEN_17666; // @[FanCtrl.scala 94:39]
  wire  _T_1732 = _GEN_16968 == _GEN_17666; // @[FanCtrl.scala 99:46]
  wire  _T_1779 = _T_1713 & _T_1656; // @[FanCtrl.scala 125:65]
  wire  _T_1789 = _T_1779 & _T_1665; // @[FanCtrl.scala 126:65]
  wire  _T_1808 = _T_1732 & _T_1656; // @[FanCtrl.scala 131:70]
  wire  _T_1818 = _T_1808 & _T_1665; // @[FanCtrl.scala 132:72]
  wire  _T_1837 = _T_1713 & _T_1675; // @[FanCtrl.scala 137:72]
  wire  _T_1847 = _T_1837 & _T_1665; // @[FanCtrl.scala 138:71]
  wire [1:0] _GEN_18688 = _T_1847 ? 2'h3 : 2'h1; // @[FanCtrl.scala 139:73 141:34 144:35]
  wire [2:0] _GEN_18689 = _T_1818 ? 3'h4 : {{1'd0}, _GEN_18688}; // @[FanCtrl.scala 133:73 135:35]
  wire [2:0] _GEN_18690 = _T_1789 ? 3'h5 : _GEN_18689; // @[FanCtrl.scala 127:66 129:35]
  wire [2:0] _GEN_18753 = r_valid_1 ? _GEN_18690 : 3'h0; // @[FanCtrl.scala 117:32 148:33]
  wire [5:0] _T_1852 = 2'h2 * 4'ha; // @[FanCtrl.scala 48:25]
  wire [6:0] _T_1853 = {{1'd0}, _T_1852}; // @[FanCtrl.scala 48:31]
  wire [5:0] _T_1858 = _T_1852 + 6'h1; // @[FanCtrl.scala 48:58]
  wire [4:0] _GEN_18822 = 5'h3 == _T_1853[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_18823 = 5'h4 == _T_1853[4:0] ? w_vn_4 : _GEN_18822; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_18824 = 5'h5 == _T_1853[4:0] ? 5'h0 : _GEN_18823; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_18825 = 5'h6 == _T_1853[4:0] ? 5'h0 : _GEN_18824; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_18826 = 5'h7 == _T_1853[4:0] ? w_vn_7 : _GEN_18825; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_18827 = 5'h8 == _T_1853[4:0] ? w_vn_8 : _GEN_18826; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_18828 = 5'h9 == _T_1853[4:0] ? 5'h0 : _GEN_18827; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_18829 = 5'ha == _T_1853[4:0] ? 5'h0 : _GEN_18828; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_18830 = 5'hb == _T_1853[4:0] ? w_vn_11 : _GEN_18829; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_18831 = 5'hc == _T_1853[4:0] ? w_vn_12 : _GEN_18830; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_18832 = 5'hd == _T_1853[4:0] ? w_vn_13 : _GEN_18831; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_18833 = 5'he == _T_1853[4:0] ? 5'h0 : _GEN_18832; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_18834 = 5'hf == _T_1853[4:0] ? w_vn_15 : _GEN_18833; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_18835 = 5'h10 == _T_1853[4:0] ? w_vn_16 : _GEN_18834; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_18836 = 5'h11 == _T_1853[4:0] ? 5'h0 : _GEN_18835; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_18837 = 5'h12 == _T_1853[4:0] ? w_vn_18 : _GEN_18836; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_18838 = 5'h13 == _T_1853[4:0] ? 5'h0 : _GEN_18837; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_18839 = 5'h14 == _T_1853[4:0] ? 5'h0 : _GEN_18838; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_18840 = 5'h15 == _T_1853[4:0] ? 5'h0 : _GEN_18839; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_18841 = 5'h16 == _T_1853[4:0] ? 5'h0 : _GEN_18840; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_18842 = 5'h17 == _T_1853[4:0] ? w_vn_23 : _GEN_18841; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_18843 = 5'h18 == _T_1853[4:0] ? w_vn_24 : _GEN_18842; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_18844 = 5'h19 == _T_1853[4:0] ? 5'h0 : _GEN_18843; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_18845 = 5'h1a == _T_1853[4:0] ? 5'h0 : _GEN_18844; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_18846 = 5'h1b == _T_1853[4:0] ? 5'h0 : _GEN_18845; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_18847 = 5'h1c == _T_1853[4:0] ? 5'h0 : _GEN_18846; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_18848 = 5'h1d == _T_1853[4:0] ? 5'h0 : _GEN_18847; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_18849 = 5'h1e == _T_1853[4:0] ? 5'h0 : _GEN_18848; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_18850 = 5'h1f == _T_1853[4:0] ? 5'h0 : _GEN_18849; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_18854 = 5'h3 == _T_1858[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_18855 = 5'h4 == _T_1858[4:0] ? w_vn_4 : _GEN_18854; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_18856 = 5'h5 == _T_1858[4:0] ? 5'h0 : _GEN_18855; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_18857 = 5'h6 == _T_1858[4:0] ? 5'h0 : _GEN_18856; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_18858 = 5'h7 == _T_1858[4:0] ? w_vn_7 : _GEN_18857; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_18859 = 5'h8 == _T_1858[4:0] ? w_vn_8 : _GEN_18858; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_18860 = 5'h9 == _T_1858[4:0] ? 5'h0 : _GEN_18859; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_18861 = 5'ha == _T_1858[4:0] ? 5'h0 : _GEN_18860; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_18862 = 5'hb == _T_1858[4:0] ? w_vn_11 : _GEN_18861; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_18863 = 5'hc == _T_1858[4:0] ? w_vn_12 : _GEN_18862; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_18864 = 5'hd == _T_1858[4:0] ? w_vn_13 : _GEN_18863; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_18865 = 5'he == _T_1858[4:0] ? 5'h0 : _GEN_18864; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_18866 = 5'hf == _T_1858[4:0] ? w_vn_15 : _GEN_18865; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_18867 = 5'h10 == _T_1858[4:0] ? w_vn_16 : _GEN_18866; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_18868 = 5'h11 == _T_1858[4:0] ? 5'h0 : _GEN_18867; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_18869 = 5'h12 == _T_1858[4:0] ? w_vn_18 : _GEN_18868; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_18870 = 5'h13 == _T_1858[4:0] ? 5'h0 : _GEN_18869; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_18871 = 5'h14 == _T_1858[4:0] ? 5'h0 : _GEN_18870; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_18872 = 5'h15 == _T_1858[4:0] ? 5'h0 : _GEN_18871; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_18873 = 5'h16 == _T_1858[4:0] ? 5'h0 : _GEN_18872; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_18874 = 5'h17 == _T_1858[4:0] ? w_vn_23 : _GEN_18873; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_18875 = 5'h18 == _T_1858[4:0] ? w_vn_24 : _GEN_18874; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_18876 = 5'h19 == _T_1858[4:0] ? 5'h0 : _GEN_18875; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_18877 = 5'h1a == _T_1858[4:0] ? 5'h0 : _GEN_18876; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_18878 = 5'h1b == _T_1858[4:0] ? 5'h0 : _GEN_18877; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_18879 = 5'h1c == _T_1858[4:0] ? 5'h0 : _GEN_18878; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_18880 = 5'h1d == _T_1858[4:0] ? 5'h0 : _GEN_18879; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_18881 = 5'h1e == _T_1858[4:0] ? 5'h0 : _GEN_18880; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_18882 = 5'h1f == _T_1858[4:0] ? 5'h0 : _GEN_18881; // @[FanCtrl.scala 48:{39,39}]
  wire  _T_1860 = _GEN_18850 == _GEN_18882; // @[FanCtrl.scala 48:39]
  wire [5:0] _T_1871 = _T_1852 + 6'h2; // @[FanCtrl.scala 55:32]
  wire [4:0] _GEN_19011 = 5'h3 == _T_1871[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_19012 = 5'h4 == _T_1871[4:0] ? w_vn_4 : _GEN_19011; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_19013 = 5'h5 == _T_1871[4:0] ? 5'h0 : _GEN_19012; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_19014 = 5'h6 == _T_1871[4:0] ? 5'h0 : _GEN_19013; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_19015 = 5'h7 == _T_1871[4:0] ? w_vn_7 : _GEN_19014; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_19016 = 5'h8 == _T_1871[4:0] ? w_vn_8 : _GEN_19015; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_19017 = 5'h9 == _T_1871[4:0] ? 5'h0 : _GEN_19016; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_19018 = 5'ha == _T_1871[4:0] ? 5'h0 : _GEN_19017; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_19019 = 5'hb == _T_1871[4:0] ? w_vn_11 : _GEN_19018; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_19020 = 5'hc == _T_1871[4:0] ? w_vn_12 : _GEN_19019; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_19021 = 5'hd == _T_1871[4:0] ? w_vn_13 : _GEN_19020; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_19022 = 5'he == _T_1871[4:0] ? 5'h0 : _GEN_19021; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_19023 = 5'hf == _T_1871[4:0] ? w_vn_15 : _GEN_19022; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_19024 = 5'h10 == _T_1871[4:0] ? w_vn_16 : _GEN_19023; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_19025 = 5'h11 == _T_1871[4:0] ? 5'h0 : _GEN_19024; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_19026 = 5'h12 == _T_1871[4:0] ? w_vn_18 : _GEN_19025; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_19027 = 5'h13 == _T_1871[4:0] ? 5'h0 : _GEN_19026; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_19028 = 5'h14 == _T_1871[4:0] ? 5'h0 : _GEN_19027; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_19029 = 5'h15 == _T_1871[4:0] ? 5'h0 : _GEN_19028; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_19030 = 5'h16 == _T_1871[4:0] ? 5'h0 : _GEN_19029; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_19031 = 5'h17 == _T_1871[4:0] ? w_vn_23 : _GEN_19030; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_19032 = 5'h18 == _T_1871[4:0] ? w_vn_24 : _GEN_19031; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_19033 = 5'h19 == _T_1871[4:0] ? 5'h0 : _GEN_19032; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_19034 = 5'h1a == _T_1871[4:0] ? 5'h0 : _GEN_19033; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_19035 = 5'h1b == _T_1871[4:0] ? 5'h0 : _GEN_19034; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_19036 = 5'h1c == _T_1871[4:0] ? 5'h0 : _GEN_19035; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_19037 = 5'h1d == _T_1871[4:0] ? 5'h0 : _GEN_19036; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_19038 = 5'h1e == _T_1871[4:0] ? 5'h0 : _GEN_19037; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_19039 = 5'h1f == _T_1871[4:0] ? 5'h0 : _GEN_19038; // @[FanCtrl.scala 54:{41,41}]
  wire  _T_1873 = _GEN_18882 != _GEN_19039; // @[FanCtrl.scala 54:41]
  wire  _T_1882 = _GEN_18850 != _GEN_18882; // @[FanCtrl.scala 56:41]
  wire  _T_1892 = _GEN_18882 == _GEN_19039; // @[FanCtrl.scala 61:48]
  wire  _GEN_19275 = r_valid_1 & _T_1860; // @[FanCtrl.scala 47:34]
  wire [5:0] _T_1928 = _T_1852 - 6'h1; // @[FanCtrl.scala 94:58]
  wire [4:0] _GEN_19520 = 5'h3 == _T_1928[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_19521 = 5'h4 == _T_1928[4:0] ? w_vn_4 : _GEN_19520; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_19522 = 5'h5 == _T_1928[4:0] ? 5'h0 : _GEN_19521; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_19523 = 5'h6 == _T_1928[4:0] ? 5'h0 : _GEN_19522; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_19524 = 5'h7 == _T_1928[4:0] ? w_vn_7 : _GEN_19523; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_19525 = 5'h8 == _T_1928[4:0] ? w_vn_8 : _GEN_19524; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_19526 = 5'h9 == _T_1928[4:0] ? 5'h0 : _GEN_19525; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_19527 = 5'ha == _T_1928[4:0] ? 5'h0 : _GEN_19526; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_19528 = 5'hb == _T_1928[4:0] ? w_vn_11 : _GEN_19527; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_19529 = 5'hc == _T_1928[4:0] ? w_vn_12 : _GEN_19528; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_19530 = 5'hd == _T_1928[4:0] ? w_vn_13 : _GEN_19529; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_19531 = 5'he == _T_1928[4:0] ? 5'h0 : _GEN_19530; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_19532 = 5'hf == _T_1928[4:0] ? w_vn_15 : _GEN_19531; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_19533 = 5'h10 == _T_1928[4:0] ? w_vn_16 : _GEN_19532; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_19534 = 5'h11 == _T_1928[4:0] ? 5'h0 : _GEN_19533; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_19535 = 5'h12 == _T_1928[4:0] ? w_vn_18 : _GEN_19534; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_19536 = 5'h13 == _T_1928[4:0] ? 5'h0 : _GEN_19535; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_19537 = 5'h14 == _T_1928[4:0] ? 5'h0 : _GEN_19536; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_19538 = 5'h15 == _T_1928[4:0] ? 5'h0 : _GEN_19537; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_19539 = 5'h16 == _T_1928[4:0] ? 5'h0 : _GEN_19538; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_19540 = 5'h17 == _T_1928[4:0] ? w_vn_23 : _GEN_19539; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_19541 = 5'h18 == _T_1928[4:0] ? w_vn_24 : _GEN_19540; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_19542 = 5'h19 == _T_1928[4:0] ? 5'h0 : _GEN_19541; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_19543 = 5'h1a == _T_1928[4:0] ? 5'h0 : _GEN_19542; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_19544 = 5'h1b == _T_1928[4:0] ? 5'h0 : _GEN_19543; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_19545 = 5'h1c == _T_1928[4:0] ? 5'h0 : _GEN_19544; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_19546 = 5'h1d == _T_1928[4:0] ? 5'h0 : _GEN_19545; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_19547 = 5'h1e == _T_1928[4:0] ? 5'h0 : _GEN_19546; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_19548 = 5'h1f == _T_1928[4:0] ? 5'h0 : _GEN_19547; // @[FanCtrl.scala 94:{39,39}]
  wire  _T_1930 = _GEN_18850 != _GEN_19548; // @[FanCtrl.scala 94:39]
  wire  _T_1949 = _GEN_18850 == _GEN_19548; // @[FanCtrl.scala 99:46]
  wire  _T_1996 = _T_1930 & _T_1873; // @[FanCtrl.scala 125:65]
  wire  _T_2006 = _T_1996 & _T_1882; // @[FanCtrl.scala 126:65]
  wire  _T_2025 = _T_1949 & _T_1873; // @[FanCtrl.scala 131:70]
  wire  _T_2035 = _T_2025 & _T_1882; // @[FanCtrl.scala 132:72]
  wire  _T_2054 = _T_1930 & _T_1892; // @[FanCtrl.scala 137:72]
  wire  _T_2064 = _T_2054 & _T_1882; // @[FanCtrl.scala 138:71]
  wire [1:0] _GEN_20570 = _T_2064 ? 2'h3 : 2'h1; // @[FanCtrl.scala 139:73 141:34 144:35]
  wire [2:0] _GEN_20571 = _T_2035 ? 3'h4 : {{1'd0}, _GEN_20570}; // @[FanCtrl.scala 133:73 135:35]
  wire [2:0] _GEN_20572 = _T_2006 ? 3'h5 : _GEN_20571; // @[FanCtrl.scala 127:66 129:35]
  wire [2:0] _GEN_20635 = r_valid_1 ? _GEN_20572 : 3'h0; // @[FanCtrl.scala 117:32 148:33]
  wire [5:0] _T_2069 = 2'h2 * 4'hb; // @[FanCtrl.scala 48:25]
  wire [6:0] _T_2070 = {{1'd0}, _T_2069}; // @[FanCtrl.scala 48:31]
  wire [5:0] _T_2075 = _T_2069 + 6'h1; // @[FanCtrl.scala 48:58]
  wire [4:0] _GEN_20704 = 5'h3 == _T_2070[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_20705 = 5'h4 == _T_2070[4:0] ? w_vn_4 : _GEN_20704; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_20706 = 5'h5 == _T_2070[4:0] ? 5'h0 : _GEN_20705; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_20707 = 5'h6 == _T_2070[4:0] ? 5'h0 : _GEN_20706; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_20708 = 5'h7 == _T_2070[4:0] ? w_vn_7 : _GEN_20707; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_20709 = 5'h8 == _T_2070[4:0] ? w_vn_8 : _GEN_20708; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_20710 = 5'h9 == _T_2070[4:0] ? 5'h0 : _GEN_20709; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_20711 = 5'ha == _T_2070[4:0] ? 5'h0 : _GEN_20710; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_20712 = 5'hb == _T_2070[4:0] ? w_vn_11 : _GEN_20711; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_20713 = 5'hc == _T_2070[4:0] ? w_vn_12 : _GEN_20712; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_20714 = 5'hd == _T_2070[4:0] ? w_vn_13 : _GEN_20713; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_20715 = 5'he == _T_2070[4:0] ? 5'h0 : _GEN_20714; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_20716 = 5'hf == _T_2070[4:0] ? w_vn_15 : _GEN_20715; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_20717 = 5'h10 == _T_2070[4:0] ? w_vn_16 : _GEN_20716; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_20718 = 5'h11 == _T_2070[4:0] ? 5'h0 : _GEN_20717; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_20719 = 5'h12 == _T_2070[4:0] ? w_vn_18 : _GEN_20718; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_20720 = 5'h13 == _T_2070[4:0] ? 5'h0 : _GEN_20719; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_20721 = 5'h14 == _T_2070[4:0] ? 5'h0 : _GEN_20720; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_20722 = 5'h15 == _T_2070[4:0] ? 5'h0 : _GEN_20721; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_20723 = 5'h16 == _T_2070[4:0] ? 5'h0 : _GEN_20722; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_20724 = 5'h17 == _T_2070[4:0] ? w_vn_23 : _GEN_20723; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_20725 = 5'h18 == _T_2070[4:0] ? w_vn_24 : _GEN_20724; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_20726 = 5'h19 == _T_2070[4:0] ? 5'h0 : _GEN_20725; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_20727 = 5'h1a == _T_2070[4:0] ? 5'h0 : _GEN_20726; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_20728 = 5'h1b == _T_2070[4:0] ? 5'h0 : _GEN_20727; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_20729 = 5'h1c == _T_2070[4:0] ? 5'h0 : _GEN_20728; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_20730 = 5'h1d == _T_2070[4:0] ? 5'h0 : _GEN_20729; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_20731 = 5'h1e == _T_2070[4:0] ? 5'h0 : _GEN_20730; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_20732 = 5'h1f == _T_2070[4:0] ? 5'h0 : _GEN_20731; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_20736 = 5'h3 == _T_2075[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_20737 = 5'h4 == _T_2075[4:0] ? w_vn_4 : _GEN_20736; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_20738 = 5'h5 == _T_2075[4:0] ? 5'h0 : _GEN_20737; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_20739 = 5'h6 == _T_2075[4:0] ? 5'h0 : _GEN_20738; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_20740 = 5'h7 == _T_2075[4:0] ? w_vn_7 : _GEN_20739; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_20741 = 5'h8 == _T_2075[4:0] ? w_vn_8 : _GEN_20740; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_20742 = 5'h9 == _T_2075[4:0] ? 5'h0 : _GEN_20741; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_20743 = 5'ha == _T_2075[4:0] ? 5'h0 : _GEN_20742; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_20744 = 5'hb == _T_2075[4:0] ? w_vn_11 : _GEN_20743; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_20745 = 5'hc == _T_2075[4:0] ? w_vn_12 : _GEN_20744; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_20746 = 5'hd == _T_2075[4:0] ? w_vn_13 : _GEN_20745; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_20747 = 5'he == _T_2075[4:0] ? 5'h0 : _GEN_20746; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_20748 = 5'hf == _T_2075[4:0] ? w_vn_15 : _GEN_20747; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_20749 = 5'h10 == _T_2075[4:0] ? w_vn_16 : _GEN_20748; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_20750 = 5'h11 == _T_2075[4:0] ? 5'h0 : _GEN_20749; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_20751 = 5'h12 == _T_2075[4:0] ? w_vn_18 : _GEN_20750; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_20752 = 5'h13 == _T_2075[4:0] ? 5'h0 : _GEN_20751; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_20753 = 5'h14 == _T_2075[4:0] ? 5'h0 : _GEN_20752; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_20754 = 5'h15 == _T_2075[4:0] ? 5'h0 : _GEN_20753; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_20755 = 5'h16 == _T_2075[4:0] ? 5'h0 : _GEN_20754; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_20756 = 5'h17 == _T_2075[4:0] ? w_vn_23 : _GEN_20755; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_20757 = 5'h18 == _T_2075[4:0] ? w_vn_24 : _GEN_20756; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_20758 = 5'h19 == _T_2075[4:0] ? 5'h0 : _GEN_20757; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_20759 = 5'h1a == _T_2075[4:0] ? 5'h0 : _GEN_20758; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_20760 = 5'h1b == _T_2075[4:0] ? 5'h0 : _GEN_20759; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_20761 = 5'h1c == _T_2075[4:0] ? 5'h0 : _GEN_20760; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_20762 = 5'h1d == _T_2075[4:0] ? 5'h0 : _GEN_20761; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_20763 = 5'h1e == _T_2075[4:0] ? 5'h0 : _GEN_20762; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_20764 = 5'h1f == _T_2075[4:0] ? 5'h0 : _GEN_20763; // @[FanCtrl.scala 48:{39,39}]
  wire  _T_2077 = _GEN_20732 == _GEN_20764; // @[FanCtrl.scala 48:39]
  wire [5:0] _T_2088 = _T_2069 + 6'h2; // @[FanCtrl.scala 55:32]
  wire [4:0] _GEN_20893 = 5'h3 == _T_2088[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_20894 = 5'h4 == _T_2088[4:0] ? w_vn_4 : _GEN_20893; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_20895 = 5'h5 == _T_2088[4:0] ? 5'h0 : _GEN_20894; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_20896 = 5'h6 == _T_2088[4:0] ? 5'h0 : _GEN_20895; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_20897 = 5'h7 == _T_2088[4:0] ? w_vn_7 : _GEN_20896; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_20898 = 5'h8 == _T_2088[4:0] ? w_vn_8 : _GEN_20897; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_20899 = 5'h9 == _T_2088[4:0] ? 5'h0 : _GEN_20898; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_20900 = 5'ha == _T_2088[4:0] ? 5'h0 : _GEN_20899; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_20901 = 5'hb == _T_2088[4:0] ? w_vn_11 : _GEN_20900; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_20902 = 5'hc == _T_2088[4:0] ? w_vn_12 : _GEN_20901; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_20903 = 5'hd == _T_2088[4:0] ? w_vn_13 : _GEN_20902; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_20904 = 5'he == _T_2088[4:0] ? 5'h0 : _GEN_20903; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_20905 = 5'hf == _T_2088[4:0] ? w_vn_15 : _GEN_20904; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_20906 = 5'h10 == _T_2088[4:0] ? w_vn_16 : _GEN_20905; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_20907 = 5'h11 == _T_2088[4:0] ? 5'h0 : _GEN_20906; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_20908 = 5'h12 == _T_2088[4:0] ? w_vn_18 : _GEN_20907; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_20909 = 5'h13 == _T_2088[4:0] ? 5'h0 : _GEN_20908; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_20910 = 5'h14 == _T_2088[4:0] ? 5'h0 : _GEN_20909; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_20911 = 5'h15 == _T_2088[4:0] ? 5'h0 : _GEN_20910; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_20912 = 5'h16 == _T_2088[4:0] ? 5'h0 : _GEN_20911; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_20913 = 5'h17 == _T_2088[4:0] ? w_vn_23 : _GEN_20912; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_20914 = 5'h18 == _T_2088[4:0] ? w_vn_24 : _GEN_20913; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_20915 = 5'h19 == _T_2088[4:0] ? 5'h0 : _GEN_20914; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_20916 = 5'h1a == _T_2088[4:0] ? 5'h0 : _GEN_20915; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_20917 = 5'h1b == _T_2088[4:0] ? 5'h0 : _GEN_20916; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_20918 = 5'h1c == _T_2088[4:0] ? 5'h0 : _GEN_20917; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_20919 = 5'h1d == _T_2088[4:0] ? 5'h0 : _GEN_20918; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_20920 = 5'h1e == _T_2088[4:0] ? 5'h0 : _GEN_20919; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_20921 = 5'h1f == _T_2088[4:0] ? 5'h0 : _GEN_20920; // @[FanCtrl.scala 54:{41,41}]
  wire  _T_2090 = _GEN_20764 != _GEN_20921; // @[FanCtrl.scala 54:41]
  wire  _T_2099 = _GEN_20732 != _GEN_20764; // @[FanCtrl.scala 56:41]
  wire  _T_2109 = _GEN_20764 == _GEN_20921; // @[FanCtrl.scala 61:48]
  wire  _GEN_21158 = r_valid_1 & _T_2077; // @[FanCtrl.scala 47:34]
  wire [5:0] _T_2145 = _T_2069 - 6'h1; // @[FanCtrl.scala 94:58]
  wire [4:0] _GEN_21402 = 5'h3 == _T_2145[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_21403 = 5'h4 == _T_2145[4:0] ? w_vn_4 : _GEN_21402; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_21404 = 5'h5 == _T_2145[4:0] ? 5'h0 : _GEN_21403; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_21405 = 5'h6 == _T_2145[4:0] ? 5'h0 : _GEN_21404; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_21406 = 5'h7 == _T_2145[4:0] ? w_vn_7 : _GEN_21405; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_21407 = 5'h8 == _T_2145[4:0] ? w_vn_8 : _GEN_21406; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_21408 = 5'h9 == _T_2145[4:0] ? 5'h0 : _GEN_21407; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_21409 = 5'ha == _T_2145[4:0] ? 5'h0 : _GEN_21408; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_21410 = 5'hb == _T_2145[4:0] ? w_vn_11 : _GEN_21409; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_21411 = 5'hc == _T_2145[4:0] ? w_vn_12 : _GEN_21410; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_21412 = 5'hd == _T_2145[4:0] ? w_vn_13 : _GEN_21411; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_21413 = 5'he == _T_2145[4:0] ? 5'h0 : _GEN_21412; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_21414 = 5'hf == _T_2145[4:0] ? w_vn_15 : _GEN_21413; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_21415 = 5'h10 == _T_2145[4:0] ? w_vn_16 : _GEN_21414; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_21416 = 5'h11 == _T_2145[4:0] ? 5'h0 : _GEN_21415; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_21417 = 5'h12 == _T_2145[4:0] ? w_vn_18 : _GEN_21416; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_21418 = 5'h13 == _T_2145[4:0] ? 5'h0 : _GEN_21417; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_21419 = 5'h14 == _T_2145[4:0] ? 5'h0 : _GEN_21418; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_21420 = 5'h15 == _T_2145[4:0] ? 5'h0 : _GEN_21419; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_21421 = 5'h16 == _T_2145[4:0] ? 5'h0 : _GEN_21420; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_21422 = 5'h17 == _T_2145[4:0] ? w_vn_23 : _GEN_21421; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_21423 = 5'h18 == _T_2145[4:0] ? w_vn_24 : _GEN_21422; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_21424 = 5'h19 == _T_2145[4:0] ? 5'h0 : _GEN_21423; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_21425 = 5'h1a == _T_2145[4:0] ? 5'h0 : _GEN_21424; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_21426 = 5'h1b == _T_2145[4:0] ? 5'h0 : _GEN_21425; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_21427 = 5'h1c == _T_2145[4:0] ? 5'h0 : _GEN_21426; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_21428 = 5'h1d == _T_2145[4:0] ? 5'h0 : _GEN_21427; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_21429 = 5'h1e == _T_2145[4:0] ? 5'h0 : _GEN_21428; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_21430 = 5'h1f == _T_2145[4:0] ? 5'h0 : _GEN_21429; // @[FanCtrl.scala 94:{39,39}]
  wire  _T_2147 = _GEN_20732 != _GEN_21430; // @[FanCtrl.scala 94:39]
  wire  _T_2166 = _GEN_20732 == _GEN_21430; // @[FanCtrl.scala 99:46]
  wire  _T_2213 = _T_2147 & _T_2090; // @[FanCtrl.scala 125:65]
  wire  _T_2223 = _T_2213 & _T_2099; // @[FanCtrl.scala 126:65]
  wire  _T_2242 = _T_2166 & _T_2090; // @[FanCtrl.scala 131:70]
  wire  _T_2252 = _T_2242 & _T_2099; // @[FanCtrl.scala 132:72]
  wire  _T_2271 = _T_2147 & _T_2109; // @[FanCtrl.scala 137:72]
  wire  _T_2281 = _T_2271 & _T_2099; // @[FanCtrl.scala 138:71]
  wire [1:0] _GEN_22452 = _T_2281 ? 2'h3 : 2'h1; // @[FanCtrl.scala 139:73 141:34 144:35]
  wire [2:0] _GEN_22453 = _T_2252 ? 3'h4 : {{1'd0}, _GEN_22452}; // @[FanCtrl.scala 133:73 135:35]
  wire [2:0] _GEN_22454 = _T_2223 ? 3'h5 : _GEN_22453; // @[FanCtrl.scala 127:66 129:35]
  wire [2:0] _GEN_22517 = r_valid_1 ? _GEN_22454 : 3'h0; // @[FanCtrl.scala 117:32 148:33]
  wire [5:0] _T_2286 = 2'h2 * 4'hc; // @[FanCtrl.scala 48:25]
  wire [6:0] _T_2287 = {{1'd0}, _T_2286}; // @[FanCtrl.scala 48:31]
  wire [5:0] _T_2292 = _T_2286 + 6'h1; // @[FanCtrl.scala 48:58]
  wire [4:0] _GEN_22586 = 5'h3 == _T_2287[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_22587 = 5'h4 == _T_2287[4:0] ? w_vn_4 : _GEN_22586; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_22588 = 5'h5 == _T_2287[4:0] ? 5'h0 : _GEN_22587; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_22589 = 5'h6 == _T_2287[4:0] ? 5'h0 : _GEN_22588; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_22590 = 5'h7 == _T_2287[4:0] ? w_vn_7 : _GEN_22589; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_22591 = 5'h8 == _T_2287[4:0] ? w_vn_8 : _GEN_22590; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_22592 = 5'h9 == _T_2287[4:0] ? 5'h0 : _GEN_22591; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_22593 = 5'ha == _T_2287[4:0] ? 5'h0 : _GEN_22592; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_22594 = 5'hb == _T_2287[4:0] ? w_vn_11 : _GEN_22593; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_22595 = 5'hc == _T_2287[4:0] ? w_vn_12 : _GEN_22594; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_22596 = 5'hd == _T_2287[4:0] ? w_vn_13 : _GEN_22595; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_22597 = 5'he == _T_2287[4:0] ? 5'h0 : _GEN_22596; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_22598 = 5'hf == _T_2287[4:0] ? w_vn_15 : _GEN_22597; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_22599 = 5'h10 == _T_2287[4:0] ? w_vn_16 : _GEN_22598; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_22600 = 5'h11 == _T_2287[4:0] ? 5'h0 : _GEN_22599; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_22601 = 5'h12 == _T_2287[4:0] ? w_vn_18 : _GEN_22600; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_22602 = 5'h13 == _T_2287[4:0] ? 5'h0 : _GEN_22601; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_22603 = 5'h14 == _T_2287[4:0] ? 5'h0 : _GEN_22602; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_22604 = 5'h15 == _T_2287[4:0] ? 5'h0 : _GEN_22603; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_22605 = 5'h16 == _T_2287[4:0] ? 5'h0 : _GEN_22604; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_22606 = 5'h17 == _T_2287[4:0] ? w_vn_23 : _GEN_22605; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_22607 = 5'h18 == _T_2287[4:0] ? w_vn_24 : _GEN_22606; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_22608 = 5'h19 == _T_2287[4:0] ? 5'h0 : _GEN_22607; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_22609 = 5'h1a == _T_2287[4:0] ? 5'h0 : _GEN_22608; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_22610 = 5'h1b == _T_2287[4:0] ? 5'h0 : _GEN_22609; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_22611 = 5'h1c == _T_2287[4:0] ? 5'h0 : _GEN_22610; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_22612 = 5'h1d == _T_2287[4:0] ? 5'h0 : _GEN_22611; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_22613 = 5'h1e == _T_2287[4:0] ? 5'h0 : _GEN_22612; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_22614 = 5'h1f == _T_2287[4:0] ? 5'h0 : _GEN_22613; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_22618 = 5'h3 == _T_2292[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_22619 = 5'h4 == _T_2292[4:0] ? w_vn_4 : _GEN_22618; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_22620 = 5'h5 == _T_2292[4:0] ? 5'h0 : _GEN_22619; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_22621 = 5'h6 == _T_2292[4:0] ? 5'h0 : _GEN_22620; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_22622 = 5'h7 == _T_2292[4:0] ? w_vn_7 : _GEN_22621; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_22623 = 5'h8 == _T_2292[4:0] ? w_vn_8 : _GEN_22622; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_22624 = 5'h9 == _T_2292[4:0] ? 5'h0 : _GEN_22623; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_22625 = 5'ha == _T_2292[4:0] ? 5'h0 : _GEN_22624; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_22626 = 5'hb == _T_2292[4:0] ? w_vn_11 : _GEN_22625; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_22627 = 5'hc == _T_2292[4:0] ? w_vn_12 : _GEN_22626; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_22628 = 5'hd == _T_2292[4:0] ? w_vn_13 : _GEN_22627; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_22629 = 5'he == _T_2292[4:0] ? 5'h0 : _GEN_22628; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_22630 = 5'hf == _T_2292[4:0] ? w_vn_15 : _GEN_22629; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_22631 = 5'h10 == _T_2292[4:0] ? w_vn_16 : _GEN_22630; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_22632 = 5'h11 == _T_2292[4:0] ? 5'h0 : _GEN_22631; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_22633 = 5'h12 == _T_2292[4:0] ? w_vn_18 : _GEN_22632; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_22634 = 5'h13 == _T_2292[4:0] ? 5'h0 : _GEN_22633; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_22635 = 5'h14 == _T_2292[4:0] ? 5'h0 : _GEN_22634; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_22636 = 5'h15 == _T_2292[4:0] ? 5'h0 : _GEN_22635; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_22637 = 5'h16 == _T_2292[4:0] ? 5'h0 : _GEN_22636; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_22638 = 5'h17 == _T_2292[4:0] ? w_vn_23 : _GEN_22637; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_22639 = 5'h18 == _T_2292[4:0] ? w_vn_24 : _GEN_22638; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_22640 = 5'h19 == _T_2292[4:0] ? 5'h0 : _GEN_22639; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_22641 = 5'h1a == _T_2292[4:0] ? 5'h0 : _GEN_22640; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_22642 = 5'h1b == _T_2292[4:0] ? 5'h0 : _GEN_22641; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_22643 = 5'h1c == _T_2292[4:0] ? 5'h0 : _GEN_22642; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_22644 = 5'h1d == _T_2292[4:0] ? 5'h0 : _GEN_22643; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_22645 = 5'h1e == _T_2292[4:0] ? 5'h0 : _GEN_22644; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_22646 = 5'h1f == _T_2292[4:0] ? 5'h0 : _GEN_22645; // @[FanCtrl.scala 48:{39,39}]
  wire  _T_2294 = _GEN_22614 == _GEN_22646; // @[FanCtrl.scala 48:39]
  wire [5:0] _T_2305 = _T_2286 + 6'h2; // @[FanCtrl.scala 55:32]
  wire [4:0] _GEN_22775 = 5'h3 == _T_2305[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_22776 = 5'h4 == _T_2305[4:0] ? w_vn_4 : _GEN_22775; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_22777 = 5'h5 == _T_2305[4:0] ? 5'h0 : _GEN_22776; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_22778 = 5'h6 == _T_2305[4:0] ? 5'h0 : _GEN_22777; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_22779 = 5'h7 == _T_2305[4:0] ? w_vn_7 : _GEN_22778; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_22780 = 5'h8 == _T_2305[4:0] ? w_vn_8 : _GEN_22779; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_22781 = 5'h9 == _T_2305[4:0] ? 5'h0 : _GEN_22780; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_22782 = 5'ha == _T_2305[4:0] ? 5'h0 : _GEN_22781; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_22783 = 5'hb == _T_2305[4:0] ? w_vn_11 : _GEN_22782; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_22784 = 5'hc == _T_2305[4:0] ? w_vn_12 : _GEN_22783; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_22785 = 5'hd == _T_2305[4:0] ? w_vn_13 : _GEN_22784; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_22786 = 5'he == _T_2305[4:0] ? 5'h0 : _GEN_22785; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_22787 = 5'hf == _T_2305[4:0] ? w_vn_15 : _GEN_22786; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_22788 = 5'h10 == _T_2305[4:0] ? w_vn_16 : _GEN_22787; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_22789 = 5'h11 == _T_2305[4:0] ? 5'h0 : _GEN_22788; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_22790 = 5'h12 == _T_2305[4:0] ? w_vn_18 : _GEN_22789; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_22791 = 5'h13 == _T_2305[4:0] ? 5'h0 : _GEN_22790; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_22792 = 5'h14 == _T_2305[4:0] ? 5'h0 : _GEN_22791; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_22793 = 5'h15 == _T_2305[4:0] ? 5'h0 : _GEN_22792; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_22794 = 5'h16 == _T_2305[4:0] ? 5'h0 : _GEN_22793; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_22795 = 5'h17 == _T_2305[4:0] ? w_vn_23 : _GEN_22794; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_22796 = 5'h18 == _T_2305[4:0] ? w_vn_24 : _GEN_22795; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_22797 = 5'h19 == _T_2305[4:0] ? 5'h0 : _GEN_22796; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_22798 = 5'h1a == _T_2305[4:0] ? 5'h0 : _GEN_22797; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_22799 = 5'h1b == _T_2305[4:0] ? 5'h0 : _GEN_22798; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_22800 = 5'h1c == _T_2305[4:0] ? 5'h0 : _GEN_22799; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_22801 = 5'h1d == _T_2305[4:0] ? 5'h0 : _GEN_22800; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_22802 = 5'h1e == _T_2305[4:0] ? 5'h0 : _GEN_22801; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_22803 = 5'h1f == _T_2305[4:0] ? 5'h0 : _GEN_22802; // @[FanCtrl.scala 54:{41,41}]
  wire  _T_2307 = _GEN_22646 != _GEN_22803; // @[FanCtrl.scala 54:41]
  wire  _T_2316 = _GEN_22614 != _GEN_22646; // @[FanCtrl.scala 56:41]
  wire  _T_2326 = _GEN_22646 == _GEN_22803; // @[FanCtrl.scala 61:48]
  wire  _GEN_23041 = r_valid_1 & _T_2294; // @[FanCtrl.scala 47:34]
  wire [5:0] _T_2362 = _T_2286 - 6'h1; // @[FanCtrl.scala 94:58]
  wire [4:0] _GEN_23284 = 5'h3 == _T_2362[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_23285 = 5'h4 == _T_2362[4:0] ? w_vn_4 : _GEN_23284; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_23286 = 5'h5 == _T_2362[4:0] ? 5'h0 : _GEN_23285; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_23287 = 5'h6 == _T_2362[4:0] ? 5'h0 : _GEN_23286; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_23288 = 5'h7 == _T_2362[4:0] ? w_vn_7 : _GEN_23287; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_23289 = 5'h8 == _T_2362[4:0] ? w_vn_8 : _GEN_23288; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_23290 = 5'h9 == _T_2362[4:0] ? 5'h0 : _GEN_23289; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_23291 = 5'ha == _T_2362[4:0] ? 5'h0 : _GEN_23290; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_23292 = 5'hb == _T_2362[4:0] ? w_vn_11 : _GEN_23291; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_23293 = 5'hc == _T_2362[4:0] ? w_vn_12 : _GEN_23292; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_23294 = 5'hd == _T_2362[4:0] ? w_vn_13 : _GEN_23293; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_23295 = 5'he == _T_2362[4:0] ? 5'h0 : _GEN_23294; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_23296 = 5'hf == _T_2362[4:0] ? w_vn_15 : _GEN_23295; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_23297 = 5'h10 == _T_2362[4:0] ? w_vn_16 : _GEN_23296; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_23298 = 5'h11 == _T_2362[4:0] ? 5'h0 : _GEN_23297; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_23299 = 5'h12 == _T_2362[4:0] ? w_vn_18 : _GEN_23298; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_23300 = 5'h13 == _T_2362[4:0] ? 5'h0 : _GEN_23299; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_23301 = 5'h14 == _T_2362[4:0] ? 5'h0 : _GEN_23300; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_23302 = 5'h15 == _T_2362[4:0] ? 5'h0 : _GEN_23301; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_23303 = 5'h16 == _T_2362[4:0] ? 5'h0 : _GEN_23302; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_23304 = 5'h17 == _T_2362[4:0] ? w_vn_23 : _GEN_23303; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_23305 = 5'h18 == _T_2362[4:0] ? w_vn_24 : _GEN_23304; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_23306 = 5'h19 == _T_2362[4:0] ? 5'h0 : _GEN_23305; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_23307 = 5'h1a == _T_2362[4:0] ? 5'h0 : _GEN_23306; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_23308 = 5'h1b == _T_2362[4:0] ? 5'h0 : _GEN_23307; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_23309 = 5'h1c == _T_2362[4:0] ? 5'h0 : _GEN_23308; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_23310 = 5'h1d == _T_2362[4:0] ? 5'h0 : _GEN_23309; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_23311 = 5'h1e == _T_2362[4:0] ? 5'h0 : _GEN_23310; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_23312 = 5'h1f == _T_2362[4:0] ? 5'h0 : _GEN_23311; // @[FanCtrl.scala 94:{39,39}]
  wire  _T_2364 = _GEN_22614 != _GEN_23312; // @[FanCtrl.scala 94:39]
  wire  _T_2383 = _GEN_22614 == _GEN_23312; // @[FanCtrl.scala 99:46]
  wire  _T_2430 = _T_2364 & _T_2307; // @[FanCtrl.scala 125:65]
  wire  _T_2440 = _T_2430 & _T_2316; // @[FanCtrl.scala 126:65]
  wire  _T_2459 = _T_2383 & _T_2307; // @[FanCtrl.scala 131:70]
  wire  _T_2469 = _T_2459 & _T_2316; // @[FanCtrl.scala 132:72]
  wire  _T_2488 = _T_2364 & _T_2326; // @[FanCtrl.scala 137:72]
  wire  _T_2498 = _T_2488 & _T_2316; // @[FanCtrl.scala 138:71]
  wire [1:0] _GEN_24334 = _T_2498 ? 2'h3 : 2'h1; // @[FanCtrl.scala 139:73 141:34 144:35]
  wire [2:0] _GEN_24335 = _T_2469 ? 3'h4 : {{1'd0}, _GEN_24334}; // @[FanCtrl.scala 133:73 135:35]
  wire [2:0] _GEN_24336 = _T_2440 ? 3'h5 : _GEN_24335; // @[FanCtrl.scala 127:66 129:35]
  wire [2:0] _GEN_24399 = r_valid_1 ? _GEN_24336 : 3'h0; // @[FanCtrl.scala 117:32 148:33]
  wire [5:0] _T_2503 = 2'h2 * 4'hd; // @[FanCtrl.scala 48:25]
  wire [6:0] _T_2504 = {{1'd0}, _T_2503}; // @[FanCtrl.scala 48:31]
  wire [5:0] _T_2509 = _T_2503 + 6'h1; // @[FanCtrl.scala 48:58]
  wire [4:0] _GEN_24468 = 5'h3 == _T_2504[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_24469 = 5'h4 == _T_2504[4:0] ? w_vn_4 : _GEN_24468; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_24470 = 5'h5 == _T_2504[4:0] ? 5'h0 : _GEN_24469; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_24471 = 5'h6 == _T_2504[4:0] ? 5'h0 : _GEN_24470; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_24472 = 5'h7 == _T_2504[4:0] ? w_vn_7 : _GEN_24471; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_24473 = 5'h8 == _T_2504[4:0] ? w_vn_8 : _GEN_24472; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_24474 = 5'h9 == _T_2504[4:0] ? 5'h0 : _GEN_24473; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_24475 = 5'ha == _T_2504[4:0] ? 5'h0 : _GEN_24474; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_24476 = 5'hb == _T_2504[4:0] ? w_vn_11 : _GEN_24475; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_24477 = 5'hc == _T_2504[4:0] ? w_vn_12 : _GEN_24476; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_24478 = 5'hd == _T_2504[4:0] ? w_vn_13 : _GEN_24477; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_24479 = 5'he == _T_2504[4:0] ? 5'h0 : _GEN_24478; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_24480 = 5'hf == _T_2504[4:0] ? w_vn_15 : _GEN_24479; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_24481 = 5'h10 == _T_2504[4:0] ? w_vn_16 : _GEN_24480; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_24482 = 5'h11 == _T_2504[4:0] ? 5'h0 : _GEN_24481; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_24483 = 5'h12 == _T_2504[4:0] ? w_vn_18 : _GEN_24482; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_24484 = 5'h13 == _T_2504[4:0] ? 5'h0 : _GEN_24483; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_24485 = 5'h14 == _T_2504[4:0] ? 5'h0 : _GEN_24484; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_24486 = 5'h15 == _T_2504[4:0] ? 5'h0 : _GEN_24485; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_24487 = 5'h16 == _T_2504[4:0] ? 5'h0 : _GEN_24486; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_24488 = 5'h17 == _T_2504[4:0] ? w_vn_23 : _GEN_24487; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_24489 = 5'h18 == _T_2504[4:0] ? w_vn_24 : _GEN_24488; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_24490 = 5'h19 == _T_2504[4:0] ? 5'h0 : _GEN_24489; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_24491 = 5'h1a == _T_2504[4:0] ? 5'h0 : _GEN_24490; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_24492 = 5'h1b == _T_2504[4:0] ? 5'h0 : _GEN_24491; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_24493 = 5'h1c == _T_2504[4:0] ? 5'h0 : _GEN_24492; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_24494 = 5'h1d == _T_2504[4:0] ? 5'h0 : _GEN_24493; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_24495 = 5'h1e == _T_2504[4:0] ? 5'h0 : _GEN_24494; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_24496 = 5'h1f == _T_2504[4:0] ? 5'h0 : _GEN_24495; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_24500 = 5'h3 == _T_2509[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_24501 = 5'h4 == _T_2509[4:0] ? w_vn_4 : _GEN_24500; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_24502 = 5'h5 == _T_2509[4:0] ? 5'h0 : _GEN_24501; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_24503 = 5'h6 == _T_2509[4:0] ? 5'h0 : _GEN_24502; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_24504 = 5'h7 == _T_2509[4:0] ? w_vn_7 : _GEN_24503; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_24505 = 5'h8 == _T_2509[4:0] ? w_vn_8 : _GEN_24504; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_24506 = 5'h9 == _T_2509[4:0] ? 5'h0 : _GEN_24505; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_24507 = 5'ha == _T_2509[4:0] ? 5'h0 : _GEN_24506; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_24508 = 5'hb == _T_2509[4:0] ? w_vn_11 : _GEN_24507; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_24509 = 5'hc == _T_2509[4:0] ? w_vn_12 : _GEN_24508; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_24510 = 5'hd == _T_2509[4:0] ? w_vn_13 : _GEN_24509; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_24511 = 5'he == _T_2509[4:0] ? 5'h0 : _GEN_24510; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_24512 = 5'hf == _T_2509[4:0] ? w_vn_15 : _GEN_24511; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_24513 = 5'h10 == _T_2509[4:0] ? w_vn_16 : _GEN_24512; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_24514 = 5'h11 == _T_2509[4:0] ? 5'h0 : _GEN_24513; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_24515 = 5'h12 == _T_2509[4:0] ? w_vn_18 : _GEN_24514; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_24516 = 5'h13 == _T_2509[4:0] ? 5'h0 : _GEN_24515; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_24517 = 5'h14 == _T_2509[4:0] ? 5'h0 : _GEN_24516; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_24518 = 5'h15 == _T_2509[4:0] ? 5'h0 : _GEN_24517; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_24519 = 5'h16 == _T_2509[4:0] ? 5'h0 : _GEN_24518; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_24520 = 5'h17 == _T_2509[4:0] ? w_vn_23 : _GEN_24519; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_24521 = 5'h18 == _T_2509[4:0] ? w_vn_24 : _GEN_24520; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_24522 = 5'h19 == _T_2509[4:0] ? 5'h0 : _GEN_24521; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_24523 = 5'h1a == _T_2509[4:0] ? 5'h0 : _GEN_24522; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_24524 = 5'h1b == _T_2509[4:0] ? 5'h0 : _GEN_24523; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_24525 = 5'h1c == _T_2509[4:0] ? 5'h0 : _GEN_24524; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_24526 = 5'h1d == _T_2509[4:0] ? 5'h0 : _GEN_24525; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_24527 = 5'h1e == _T_2509[4:0] ? 5'h0 : _GEN_24526; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_24528 = 5'h1f == _T_2509[4:0] ? 5'h0 : _GEN_24527; // @[FanCtrl.scala 48:{39,39}]
  wire  _T_2511 = _GEN_24496 == _GEN_24528; // @[FanCtrl.scala 48:39]
  wire [5:0] _T_2522 = _T_2503 + 6'h2; // @[FanCtrl.scala 55:32]
  wire [4:0] _GEN_24657 = 5'h3 == _T_2522[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_24658 = 5'h4 == _T_2522[4:0] ? w_vn_4 : _GEN_24657; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_24659 = 5'h5 == _T_2522[4:0] ? 5'h0 : _GEN_24658; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_24660 = 5'h6 == _T_2522[4:0] ? 5'h0 : _GEN_24659; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_24661 = 5'h7 == _T_2522[4:0] ? w_vn_7 : _GEN_24660; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_24662 = 5'h8 == _T_2522[4:0] ? w_vn_8 : _GEN_24661; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_24663 = 5'h9 == _T_2522[4:0] ? 5'h0 : _GEN_24662; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_24664 = 5'ha == _T_2522[4:0] ? 5'h0 : _GEN_24663; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_24665 = 5'hb == _T_2522[4:0] ? w_vn_11 : _GEN_24664; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_24666 = 5'hc == _T_2522[4:0] ? w_vn_12 : _GEN_24665; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_24667 = 5'hd == _T_2522[4:0] ? w_vn_13 : _GEN_24666; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_24668 = 5'he == _T_2522[4:0] ? 5'h0 : _GEN_24667; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_24669 = 5'hf == _T_2522[4:0] ? w_vn_15 : _GEN_24668; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_24670 = 5'h10 == _T_2522[4:0] ? w_vn_16 : _GEN_24669; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_24671 = 5'h11 == _T_2522[4:0] ? 5'h0 : _GEN_24670; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_24672 = 5'h12 == _T_2522[4:0] ? w_vn_18 : _GEN_24671; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_24673 = 5'h13 == _T_2522[4:0] ? 5'h0 : _GEN_24672; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_24674 = 5'h14 == _T_2522[4:0] ? 5'h0 : _GEN_24673; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_24675 = 5'h15 == _T_2522[4:0] ? 5'h0 : _GEN_24674; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_24676 = 5'h16 == _T_2522[4:0] ? 5'h0 : _GEN_24675; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_24677 = 5'h17 == _T_2522[4:0] ? w_vn_23 : _GEN_24676; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_24678 = 5'h18 == _T_2522[4:0] ? w_vn_24 : _GEN_24677; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_24679 = 5'h19 == _T_2522[4:0] ? 5'h0 : _GEN_24678; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_24680 = 5'h1a == _T_2522[4:0] ? 5'h0 : _GEN_24679; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_24681 = 5'h1b == _T_2522[4:0] ? 5'h0 : _GEN_24680; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_24682 = 5'h1c == _T_2522[4:0] ? 5'h0 : _GEN_24681; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_24683 = 5'h1d == _T_2522[4:0] ? 5'h0 : _GEN_24682; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_24684 = 5'h1e == _T_2522[4:0] ? 5'h0 : _GEN_24683; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_24685 = 5'h1f == _T_2522[4:0] ? 5'h0 : _GEN_24684; // @[FanCtrl.scala 54:{41,41}]
  wire  _T_2524 = _GEN_24528 != _GEN_24685; // @[FanCtrl.scala 54:41]
  wire  _T_2533 = _GEN_24496 != _GEN_24528; // @[FanCtrl.scala 56:41]
  wire  _T_2543 = _GEN_24528 == _GEN_24685; // @[FanCtrl.scala 61:48]
  wire  _GEN_24924 = r_valid_1 & _T_2511; // @[FanCtrl.scala 47:34]
  wire [5:0] _T_2579 = _T_2503 - 6'h1; // @[FanCtrl.scala 94:58]
  wire [4:0] _GEN_25166 = 5'h3 == _T_2579[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_25167 = 5'h4 == _T_2579[4:0] ? w_vn_4 : _GEN_25166; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_25168 = 5'h5 == _T_2579[4:0] ? 5'h0 : _GEN_25167; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_25169 = 5'h6 == _T_2579[4:0] ? 5'h0 : _GEN_25168; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_25170 = 5'h7 == _T_2579[4:0] ? w_vn_7 : _GEN_25169; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_25171 = 5'h8 == _T_2579[4:0] ? w_vn_8 : _GEN_25170; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_25172 = 5'h9 == _T_2579[4:0] ? 5'h0 : _GEN_25171; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_25173 = 5'ha == _T_2579[4:0] ? 5'h0 : _GEN_25172; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_25174 = 5'hb == _T_2579[4:0] ? w_vn_11 : _GEN_25173; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_25175 = 5'hc == _T_2579[4:0] ? w_vn_12 : _GEN_25174; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_25176 = 5'hd == _T_2579[4:0] ? w_vn_13 : _GEN_25175; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_25177 = 5'he == _T_2579[4:0] ? 5'h0 : _GEN_25176; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_25178 = 5'hf == _T_2579[4:0] ? w_vn_15 : _GEN_25177; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_25179 = 5'h10 == _T_2579[4:0] ? w_vn_16 : _GEN_25178; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_25180 = 5'h11 == _T_2579[4:0] ? 5'h0 : _GEN_25179; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_25181 = 5'h12 == _T_2579[4:0] ? w_vn_18 : _GEN_25180; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_25182 = 5'h13 == _T_2579[4:0] ? 5'h0 : _GEN_25181; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_25183 = 5'h14 == _T_2579[4:0] ? 5'h0 : _GEN_25182; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_25184 = 5'h15 == _T_2579[4:0] ? 5'h0 : _GEN_25183; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_25185 = 5'h16 == _T_2579[4:0] ? 5'h0 : _GEN_25184; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_25186 = 5'h17 == _T_2579[4:0] ? w_vn_23 : _GEN_25185; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_25187 = 5'h18 == _T_2579[4:0] ? w_vn_24 : _GEN_25186; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_25188 = 5'h19 == _T_2579[4:0] ? 5'h0 : _GEN_25187; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_25189 = 5'h1a == _T_2579[4:0] ? 5'h0 : _GEN_25188; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_25190 = 5'h1b == _T_2579[4:0] ? 5'h0 : _GEN_25189; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_25191 = 5'h1c == _T_2579[4:0] ? 5'h0 : _GEN_25190; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_25192 = 5'h1d == _T_2579[4:0] ? 5'h0 : _GEN_25191; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_25193 = 5'h1e == _T_2579[4:0] ? 5'h0 : _GEN_25192; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_25194 = 5'h1f == _T_2579[4:0] ? 5'h0 : _GEN_25193; // @[FanCtrl.scala 94:{39,39}]
  wire  _T_2581 = _GEN_24496 != _GEN_25194; // @[FanCtrl.scala 94:39]
  wire  _T_2600 = _GEN_24496 == _GEN_25194; // @[FanCtrl.scala 99:46]
  wire  _T_2647 = _T_2581 & _T_2524; // @[FanCtrl.scala 125:65]
  wire  _T_2657 = _T_2647 & _T_2533; // @[FanCtrl.scala 126:65]
  wire  _T_2676 = _T_2600 & _T_2524; // @[FanCtrl.scala 131:70]
  wire  _T_2686 = _T_2676 & _T_2533; // @[FanCtrl.scala 132:72]
  wire  _T_2705 = _T_2581 & _T_2543; // @[FanCtrl.scala 137:72]
  wire  _T_2715 = _T_2705 & _T_2533; // @[FanCtrl.scala 138:71]
  wire [1:0] _GEN_26216 = _T_2715 ? 2'h3 : 2'h1; // @[FanCtrl.scala 139:73 141:34 144:35]
  wire [2:0] _GEN_26217 = _T_2686 ? 3'h4 : {{1'd0}, _GEN_26216}; // @[FanCtrl.scala 133:73 135:35]
  wire [2:0] _GEN_26218 = _T_2657 ? 3'h5 : _GEN_26217; // @[FanCtrl.scala 127:66 129:35]
  wire [2:0] _GEN_26281 = r_valid_1 ? _GEN_26218 : 3'h0; // @[FanCtrl.scala 117:32 148:33]
  wire [5:0] _T_2720 = 2'h2 * 4'he; // @[FanCtrl.scala 48:25]
  wire [6:0] _T_2721 = {{1'd0}, _T_2720}; // @[FanCtrl.scala 48:31]
  wire [5:0] _T_2726 = _T_2720 + 6'h1; // @[FanCtrl.scala 48:58]
  wire [4:0] _GEN_26350 = 5'h3 == _T_2721[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_26351 = 5'h4 == _T_2721[4:0] ? w_vn_4 : _GEN_26350; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_26352 = 5'h5 == _T_2721[4:0] ? 5'h0 : _GEN_26351; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_26353 = 5'h6 == _T_2721[4:0] ? 5'h0 : _GEN_26352; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_26354 = 5'h7 == _T_2721[4:0] ? w_vn_7 : _GEN_26353; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_26355 = 5'h8 == _T_2721[4:0] ? w_vn_8 : _GEN_26354; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_26356 = 5'h9 == _T_2721[4:0] ? 5'h0 : _GEN_26355; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_26357 = 5'ha == _T_2721[4:0] ? 5'h0 : _GEN_26356; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_26358 = 5'hb == _T_2721[4:0] ? w_vn_11 : _GEN_26357; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_26359 = 5'hc == _T_2721[4:0] ? w_vn_12 : _GEN_26358; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_26360 = 5'hd == _T_2721[4:0] ? w_vn_13 : _GEN_26359; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_26361 = 5'he == _T_2721[4:0] ? 5'h0 : _GEN_26360; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_26362 = 5'hf == _T_2721[4:0] ? w_vn_15 : _GEN_26361; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_26363 = 5'h10 == _T_2721[4:0] ? w_vn_16 : _GEN_26362; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_26364 = 5'h11 == _T_2721[4:0] ? 5'h0 : _GEN_26363; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_26365 = 5'h12 == _T_2721[4:0] ? w_vn_18 : _GEN_26364; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_26366 = 5'h13 == _T_2721[4:0] ? 5'h0 : _GEN_26365; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_26367 = 5'h14 == _T_2721[4:0] ? 5'h0 : _GEN_26366; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_26368 = 5'h15 == _T_2721[4:0] ? 5'h0 : _GEN_26367; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_26369 = 5'h16 == _T_2721[4:0] ? 5'h0 : _GEN_26368; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_26370 = 5'h17 == _T_2721[4:0] ? w_vn_23 : _GEN_26369; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_26371 = 5'h18 == _T_2721[4:0] ? w_vn_24 : _GEN_26370; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_26372 = 5'h19 == _T_2721[4:0] ? 5'h0 : _GEN_26371; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_26373 = 5'h1a == _T_2721[4:0] ? 5'h0 : _GEN_26372; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_26374 = 5'h1b == _T_2721[4:0] ? 5'h0 : _GEN_26373; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_26375 = 5'h1c == _T_2721[4:0] ? 5'h0 : _GEN_26374; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_26376 = 5'h1d == _T_2721[4:0] ? 5'h0 : _GEN_26375; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_26377 = 5'h1e == _T_2721[4:0] ? 5'h0 : _GEN_26376; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_26378 = 5'h1f == _T_2721[4:0] ? 5'h0 : _GEN_26377; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_26382 = 5'h3 == _T_2726[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_26383 = 5'h4 == _T_2726[4:0] ? w_vn_4 : _GEN_26382; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_26384 = 5'h5 == _T_2726[4:0] ? 5'h0 : _GEN_26383; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_26385 = 5'h6 == _T_2726[4:0] ? 5'h0 : _GEN_26384; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_26386 = 5'h7 == _T_2726[4:0] ? w_vn_7 : _GEN_26385; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_26387 = 5'h8 == _T_2726[4:0] ? w_vn_8 : _GEN_26386; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_26388 = 5'h9 == _T_2726[4:0] ? 5'h0 : _GEN_26387; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_26389 = 5'ha == _T_2726[4:0] ? 5'h0 : _GEN_26388; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_26390 = 5'hb == _T_2726[4:0] ? w_vn_11 : _GEN_26389; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_26391 = 5'hc == _T_2726[4:0] ? w_vn_12 : _GEN_26390; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_26392 = 5'hd == _T_2726[4:0] ? w_vn_13 : _GEN_26391; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_26393 = 5'he == _T_2726[4:0] ? 5'h0 : _GEN_26392; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_26394 = 5'hf == _T_2726[4:0] ? w_vn_15 : _GEN_26393; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_26395 = 5'h10 == _T_2726[4:0] ? w_vn_16 : _GEN_26394; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_26396 = 5'h11 == _T_2726[4:0] ? 5'h0 : _GEN_26395; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_26397 = 5'h12 == _T_2726[4:0] ? w_vn_18 : _GEN_26396; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_26398 = 5'h13 == _T_2726[4:0] ? 5'h0 : _GEN_26397; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_26399 = 5'h14 == _T_2726[4:0] ? 5'h0 : _GEN_26398; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_26400 = 5'h15 == _T_2726[4:0] ? 5'h0 : _GEN_26399; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_26401 = 5'h16 == _T_2726[4:0] ? 5'h0 : _GEN_26400; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_26402 = 5'h17 == _T_2726[4:0] ? w_vn_23 : _GEN_26401; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_26403 = 5'h18 == _T_2726[4:0] ? w_vn_24 : _GEN_26402; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_26404 = 5'h19 == _T_2726[4:0] ? 5'h0 : _GEN_26403; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_26405 = 5'h1a == _T_2726[4:0] ? 5'h0 : _GEN_26404; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_26406 = 5'h1b == _T_2726[4:0] ? 5'h0 : _GEN_26405; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_26407 = 5'h1c == _T_2726[4:0] ? 5'h0 : _GEN_26406; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_26408 = 5'h1d == _T_2726[4:0] ? 5'h0 : _GEN_26407; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_26409 = 5'h1e == _T_2726[4:0] ? 5'h0 : _GEN_26408; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_26410 = 5'h1f == _T_2726[4:0] ? 5'h0 : _GEN_26409; // @[FanCtrl.scala 48:{39,39}]
  wire  _T_2728 = _GEN_26378 == _GEN_26410; // @[FanCtrl.scala 48:39]
  wire [5:0] _T_2739 = _T_2720 + 6'h2; // @[FanCtrl.scala 55:32]
  wire [4:0] _GEN_26539 = 5'h3 == _T_2739[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_26540 = 5'h4 == _T_2739[4:0] ? w_vn_4 : _GEN_26539; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_26541 = 5'h5 == _T_2739[4:0] ? 5'h0 : _GEN_26540; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_26542 = 5'h6 == _T_2739[4:0] ? 5'h0 : _GEN_26541; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_26543 = 5'h7 == _T_2739[4:0] ? w_vn_7 : _GEN_26542; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_26544 = 5'h8 == _T_2739[4:0] ? w_vn_8 : _GEN_26543; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_26545 = 5'h9 == _T_2739[4:0] ? 5'h0 : _GEN_26544; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_26546 = 5'ha == _T_2739[4:0] ? 5'h0 : _GEN_26545; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_26547 = 5'hb == _T_2739[4:0] ? w_vn_11 : _GEN_26546; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_26548 = 5'hc == _T_2739[4:0] ? w_vn_12 : _GEN_26547; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_26549 = 5'hd == _T_2739[4:0] ? w_vn_13 : _GEN_26548; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_26550 = 5'he == _T_2739[4:0] ? 5'h0 : _GEN_26549; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_26551 = 5'hf == _T_2739[4:0] ? w_vn_15 : _GEN_26550; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_26552 = 5'h10 == _T_2739[4:0] ? w_vn_16 : _GEN_26551; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_26553 = 5'h11 == _T_2739[4:0] ? 5'h0 : _GEN_26552; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_26554 = 5'h12 == _T_2739[4:0] ? w_vn_18 : _GEN_26553; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_26555 = 5'h13 == _T_2739[4:0] ? 5'h0 : _GEN_26554; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_26556 = 5'h14 == _T_2739[4:0] ? 5'h0 : _GEN_26555; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_26557 = 5'h15 == _T_2739[4:0] ? 5'h0 : _GEN_26556; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_26558 = 5'h16 == _T_2739[4:0] ? 5'h0 : _GEN_26557; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_26559 = 5'h17 == _T_2739[4:0] ? w_vn_23 : _GEN_26558; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_26560 = 5'h18 == _T_2739[4:0] ? w_vn_24 : _GEN_26559; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_26561 = 5'h19 == _T_2739[4:0] ? 5'h0 : _GEN_26560; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_26562 = 5'h1a == _T_2739[4:0] ? 5'h0 : _GEN_26561; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_26563 = 5'h1b == _T_2739[4:0] ? 5'h0 : _GEN_26562; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_26564 = 5'h1c == _T_2739[4:0] ? 5'h0 : _GEN_26563; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_26565 = 5'h1d == _T_2739[4:0] ? 5'h0 : _GEN_26564; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_26566 = 5'h1e == _T_2739[4:0] ? 5'h0 : _GEN_26565; // @[FanCtrl.scala 54:{41,41}]
  wire [4:0] _GEN_26567 = 5'h1f == _T_2739[4:0] ? 5'h0 : _GEN_26566; // @[FanCtrl.scala 54:{41,41}]
  wire  _T_2741 = _GEN_26410 != _GEN_26567; // @[FanCtrl.scala 54:41]
  wire  _T_2750 = _GEN_26378 != _GEN_26410; // @[FanCtrl.scala 56:41]
  wire  _T_2760 = _GEN_26410 == _GEN_26567; // @[FanCtrl.scala 61:48]
  wire  _GEN_26807 = r_valid_1 & _T_2728; // @[FanCtrl.scala 47:34]
  wire [5:0] _T_2796 = _T_2720 - 6'h1; // @[FanCtrl.scala 94:58]
  wire [4:0] _GEN_27048 = 5'h3 == _T_2796[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_27049 = 5'h4 == _T_2796[4:0] ? w_vn_4 : _GEN_27048; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_27050 = 5'h5 == _T_2796[4:0] ? 5'h0 : _GEN_27049; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_27051 = 5'h6 == _T_2796[4:0] ? 5'h0 : _GEN_27050; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_27052 = 5'h7 == _T_2796[4:0] ? w_vn_7 : _GEN_27051; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_27053 = 5'h8 == _T_2796[4:0] ? w_vn_8 : _GEN_27052; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_27054 = 5'h9 == _T_2796[4:0] ? 5'h0 : _GEN_27053; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_27055 = 5'ha == _T_2796[4:0] ? 5'h0 : _GEN_27054; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_27056 = 5'hb == _T_2796[4:0] ? w_vn_11 : _GEN_27055; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_27057 = 5'hc == _T_2796[4:0] ? w_vn_12 : _GEN_27056; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_27058 = 5'hd == _T_2796[4:0] ? w_vn_13 : _GEN_27057; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_27059 = 5'he == _T_2796[4:0] ? 5'h0 : _GEN_27058; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_27060 = 5'hf == _T_2796[4:0] ? w_vn_15 : _GEN_27059; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_27061 = 5'h10 == _T_2796[4:0] ? w_vn_16 : _GEN_27060; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_27062 = 5'h11 == _T_2796[4:0] ? 5'h0 : _GEN_27061; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_27063 = 5'h12 == _T_2796[4:0] ? w_vn_18 : _GEN_27062; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_27064 = 5'h13 == _T_2796[4:0] ? 5'h0 : _GEN_27063; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_27065 = 5'h14 == _T_2796[4:0] ? 5'h0 : _GEN_27064; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_27066 = 5'h15 == _T_2796[4:0] ? 5'h0 : _GEN_27065; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_27067 = 5'h16 == _T_2796[4:0] ? 5'h0 : _GEN_27066; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_27068 = 5'h17 == _T_2796[4:0] ? w_vn_23 : _GEN_27067; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_27069 = 5'h18 == _T_2796[4:0] ? w_vn_24 : _GEN_27068; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_27070 = 5'h19 == _T_2796[4:0] ? 5'h0 : _GEN_27069; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_27071 = 5'h1a == _T_2796[4:0] ? 5'h0 : _GEN_27070; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_27072 = 5'h1b == _T_2796[4:0] ? 5'h0 : _GEN_27071; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_27073 = 5'h1c == _T_2796[4:0] ? 5'h0 : _GEN_27072; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_27074 = 5'h1d == _T_2796[4:0] ? 5'h0 : _GEN_27073; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_27075 = 5'h1e == _T_2796[4:0] ? 5'h0 : _GEN_27074; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_27076 = 5'h1f == _T_2796[4:0] ? 5'h0 : _GEN_27075; // @[FanCtrl.scala 94:{39,39}]
  wire  _T_2798 = _GEN_26378 != _GEN_27076; // @[FanCtrl.scala 94:39]
  wire  _T_2817 = _GEN_26378 == _GEN_27076; // @[FanCtrl.scala 99:46]
  wire  _T_2864 = _T_2798 & _T_2741; // @[FanCtrl.scala 125:65]
  wire  _T_2874 = _T_2864 & _T_2750; // @[FanCtrl.scala 126:65]
  wire  _T_2893 = _T_2817 & _T_2741; // @[FanCtrl.scala 131:70]
  wire  _T_2903 = _T_2893 & _T_2750; // @[FanCtrl.scala 132:72]
  wire  _T_2922 = _T_2798 & _T_2760; // @[FanCtrl.scala 137:72]
  wire  _T_2932 = _T_2922 & _T_2750; // @[FanCtrl.scala 138:71]
  wire [1:0] _GEN_28098 = _T_2932 ? 2'h3 : 2'h1; // @[FanCtrl.scala 139:73 141:34 144:35]
  wire [2:0] _GEN_28099 = _T_2903 ? 3'h4 : {{1'd0}, _GEN_28098}; // @[FanCtrl.scala 133:73 135:35]
  wire [2:0] _GEN_28100 = _T_2874 ? 3'h5 : _GEN_28099; // @[FanCtrl.scala 127:66 129:35]
  wire [2:0] _GEN_28163 = r_valid_1 ? _GEN_28100 : 3'h0; // @[FanCtrl.scala 117:32 148:33]
  wire [5:0] _T_2937 = 2'h2 * 4'hf; // @[FanCtrl.scala 48:25]
  wire [6:0] _T_2938 = {{1'd0}, _T_2937}; // @[FanCtrl.scala 48:31]
  wire [5:0] _T_2943 = _T_2937 + 6'h1; // @[FanCtrl.scala 48:58]
  wire [4:0] _GEN_28232 = 5'h3 == _T_2938[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_28233 = 5'h4 == _T_2938[4:0] ? w_vn_4 : _GEN_28232; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_28234 = 5'h5 == _T_2938[4:0] ? 5'h0 : _GEN_28233; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_28235 = 5'h6 == _T_2938[4:0] ? 5'h0 : _GEN_28234; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_28236 = 5'h7 == _T_2938[4:0] ? w_vn_7 : _GEN_28235; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_28237 = 5'h8 == _T_2938[4:0] ? w_vn_8 : _GEN_28236; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_28238 = 5'h9 == _T_2938[4:0] ? 5'h0 : _GEN_28237; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_28239 = 5'ha == _T_2938[4:0] ? 5'h0 : _GEN_28238; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_28240 = 5'hb == _T_2938[4:0] ? w_vn_11 : _GEN_28239; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_28241 = 5'hc == _T_2938[4:0] ? w_vn_12 : _GEN_28240; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_28242 = 5'hd == _T_2938[4:0] ? w_vn_13 : _GEN_28241; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_28243 = 5'he == _T_2938[4:0] ? 5'h0 : _GEN_28242; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_28244 = 5'hf == _T_2938[4:0] ? w_vn_15 : _GEN_28243; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_28245 = 5'h10 == _T_2938[4:0] ? w_vn_16 : _GEN_28244; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_28246 = 5'h11 == _T_2938[4:0] ? 5'h0 : _GEN_28245; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_28247 = 5'h12 == _T_2938[4:0] ? w_vn_18 : _GEN_28246; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_28248 = 5'h13 == _T_2938[4:0] ? 5'h0 : _GEN_28247; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_28249 = 5'h14 == _T_2938[4:0] ? 5'h0 : _GEN_28248; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_28250 = 5'h15 == _T_2938[4:0] ? 5'h0 : _GEN_28249; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_28251 = 5'h16 == _T_2938[4:0] ? 5'h0 : _GEN_28250; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_28252 = 5'h17 == _T_2938[4:0] ? w_vn_23 : _GEN_28251; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_28253 = 5'h18 == _T_2938[4:0] ? w_vn_24 : _GEN_28252; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_28254 = 5'h19 == _T_2938[4:0] ? 5'h0 : _GEN_28253; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_28255 = 5'h1a == _T_2938[4:0] ? 5'h0 : _GEN_28254; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_28256 = 5'h1b == _T_2938[4:0] ? 5'h0 : _GEN_28255; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_28257 = 5'h1c == _T_2938[4:0] ? 5'h0 : _GEN_28256; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_28258 = 5'h1d == _T_2938[4:0] ? 5'h0 : _GEN_28257; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_28259 = 5'h1e == _T_2938[4:0] ? 5'h0 : _GEN_28258; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_28260 = 5'h1f == _T_2938[4:0] ? 5'h0 : _GEN_28259; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_28264 = 5'h3 == _T_2943[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_28265 = 5'h4 == _T_2943[4:0] ? w_vn_4 : _GEN_28264; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_28266 = 5'h5 == _T_2943[4:0] ? 5'h0 : _GEN_28265; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_28267 = 5'h6 == _T_2943[4:0] ? 5'h0 : _GEN_28266; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_28268 = 5'h7 == _T_2943[4:0] ? w_vn_7 : _GEN_28267; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_28269 = 5'h8 == _T_2943[4:0] ? w_vn_8 : _GEN_28268; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_28270 = 5'h9 == _T_2943[4:0] ? 5'h0 : _GEN_28269; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_28271 = 5'ha == _T_2943[4:0] ? 5'h0 : _GEN_28270; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_28272 = 5'hb == _T_2943[4:0] ? w_vn_11 : _GEN_28271; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_28273 = 5'hc == _T_2943[4:0] ? w_vn_12 : _GEN_28272; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_28274 = 5'hd == _T_2943[4:0] ? w_vn_13 : _GEN_28273; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_28275 = 5'he == _T_2943[4:0] ? 5'h0 : _GEN_28274; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_28276 = 5'hf == _T_2943[4:0] ? w_vn_15 : _GEN_28275; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_28277 = 5'h10 == _T_2943[4:0] ? w_vn_16 : _GEN_28276; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_28278 = 5'h11 == _T_2943[4:0] ? 5'h0 : _GEN_28277; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_28279 = 5'h12 == _T_2943[4:0] ? w_vn_18 : _GEN_28278; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_28280 = 5'h13 == _T_2943[4:0] ? 5'h0 : _GEN_28279; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_28281 = 5'h14 == _T_2943[4:0] ? 5'h0 : _GEN_28280; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_28282 = 5'h15 == _T_2943[4:0] ? 5'h0 : _GEN_28281; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_28283 = 5'h16 == _T_2943[4:0] ? 5'h0 : _GEN_28282; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_28284 = 5'h17 == _T_2943[4:0] ? w_vn_23 : _GEN_28283; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_28285 = 5'h18 == _T_2943[4:0] ? w_vn_24 : _GEN_28284; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_28286 = 5'h19 == _T_2943[4:0] ? 5'h0 : _GEN_28285; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_28287 = 5'h1a == _T_2943[4:0] ? 5'h0 : _GEN_28286; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_28288 = 5'h1b == _T_2943[4:0] ? 5'h0 : _GEN_28287; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_28289 = 5'h1c == _T_2943[4:0] ? 5'h0 : _GEN_28288; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_28290 = 5'h1d == _T_2943[4:0] ? 5'h0 : _GEN_28289; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_28291 = 5'h1e == _T_2943[4:0] ? 5'h0 : _GEN_28290; // @[FanCtrl.scala 48:{39,39}]
  wire [4:0] _GEN_28292 = 5'h1f == _T_2943[4:0] ? 5'h0 : _GEN_28291; // @[FanCtrl.scala 48:{39,39}]
  wire  _T_2945 = _GEN_28260 == _GEN_28292; // @[FanCtrl.scala 48:39]
  wire  _T_2967 = _GEN_28260 != _GEN_28292; // @[FanCtrl.scala 56:41]
  wire  _GEN_28690 = r_valid_1 & _T_2945; // @[FanCtrl.scala 47:34]
  wire [5:0] _T_3013 = _T_2937 - 6'h1; // @[FanCtrl.scala 94:58]
  wire [4:0] _GEN_28930 = 5'h3 == _T_3013[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_28931 = 5'h4 == _T_3013[4:0] ? w_vn_4 : _GEN_28930; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_28932 = 5'h5 == _T_3013[4:0] ? 5'h0 : _GEN_28931; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_28933 = 5'h6 == _T_3013[4:0] ? 5'h0 : _GEN_28932; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_28934 = 5'h7 == _T_3013[4:0] ? w_vn_7 : _GEN_28933; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_28935 = 5'h8 == _T_3013[4:0] ? w_vn_8 : _GEN_28934; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_28936 = 5'h9 == _T_3013[4:0] ? 5'h0 : _GEN_28935; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_28937 = 5'ha == _T_3013[4:0] ? 5'h0 : _GEN_28936; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_28938 = 5'hb == _T_3013[4:0] ? w_vn_11 : _GEN_28937; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_28939 = 5'hc == _T_3013[4:0] ? w_vn_12 : _GEN_28938; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_28940 = 5'hd == _T_3013[4:0] ? w_vn_13 : _GEN_28939; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_28941 = 5'he == _T_3013[4:0] ? 5'h0 : _GEN_28940; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_28942 = 5'hf == _T_3013[4:0] ? w_vn_15 : _GEN_28941; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_28943 = 5'h10 == _T_3013[4:0] ? w_vn_16 : _GEN_28942; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_28944 = 5'h11 == _T_3013[4:0] ? 5'h0 : _GEN_28943; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_28945 = 5'h12 == _T_3013[4:0] ? w_vn_18 : _GEN_28944; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_28946 = 5'h13 == _T_3013[4:0] ? 5'h0 : _GEN_28945; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_28947 = 5'h14 == _T_3013[4:0] ? 5'h0 : _GEN_28946; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_28948 = 5'h15 == _T_3013[4:0] ? 5'h0 : _GEN_28947; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_28949 = 5'h16 == _T_3013[4:0] ? 5'h0 : _GEN_28948; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_28950 = 5'h17 == _T_3013[4:0] ? w_vn_23 : _GEN_28949; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_28951 = 5'h18 == _T_3013[4:0] ? w_vn_24 : _GEN_28950; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_28952 = 5'h19 == _T_3013[4:0] ? 5'h0 : _GEN_28951; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_28953 = 5'h1a == _T_3013[4:0] ? 5'h0 : _GEN_28952; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_28954 = 5'h1b == _T_3013[4:0] ? 5'h0 : _GEN_28953; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_28955 = 5'h1c == _T_3013[4:0] ? 5'h0 : _GEN_28954; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_28956 = 5'h1d == _T_3013[4:0] ? 5'h0 : _GEN_28955; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_28957 = 5'h1e == _T_3013[4:0] ? 5'h0 : _GEN_28956; // @[FanCtrl.scala 94:{39,39}]
  wire [4:0] _GEN_28958 = 5'h1f == _T_3013[4:0] ? 5'h0 : _GEN_28957; // @[FanCtrl.scala 94:{39,39}]
  wire  _T_3025 = _GEN_28260 != _GEN_28958 & _T_2967; // @[FanCtrl.scala 94:67]
  wire  _T_3044 = _GEN_28260 == _GEN_28958 & _T_2967; // @[FanCtrl.scala 99:73]
  wire [2:0] _GEN_29151 = _T_3044 ? 3'h4 : 3'h0; // @[FanCtrl.scala 100:66 102:35 105:35]
  wire [2:0] _GEN_29152 = _T_3025 ? 3'h5 : _GEN_29151; // @[FanCtrl.scala 95:66 97:36]
  wire [2:0] _GEN_29215 = r_valid_1 ? _GEN_29152 : 3'h0; // @[FanCtrl.scala 109:33 87:34]
  wire [3:0] _T_3158 = 3'h4 * 1'h0; // @[FanCtrl.scala 160:23]
  wire [3:0] _T_3160 = _T_3158 + 4'h1; // @[FanCtrl.scala 160:29]
  wire [3:0] _T_3163 = _T_3158 + 4'h2; // @[FanCtrl.scala 160:56]
  wire [4:0] _GEN_30176 = 4'h3 == _T_3160 ? w_vn_3 : 5'h0; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_30177 = 4'h4 == _T_3160 ? w_vn_4 : _GEN_30176; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_30178 = 4'h5 == _T_3160 ? 5'h0 : _GEN_30177; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_30179 = 4'h6 == _T_3160 ? 5'h0 : _GEN_30178; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_30180 = 4'h7 == _T_3160 ? w_vn_7 : _GEN_30179; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_30181 = 4'h8 == _T_3160 ? w_vn_8 : _GEN_30180; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_30182 = 4'h9 == _T_3160 ? 5'h0 : _GEN_30181; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_30183 = 4'ha == _T_3160 ? 5'h0 : _GEN_30182; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_30184 = 4'hb == _T_3160 ? w_vn_11 : _GEN_30183; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_30185 = 4'hc == _T_3160 ? w_vn_12 : _GEN_30184; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_30186 = 4'hd == _T_3160 ? w_vn_13 : _GEN_30185; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_30187 = 4'he == _T_3160 ? 5'h0 : _GEN_30186; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_30188 = 4'hf == _T_3160 ? w_vn_15 : _GEN_30187; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_95374 = {{1'd0}, _T_3160}; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_30189 = 5'h10 == _GEN_95374 ? w_vn_16 : _GEN_30188; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_30190 = 5'h11 == _GEN_95374 ? 5'h0 : _GEN_30189; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_30191 = 5'h12 == _GEN_95374 ? w_vn_18 : _GEN_30190; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_30192 = 5'h13 == _GEN_95374 ? 5'h0 : _GEN_30191; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_30193 = 5'h14 == _GEN_95374 ? 5'h0 : _GEN_30192; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_30194 = 5'h15 == _GEN_95374 ? 5'h0 : _GEN_30193; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_30195 = 5'h16 == _GEN_95374 ? 5'h0 : _GEN_30194; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_30196 = 5'h17 == _GEN_95374 ? w_vn_23 : _GEN_30195; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_30197 = 5'h18 == _GEN_95374 ? w_vn_24 : _GEN_30196; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_30198 = 5'h19 == _GEN_95374 ? 5'h0 : _GEN_30197; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_30199 = 5'h1a == _GEN_95374 ? 5'h0 : _GEN_30198; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_30200 = 5'h1b == _GEN_95374 ? 5'h0 : _GEN_30199; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_30201 = 5'h1c == _GEN_95374 ? 5'h0 : _GEN_30200; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_30202 = 5'h1d == _GEN_95374 ? 5'h0 : _GEN_30201; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_30203 = 5'h1e == _GEN_95374 ? 5'h0 : _GEN_30202; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_30204 = 5'h1f == _GEN_95374 ? 5'h0 : _GEN_30203; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_30208 = 4'h3 == _T_3163 ? w_vn_3 : 5'h0; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_30209 = 4'h4 == _T_3163 ? w_vn_4 : _GEN_30208; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_30210 = 4'h5 == _T_3163 ? 5'h0 : _GEN_30209; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_30211 = 4'h6 == _T_3163 ? 5'h0 : _GEN_30210; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_30212 = 4'h7 == _T_3163 ? w_vn_7 : _GEN_30211; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_30213 = 4'h8 == _T_3163 ? w_vn_8 : _GEN_30212; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_30214 = 4'h9 == _T_3163 ? 5'h0 : _GEN_30213; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_30215 = 4'ha == _T_3163 ? 5'h0 : _GEN_30214; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_30216 = 4'hb == _T_3163 ? w_vn_11 : _GEN_30215; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_30217 = 4'hc == _T_3163 ? w_vn_12 : _GEN_30216; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_30218 = 4'hd == _T_3163 ? w_vn_13 : _GEN_30217; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_30219 = 4'he == _T_3163 ? 5'h0 : _GEN_30218; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_30220 = 4'hf == _T_3163 ? w_vn_15 : _GEN_30219; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_95390 = {{1'd0}, _T_3163}; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_30221 = 5'h10 == _GEN_95390 ? w_vn_16 : _GEN_30220; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_30222 = 5'h11 == _GEN_95390 ? 5'h0 : _GEN_30221; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_30223 = 5'h12 == _GEN_95390 ? w_vn_18 : _GEN_30222; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_30224 = 5'h13 == _GEN_95390 ? 5'h0 : _GEN_30223; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_30225 = 5'h14 == _GEN_95390 ? 5'h0 : _GEN_30224; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_30226 = 5'h15 == _GEN_95390 ? 5'h0 : _GEN_30225; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_30227 = 5'h16 == _GEN_95390 ? 5'h0 : _GEN_30226; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_30228 = 5'h17 == _GEN_95390 ? w_vn_23 : _GEN_30227; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_30229 = 5'h18 == _GEN_95390 ? w_vn_24 : _GEN_30228; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_30230 = 5'h19 == _GEN_95390 ? 5'h0 : _GEN_30229; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_30231 = 5'h1a == _GEN_95390 ? 5'h0 : _GEN_30230; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_30232 = 5'h1b == _GEN_95390 ? 5'h0 : _GEN_30231; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_30233 = 5'h1c == _GEN_95390 ? 5'h0 : _GEN_30232; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_30234 = 5'h1d == _GEN_95390 ? 5'h0 : _GEN_30233; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_30235 = 5'h1e == _GEN_95390 ? 5'h0 : _GEN_30234; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_30236 = 5'h1f == _GEN_95390 ? 5'h0 : _GEN_30235; // @[FanCtrl.scala 160:{37,37}]
  wire  _T_3164 = _GEN_30204 == _GEN_30236; // @[FanCtrl.scala 160:37]
  wire [4:0] _T_3170 = {{1'd0}, _T_3158}; // @[FanCtrl.scala 166:30]
  wire [4:0] _GEN_30333 = 4'h3 == _T_3170[3:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_30334 = 4'h4 == _T_3170[3:0] ? w_vn_4 : _GEN_30333; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_30335 = 4'h5 == _T_3170[3:0] ? 5'h0 : _GEN_30334; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_30336 = 4'h6 == _T_3170[3:0] ? 5'h0 : _GEN_30335; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_30337 = 4'h7 == _T_3170[3:0] ? w_vn_7 : _GEN_30336; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_30338 = 4'h8 == _T_3170[3:0] ? w_vn_8 : _GEN_30337; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_30339 = 4'h9 == _T_3170[3:0] ? 5'h0 : _GEN_30338; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_30340 = 4'ha == _T_3170[3:0] ? 5'h0 : _GEN_30339; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_30341 = 4'hb == _T_3170[3:0] ? w_vn_11 : _GEN_30340; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_30342 = 4'hc == _T_3170[3:0] ? w_vn_12 : _GEN_30341; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_30343 = 4'hd == _T_3170[3:0] ? w_vn_13 : _GEN_30342; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_30344 = 4'he == _T_3170[3:0] ? 5'h0 : _GEN_30343; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_30345 = 4'hf == _T_3170[3:0] ? w_vn_15 : _GEN_30344; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_95406 = {{1'd0}, _T_3170[3:0]}; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_30346 = 5'h10 == _GEN_95406 ? w_vn_16 : _GEN_30345; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_30347 = 5'h11 == _GEN_95406 ? 5'h0 : _GEN_30346; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_30348 = 5'h12 == _GEN_95406 ? w_vn_18 : _GEN_30347; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_30349 = 5'h13 == _GEN_95406 ? 5'h0 : _GEN_30348; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_30350 = 5'h14 == _GEN_95406 ? 5'h0 : _GEN_30349; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_30351 = 5'h15 == _GEN_95406 ? 5'h0 : _GEN_30350; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_30352 = 5'h16 == _GEN_95406 ? 5'h0 : _GEN_30351; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_30353 = 5'h17 == _GEN_95406 ? w_vn_23 : _GEN_30352; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_30354 = 5'h18 == _GEN_95406 ? w_vn_24 : _GEN_30353; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_30355 = 5'h19 == _GEN_95406 ? 5'h0 : _GEN_30354; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_30356 = 5'h1a == _GEN_95406 ? 5'h0 : _GEN_30355; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_30357 = 5'h1b == _GEN_95406 ? 5'h0 : _GEN_30356; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_30358 = 5'h1c == _GEN_95406 ? 5'h0 : _GEN_30357; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_30359 = 5'h1d == _GEN_95406 ? 5'h0 : _GEN_30358; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_30360 = 5'h1e == _GEN_95406 ? 5'h0 : _GEN_30359; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_30361 = 5'h1f == _GEN_95406 ? 5'h0 : _GEN_30360; // @[FanCtrl.scala 166:{38,38}]
  wire  _T_3175 = _GEN_30361 == _GEN_30204; // @[FanCtrl.scala 166:38]
  wire [3:0] _T_3181 = _T_3158 + 4'h3; // @[FanCtrl.scala 167:55]
  wire [4:0] _GEN_30429 = 4'h3 == _T_3181 ? w_vn_3 : 5'h0; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_30430 = 4'h4 == _T_3181 ? w_vn_4 : _GEN_30429; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_30431 = 4'h5 == _T_3181 ? 5'h0 : _GEN_30430; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_30432 = 4'h6 == _T_3181 ? 5'h0 : _GEN_30431; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_30433 = 4'h7 == _T_3181 ? w_vn_7 : _GEN_30432; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_30434 = 4'h8 == _T_3181 ? w_vn_8 : _GEN_30433; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_30435 = 4'h9 == _T_3181 ? 5'h0 : _GEN_30434; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_30436 = 4'ha == _T_3181 ? 5'h0 : _GEN_30435; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_30437 = 4'hb == _T_3181 ? w_vn_11 : _GEN_30436; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_30438 = 4'hc == _T_3181 ? w_vn_12 : _GEN_30437; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_30439 = 4'hd == _T_3181 ? w_vn_13 : _GEN_30438; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_30440 = 4'he == _T_3181 ? 5'h0 : _GEN_30439; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_30441 = 4'hf == _T_3181 ? w_vn_15 : _GEN_30440; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_95454 = {{1'd0}, _T_3181}; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_30442 = 5'h10 == _GEN_95454 ? w_vn_16 : _GEN_30441; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_30443 = 5'h11 == _GEN_95454 ? 5'h0 : _GEN_30442; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_30444 = 5'h12 == _GEN_95454 ? w_vn_18 : _GEN_30443; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_30445 = 5'h13 == _GEN_95454 ? 5'h0 : _GEN_30444; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_30446 = 5'h14 == _GEN_95454 ? 5'h0 : _GEN_30445; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_30447 = 5'h15 == _GEN_95454 ? 5'h0 : _GEN_30446; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_30448 = 5'h16 == _GEN_95454 ? 5'h0 : _GEN_30447; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_30449 = 5'h17 == _GEN_95454 ? w_vn_23 : _GEN_30448; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_30450 = 5'h18 == _GEN_95454 ? w_vn_24 : _GEN_30449; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_30451 = 5'h19 == _GEN_95454 ? 5'h0 : _GEN_30450; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_30452 = 5'h1a == _GEN_95454 ? 5'h0 : _GEN_30451; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_30453 = 5'h1b == _GEN_95454 ? 5'h0 : _GEN_30452; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_30454 = 5'h1c == _GEN_95454 ? 5'h0 : _GEN_30453; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_30455 = 5'h1d == _GEN_95454 ? 5'h0 : _GEN_30454; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_30456 = 5'h1e == _GEN_95454 ? 5'h0 : _GEN_30455; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_30457 = 5'h1f == _GEN_95454 ? 5'h0 : _GEN_30456; // @[FanCtrl.scala 167:{36,36}]
  wire  _T_3182 = _GEN_30236 == _GEN_30457; // @[FanCtrl.scala 167:36]
  wire  _T_3183 = _GEN_30361 == _GEN_30204 & _T_3182; // @[FanCtrl.scala 166:65]
  wire [3:0] _T_3186 = _T_3158 + 4'h4; // @[FanCtrl.scala 168:29]
  wire [4:0] _GEN_30461 = 4'h3 == _T_3186 ? w_vn_3 : 5'h0; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_30462 = 4'h4 == _T_3186 ? w_vn_4 : _GEN_30461; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_30463 = 4'h5 == _T_3186 ? 5'h0 : _GEN_30462; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_30464 = 4'h6 == _T_3186 ? 5'h0 : _GEN_30463; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_30465 = 4'h7 == _T_3186 ? w_vn_7 : _GEN_30464; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_30466 = 4'h8 == _T_3186 ? w_vn_8 : _GEN_30465; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_30467 = 4'h9 == _T_3186 ? 5'h0 : _GEN_30466; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_30468 = 4'ha == _T_3186 ? 5'h0 : _GEN_30467; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_30469 = 4'hb == _T_3186 ? w_vn_11 : _GEN_30468; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_30470 = 4'hc == _T_3186 ? w_vn_12 : _GEN_30469; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_30471 = 4'hd == _T_3186 ? w_vn_13 : _GEN_30470; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_30472 = 4'he == _T_3186 ? 5'h0 : _GEN_30471; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_30473 = 4'hf == _T_3186 ? w_vn_15 : _GEN_30472; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_95470 = {{1'd0}, _T_3186}; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_30474 = 5'h10 == _GEN_95470 ? w_vn_16 : _GEN_30473; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_30475 = 5'h11 == _GEN_95470 ? 5'h0 : _GEN_30474; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_30476 = 5'h12 == _GEN_95470 ? w_vn_18 : _GEN_30475; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_30477 = 5'h13 == _GEN_95470 ? 5'h0 : _GEN_30476; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_30478 = 5'h14 == _GEN_95470 ? 5'h0 : _GEN_30477; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_30479 = 5'h15 == _GEN_95470 ? 5'h0 : _GEN_30478; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_30480 = 5'h16 == _GEN_95470 ? 5'h0 : _GEN_30479; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_30481 = 5'h17 == _GEN_95470 ? w_vn_23 : _GEN_30480; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_30482 = 5'h18 == _GEN_95470 ? w_vn_24 : _GEN_30481; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_30483 = 5'h19 == _GEN_95470 ? 5'h0 : _GEN_30482; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_30484 = 5'h1a == _GEN_95470 ? 5'h0 : _GEN_30483; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_30485 = 5'h1b == _GEN_95470 ? 5'h0 : _GEN_30484; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_30486 = 5'h1c == _GEN_95470 ? 5'h0 : _GEN_30485; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_30487 = 5'h1d == _GEN_95470 ? 5'h0 : _GEN_30486; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_30488 = 5'h1e == _GEN_95470 ? 5'h0 : _GEN_30487; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_30489 = 5'h1f == _GEN_95470 ? 5'h0 : _GEN_30488; // @[FanCtrl.scala 168:{37,37}]
  wire  _T_3190 = _GEN_30489 != _GEN_30457; // @[FanCtrl.scala 168:37]
  wire  _T_3191 = _T_3183 & _T_3190; // @[FanCtrl.scala 167:64]
  wire  _T_3198 = _GEN_30204 != _GEN_30236; // @[FanCtrl.scala 169:37]
  wire  _T_3199 = _T_3191 & _T_3198; // @[FanCtrl.scala 168:64]
  wire  _T_3216 = _T_3182 & _T_3190; // @[FanCtrl.scala 173:71]
  wire  _T_3224 = _T_3216 & _T_3198; // @[FanCtrl.scala 174:71]
  wire  _T_3241 = _T_3175 & _T_3198; // @[FanCtrl.scala 179:71]
  wire [2:0] _GEN_31046 = _T_3241 ? 3'h3 : 3'h0; // @[FanCtrl.scala 180:72]
  wire [2:0] _GEN_31077 = _T_3224 ? 3'h4 : _GEN_31046; // @[FanCtrl.scala 175:72]
  wire [2:0] _GEN_31108 = _T_3199 ? 3'h5 : _GEN_31077; // @[FanCtrl.scala 169:66]
  wire  _GEN_31201 = r_valid_1 & _T_3164; // @[FanCtrl.scala 159:32]
  wire [2:0] _GEN_31232 = r_valid_1 ? _GEN_31108 : 3'h0; // @[FanCtrl.scala 159:32]
  wire [3:0] _T_3467 = 3'h4 * 1'h1; // @[FanCtrl.scala 160:23]
  wire [3:0] _T_3469 = _T_3467 + 4'h1; // @[FanCtrl.scala 160:29]
  wire [3:0] _T_3472 = _T_3467 + 4'h2; // @[FanCtrl.scala 160:56]
  wire [4:0] _GEN_33836 = 4'h3 == _T_3469 ? w_vn_3 : 5'h0; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_33837 = 4'h4 == _T_3469 ? w_vn_4 : _GEN_33836; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_33838 = 4'h5 == _T_3469 ? 5'h0 : _GEN_33837; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_33839 = 4'h6 == _T_3469 ? 5'h0 : _GEN_33838; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_33840 = 4'h7 == _T_3469 ? w_vn_7 : _GEN_33839; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_33841 = 4'h8 == _T_3469 ? w_vn_8 : _GEN_33840; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_33842 = 4'h9 == _T_3469 ? 5'h0 : _GEN_33841; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_33843 = 4'ha == _T_3469 ? 5'h0 : _GEN_33842; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_33844 = 4'hb == _T_3469 ? w_vn_11 : _GEN_33843; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_33845 = 4'hc == _T_3469 ? w_vn_12 : _GEN_33844; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_33846 = 4'hd == _T_3469 ? w_vn_13 : _GEN_33845; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_33847 = 4'he == _T_3469 ? 5'h0 : _GEN_33846; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_33848 = 4'hf == _T_3469 ? w_vn_15 : _GEN_33847; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_96398 = {{1'd0}, _T_3469}; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_33849 = 5'h10 == _GEN_96398 ? w_vn_16 : _GEN_33848; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_33850 = 5'h11 == _GEN_96398 ? 5'h0 : _GEN_33849; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_33851 = 5'h12 == _GEN_96398 ? w_vn_18 : _GEN_33850; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_33852 = 5'h13 == _GEN_96398 ? 5'h0 : _GEN_33851; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_33853 = 5'h14 == _GEN_96398 ? 5'h0 : _GEN_33852; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_33854 = 5'h15 == _GEN_96398 ? 5'h0 : _GEN_33853; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_33855 = 5'h16 == _GEN_96398 ? 5'h0 : _GEN_33854; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_33856 = 5'h17 == _GEN_96398 ? w_vn_23 : _GEN_33855; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_33857 = 5'h18 == _GEN_96398 ? w_vn_24 : _GEN_33856; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_33858 = 5'h19 == _GEN_96398 ? 5'h0 : _GEN_33857; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_33859 = 5'h1a == _GEN_96398 ? 5'h0 : _GEN_33858; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_33860 = 5'h1b == _GEN_96398 ? 5'h0 : _GEN_33859; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_33861 = 5'h1c == _GEN_96398 ? 5'h0 : _GEN_33860; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_33862 = 5'h1d == _GEN_96398 ? 5'h0 : _GEN_33861; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_33863 = 5'h1e == _GEN_96398 ? 5'h0 : _GEN_33862; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_33864 = 5'h1f == _GEN_96398 ? 5'h0 : _GEN_33863; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_33868 = 4'h3 == _T_3472 ? w_vn_3 : 5'h0; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_33869 = 4'h4 == _T_3472 ? w_vn_4 : _GEN_33868; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_33870 = 4'h5 == _T_3472 ? 5'h0 : _GEN_33869; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_33871 = 4'h6 == _T_3472 ? 5'h0 : _GEN_33870; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_33872 = 4'h7 == _T_3472 ? w_vn_7 : _GEN_33871; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_33873 = 4'h8 == _T_3472 ? w_vn_8 : _GEN_33872; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_33874 = 4'h9 == _T_3472 ? 5'h0 : _GEN_33873; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_33875 = 4'ha == _T_3472 ? 5'h0 : _GEN_33874; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_33876 = 4'hb == _T_3472 ? w_vn_11 : _GEN_33875; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_33877 = 4'hc == _T_3472 ? w_vn_12 : _GEN_33876; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_33878 = 4'hd == _T_3472 ? w_vn_13 : _GEN_33877; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_33879 = 4'he == _T_3472 ? 5'h0 : _GEN_33878; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_33880 = 4'hf == _T_3472 ? w_vn_15 : _GEN_33879; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_96414 = {{1'd0}, _T_3472}; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_33881 = 5'h10 == _GEN_96414 ? w_vn_16 : _GEN_33880; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_33882 = 5'h11 == _GEN_96414 ? 5'h0 : _GEN_33881; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_33883 = 5'h12 == _GEN_96414 ? w_vn_18 : _GEN_33882; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_33884 = 5'h13 == _GEN_96414 ? 5'h0 : _GEN_33883; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_33885 = 5'h14 == _GEN_96414 ? 5'h0 : _GEN_33884; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_33886 = 5'h15 == _GEN_96414 ? 5'h0 : _GEN_33885; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_33887 = 5'h16 == _GEN_96414 ? 5'h0 : _GEN_33886; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_33888 = 5'h17 == _GEN_96414 ? w_vn_23 : _GEN_33887; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_33889 = 5'h18 == _GEN_96414 ? w_vn_24 : _GEN_33888; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_33890 = 5'h19 == _GEN_96414 ? 5'h0 : _GEN_33889; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_33891 = 5'h1a == _GEN_96414 ? 5'h0 : _GEN_33890; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_33892 = 5'h1b == _GEN_96414 ? 5'h0 : _GEN_33891; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_33893 = 5'h1c == _GEN_96414 ? 5'h0 : _GEN_33892; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_33894 = 5'h1d == _GEN_96414 ? 5'h0 : _GEN_33893; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_33895 = 5'h1e == _GEN_96414 ? 5'h0 : _GEN_33894; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_33896 = 5'h1f == _GEN_96414 ? 5'h0 : _GEN_33895; // @[FanCtrl.scala 160:{37,37}]
  wire  _T_3473 = _GEN_33864 == _GEN_33896; // @[FanCtrl.scala 160:37]
  wire [4:0] _T_3479 = {{1'd0}, _T_3467}; // @[FanCtrl.scala 166:30]
  wire [4:0] _GEN_33993 = 4'h3 == _T_3479[3:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_33994 = 4'h4 == _T_3479[3:0] ? w_vn_4 : _GEN_33993; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_33995 = 4'h5 == _T_3479[3:0] ? 5'h0 : _GEN_33994; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_33996 = 4'h6 == _T_3479[3:0] ? 5'h0 : _GEN_33995; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_33997 = 4'h7 == _T_3479[3:0] ? w_vn_7 : _GEN_33996; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_33998 = 4'h8 == _T_3479[3:0] ? w_vn_8 : _GEN_33997; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_33999 = 4'h9 == _T_3479[3:0] ? 5'h0 : _GEN_33998; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_34000 = 4'ha == _T_3479[3:0] ? 5'h0 : _GEN_33999; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_34001 = 4'hb == _T_3479[3:0] ? w_vn_11 : _GEN_34000; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_34002 = 4'hc == _T_3479[3:0] ? w_vn_12 : _GEN_34001; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_34003 = 4'hd == _T_3479[3:0] ? w_vn_13 : _GEN_34002; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_34004 = 4'he == _T_3479[3:0] ? 5'h0 : _GEN_34003; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_34005 = 4'hf == _T_3479[3:0] ? w_vn_15 : _GEN_34004; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_96430 = {{1'd0}, _T_3479[3:0]}; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_34006 = 5'h10 == _GEN_96430 ? w_vn_16 : _GEN_34005; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_34007 = 5'h11 == _GEN_96430 ? 5'h0 : _GEN_34006; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_34008 = 5'h12 == _GEN_96430 ? w_vn_18 : _GEN_34007; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_34009 = 5'h13 == _GEN_96430 ? 5'h0 : _GEN_34008; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_34010 = 5'h14 == _GEN_96430 ? 5'h0 : _GEN_34009; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_34011 = 5'h15 == _GEN_96430 ? 5'h0 : _GEN_34010; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_34012 = 5'h16 == _GEN_96430 ? 5'h0 : _GEN_34011; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_34013 = 5'h17 == _GEN_96430 ? w_vn_23 : _GEN_34012; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_34014 = 5'h18 == _GEN_96430 ? w_vn_24 : _GEN_34013; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_34015 = 5'h19 == _GEN_96430 ? 5'h0 : _GEN_34014; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_34016 = 5'h1a == _GEN_96430 ? 5'h0 : _GEN_34015; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_34017 = 5'h1b == _GEN_96430 ? 5'h0 : _GEN_34016; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_34018 = 5'h1c == _GEN_96430 ? 5'h0 : _GEN_34017; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_34019 = 5'h1d == _GEN_96430 ? 5'h0 : _GEN_34018; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_34020 = 5'h1e == _GEN_96430 ? 5'h0 : _GEN_34019; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_34021 = 5'h1f == _GEN_96430 ? 5'h0 : _GEN_34020; // @[FanCtrl.scala 166:{38,38}]
  wire  _T_3484 = _GEN_34021 == _GEN_33864; // @[FanCtrl.scala 166:38]
  wire [3:0] _T_3490 = _T_3467 + 4'h3; // @[FanCtrl.scala 167:55]
  wire [4:0] _GEN_34089 = 4'h3 == _T_3490 ? w_vn_3 : 5'h0; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_34090 = 4'h4 == _T_3490 ? w_vn_4 : _GEN_34089; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_34091 = 4'h5 == _T_3490 ? 5'h0 : _GEN_34090; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_34092 = 4'h6 == _T_3490 ? 5'h0 : _GEN_34091; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_34093 = 4'h7 == _T_3490 ? w_vn_7 : _GEN_34092; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_34094 = 4'h8 == _T_3490 ? w_vn_8 : _GEN_34093; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_34095 = 4'h9 == _T_3490 ? 5'h0 : _GEN_34094; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_34096 = 4'ha == _T_3490 ? 5'h0 : _GEN_34095; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_34097 = 4'hb == _T_3490 ? w_vn_11 : _GEN_34096; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_34098 = 4'hc == _T_3490 ? w_vn_12 : _GEN_34097; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_34099 = 4'hd == _T_3490 ? w_vn_13 : _GEN_34098; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_34100 = 4'he == _T_3490 ? 5'h0 : _GEN_34099; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_34101 = 4'hf == _T_3490 ? w_vn_15 : _GEN_34100; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_96478 = {{1'd0}, _T_3490}; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_34102 = 5'h10 == _GEN_96478 ? w_vn_16 : _GEN_34101; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_34103 = 5'h11 == _GEN_96478 ? 5'h0 : _GEN_34102; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_34104 = 5'h12 == _GEN_96478 ? w_vn_18 : _GEN_34103; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_34105 = 5'h13 == _GEN_96478 ? 5'h0 : _GEN_34104; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_34106 = 5'h14 == _GEN_96478 ? 5'h0 : _GEN_34105; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_34107 = 5'h15 == _GEN_96478 ? 5'h0 : _GEN_34106; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_34108 = 5'h16 == _GEN_96478 ? 5'h0 : _GEN_34107; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_34109 = 5'h17 == _GEN_96478 ? w_vn_23 : _GEN_34108; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_34110 = 5'h18 == _GEN_96478 ? w_vn_24 : _GEN_34109; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_34111 = 5'h19 == _GEN_96478 ? 5'h0 : _GEN_34110; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_34112 = 5'h1a == _GEN_96478 ? 5'h0 : _GEN_34111; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_34113 = 5'h1b == _GEN_96478 ? 5'h0 : _GEN_34112; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_34114 = 5'h1c == _GEN_96478 ? 5'h0 : _GEN_34113; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_34115 = 5'h1d == _GEN_96478 ? 5'h0 : _GEN_34114; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_34116 = 5'h1e == _GEN_96478 ? 5'h0 : _GEN_34115; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_34117 = 5'h1f == _GEN_96478 ? 5'h0 : _GEN_34116; // @[FanCtrl.scala 167:{36,36}]
  wire  _T_3491 = _GEN_33896 == _GEN_34117; // @[FanCtrl.scala 167:36]
  wire  _T_3492 = _GEN_34021 == _GEN_33864 & _T_3491; // @[FanCtrl.scala 166:65]
  wire [3:0] _T_3495 = _T_3467 + 4'h4; // @[FanCtrl.scala 168:29]
  wire [4:0] _GEN_34121 = 4'h3 == _T_3495 ? w_vn_3 : 5'h0; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_34122 = 4'h4 == _T_3495 ? w_vn_4 : _GEN_34121; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_34123 = 4'h5 == _T_3495 ? 5'h0 : _GEN_34122; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_34124 = 4'h6 == _T_3495 ? 5'h0 : _GEN_34123; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_34125 = 4'h7 == _T_3495 ? w_vn_7 : _GEN_34124; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_34126 = 4'h8 == _T_3495 ? w_vn_8 : _GEN_34125; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_34127 = 4'h9 == _T_3495 ? 5'h0 : _GEN_34126; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_34128 = 4'ha == _T_3495 ? 5'h0 : _GEN_34127; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_34129 = 4'hb == _T_3495 ? w_vn_11 : _GEN_34128; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_34130 = 4'hc == _T_3495 ? w_vn_12 : _GEN_34129; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_34131 = 4'hd == _T_3495 ? w_vn_13 : _GEN_34130; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_34132 = 4'he == _T_3495 ? 5'h0 : _GEN_34131; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_34133 = 4'hf == _T_3495 ? w_vn_15 : _GEN_34132; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_96494 = {{1'd0}, _T_3495}; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_34134 = 5'h10 == _GEN_96494 ? w_vn_16 : _GEN_34133; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_34135 = 5'h11 == _GEN_96494 ? 5'h0 : _GEN_34134; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_34136 = 5'h12 == _GEN_96494 ? w_vn_18 : _GEN_34135; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_34137 = 5'h13 == _GEN_96494 ? 5'h0 : _GEN_34136; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_34138 = 5'h14 == _GEN_96494 ? 5'h0 : _GEN_34137; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_34139 = 5'h15 == _GEN_96494 ? 5'h0 : _GEN_34138; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_34140 = 5'h16 == _GEN_96494 ? 5'h0 : _GEN_34139; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_34141 = 5'h17 == _GEN_96494 ? w_vn_23 : _GEN_34140; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_34142 = 5'h18 == _GEN_96494 ? w_vn_24 : _GEN_34141; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_34143 = 5'h19 == _GEN_96494 ? 5'h0 : _GEN_34142; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_34144 = 5'h1a == _GEN_96494 ? 5'h0 : _GEN_34143; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_34145 = 5'h1b == _GEN_96494 ? 5'h0 : _GEN_34144; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_34146 = 5'h1c == _GEN_96494 ? 5'h0 : _GEN_34145; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_34147 = 5'h1d == _GEN_96494 ? 5'h0 : _GEN_34146; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_34148 = 5'h1e == _GEN_96494 ? 5'h0 : _GEN_34147; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_34149 = 5'h1f == _GEN_96494 ? 5'h0 : _GEN_34148; // @[FanCtrl.scala 168:{37,37}]
  wire  _T_3499 = _GEN_34149 != _GEN_34117; // @[FanCtrl.scala 168:37]
  wire  _T_3507 = _GEN_33864 != _GEN_33896; // @[FanCtrl.scala 169:37]
  wire  _T_3525 = _T_3491 & _T_3499; // @[FanCtrl.scala 173:71]
  wire  _T_3533 = _T_3525 & _T_3507; // @[FanCtrl.scala 174:71]
  wire  _GEN_34862 = r_valid_1 & _T_3473; // @[FanCtrl.scala 159:32]
  wire [3:0] _T_3596 = _T_3467 - 4'h1; // @[FanCtrl.scala 203:56]
  wire [4:0] _GEN_35289 = 4'h3 == _T_3596 ? w_vn_3 : 5'h0; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_35290 = 4'h4 == _T_3596 ? w_vn_4 : _GEN_35289; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_35291 = 4'h5 == _T_3596 ? 5'h0 : _GEN_35290; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_35292 = 4'h6 == _T_3596 ? 5'h0 : _GEN_35291; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_35293 = 4'h7 == _T_3596 ? w_vn_7 : _GEN_35292; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_35294 = 4'h8 == _T_3596 ? w_vn_8 : _GEN_35293; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_35295 = 4'h9 == _T_3596 ? 5'h0 : _GEN_35294; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_35296 = 4'ha == _T_3596 ? 5'h0 : _GEN_35295; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_35297 = 4'hb == _T_3596 ? w_vn_11 : _GEN_35296; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_35298 = 4'hc == _T_3596 ? w_vn_12 : _GEN_35297; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_35299 = 4'hd == _T_3596 ? w_vn_13 : _GEN_35298; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_35300 = 4'he == _T_3596 ? 5'h0 : _GEN_35299; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_35301 = 4'hf == _T_3596 ? w_vn_15 : _GEN_35300; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_96830 = {{1'd0}, _T_3596}; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_35302 = 5'h10 == _GEN_96830 ? w_vn_16 : _GEN_35301; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_35303 = 5'h11 == _GEN_96830 ? 5'h0 : _GEN_35302; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_35304 = 5'h12 == _GEN_96830 ? w_vn_18 : _GEN_35303; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_35305 = 5'h13 == _GEN_96830 ? 5'h0 : _GEN_35304; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_35306 = 5'h14 == _GEN_96830 ? 5'h0 : _GEN_35305; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_35307 = 5'h15 == _GEN_96830 ? 5'h0 : _GEN_35306; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_35308 = 5'h16 == _GEN_96830 ? 5'h0 : _GEN_35307; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_35309 = 5'h17 == _GEN_96830 ? w_vn_23 : _GEN_35308; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_35310 = 5'h18 == _GEN_96830 ? w_vn_24 : _GEN_35309; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_35311 = 5'h19 == _GEN_96830 ? 5'h0 : _GEN_35310; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_35312 = 5'h1a == _GEN_96830 ? 5'h0 : _GEN_35311; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_35313 = 5'h1b == _GEN_96830 ? 5'h0 : _GEN_35312; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_35314 = 5'h1c == _GEN_96830 ? 5'h0 : _GEN_35313; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_35315 = 5'h1d == _GEN_96830 ? 5'h0 : _GEN_35314; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_35316 = 5'h1e == _GEN_96830 ? 5'h0 : _GEN_35315; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_35317 = 5'h1f == _GEN_96830 ? 5'h0 : _GEN_35316; // @[FanCtrl.scala 203:{37,37}]
  wire  _T_3597 = _GEN_34021 != _GEN_35317; // @[FanCtrl.scala 203:37]
  wire  _T_3598 = _T_3492 & _T_3597; // @[FanCtrl.scala 202:65]
  wire  _T_3623 = _T_3484 & _T_3597; // @[FanCtrl.scala 208:71]
  wire  _T_3631 = _T_3623 & _T_3507; // @[FanCtrl.scala 209:70]
  wire  _T_3703 = _T_3598 & _T_3499; // @[FanCtrl.scala 239:64]
  wire  _T_3711 = _T_3703 & _T_3507; // @[FanCtrl.scala 240:62]
  wire [2:0] _GEN_37107 = _T_3631 ? 3'h3 : 3'h0; // @[FanCtrl.scala 253:70]
  wire [2:0] _GEN_37138 = _T_3533 ? 3'h4 : _GEN_37107; // @[FanCtrl.scala 247:70]
  wire [2:0] _GEN_37169 = _T_3711 ? 3'h5 : _GEN_37138; // @[FanCtrl.scala 241:64]
  wire [2:0] _GEN_37293 = r_valid_1 ? _GEN_37169 : 3'h0; // @[FanCtrl.scala 230:30]
  wire [4:0] _T_3776 = 3'h4 * 2'h2; // @[FanCtrl.scala 160:23]
  wire [4:0] _T_3778 = _T_3776 + 5'h1; // @[FanCtrl.scala 160:29]
  wire [4:0] _T_3781 = _T_3776 + 5'h2; // @[FanCtrl.scala 160:56]
  wire [4:0] _GEN_37496 = 5'h3 == _T_3778 ? w_vn_3 : 5'h0; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_37497 = 5'h4 == _T_3778 ? w_vn_4 : _GEN_37496; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_37498 = 5'h5 == _T_3778 ? 5'h0 : _GEN_37497; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_37499 = 5'h6 == _T_3778 ? 5'h0 : _GEN_37498; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_37500 = 5'h7 == _T_3778 ? w_vn_7 : _GEN_37499; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_37501 = 5'h8 == _T_3778 ? w_vn_8 : _GEN_37500; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_37502 = 5'h9 == _T_3778 ? 5'h0 : _GEN_37501; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_37503 = 5'ha == _T_3778 ? 5'h0 : _GEN_37502; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_37504 = 5'hb == _T_3778 ? w_vn_11 : _GEN_37503; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_37505 = 5'hc == _T_3778 ? w_vn_12 : _GEN_37504; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_37506 = 5'hd == _T_3778 ? w_vn_13 : _GEN_37505; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_37507 = 5'he == _T_3778 ? 5'h0 : _GEN_37506; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_37508 = 5'hf == _T_3778 ? w_vn_15 : _GEN_37507; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_37509 = 5'h10 == _T_3778 ? w_vn_16 : _GEN_37508; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_37510 = 5'h11 == _T_3778 ? 5'h0 : _GEN_37509; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_37511 = 5'h12 == _T_3778 ? w_vn_18 : _GEN_37510; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_37512 = 5'h13 == _T_3778 ? 5'h0 : _GEN_37511; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_37513 = 5'h14 == _T_3778 ? 5'h0 : _GEN_37512; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_37514 = 5'h15 == _T_3778 ? 5'h0 : _GEN_37513; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_37515 = 5'h16 == _T_3778 ? 5'h0 : _GEN_37514; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_37516 = 5'h17 == _T_3778 ? w_vn_23 : _GEN_37515; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_37517 = 5'h18 == _T_3778 ? w_vn_24 : _GEN_37516; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_37518 = 5'h19 == _T_3778 ? 5'h0 : _GEN_37517; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_37519 = 5'h1a == _T_3778 ? 5'h0 : _GEN_37518; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_37520 = 5'h1b == _T_3778 ? 5'h0 : _GEN_37519; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_37521 = 5'h1c == _T_3778 ? 5'h0 : _GEN_37520; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_37522 = 5'h1d == _T_3778 ? 5'h0 : _GEN_37521; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_37523 = 5'h1e == _T_3778 ? 5'h0 : _GEN_37522; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_37524 = 5'h1f == _T_3778 ? 5'h0 : _GEN_37523; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_37528 = 5'h3 == _T_3781 ? w_vn_3 : 5'h0; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_37529 = 5'h4 == _T_3781 ? w_vn_4 : _GEN_37528; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_37530 = 5'h5 == _T_3781 ? 5'h0 : _GEN_37529; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_37531 = 5'h6 == _T_3781 ? 5'h0 : _GEN_37530; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_37532 = 5'h7 == _T_3781 ? w_vn_7 : _GEN_37531; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_37533 = 5'h8 == _T_3781 ? w_vn_8 : _GEN_37532; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_37534 = 5'h9 == _T_3781 ? 5'h0 : _GEN_37533; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_37535 = 5'ha == _T_3781 ? 5'h0 : _GEN_37534; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_37536 = 5'hb == _T_3781 ? w_vn_11 : _GEN_37535; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_37537 = 5'hc == _T_3781 ? w_vn_12 : _GEN_37536; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_37538 = 5'hd == _T_3781 ? w_vn_13 : _GEN_37537; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_37539 = 5'he == _T_3781 ? 5'h0 : _GEN_37538; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_37540 = 5'hf == _T_3781 ? w_vn_15 : _GEN_37539; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_37541 = 5'h10 == _T_3781 ? w_vn_16 : _GEN_37540; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_37542 = 5'h11 == _T_3781 ? 5'h0 : _GEN_37541; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_37543 = 5'h12 == _T_3781 ? w_vn_18 : _GEN_37542; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_37544 = 5'h13 == _T_3781 ? 5'h0 : _GEN_37543; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_37545 = 5'h14 == _T_3781 ? 5'h0 : _GEN_37544; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_37546 = 5'h15 == _T_3781 ? 5'h0 : _GEN_37545; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_37547 = 5'h16 == _T_3781 ? 5'h0 : _GEN_37546; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_37548 = 5'h17 == _T_3781 ? w_vn_23 : _GEN_37547; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_37549 = 5'h18 == _T_3781 ? w_vn_24 : _GEN_37548; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_37550 = 5'h19 == _T_3781 ? 5'h0 : _GEN_37549; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_37551 = 5'h1a == _T_3781 ? 5'h0 : _GEN_37550; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_37552 = 5'h1b == _T_3781 ? 5'h0 : _GEN_37551; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_37553 = 5'h1c == _T_3781 ? 5'h0 : _GEN_37552; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_37554 = 5'h1d == _T_3781 ? 5'h0 : _GEN_37553; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_37555 = 5'h1e == _T_3781 ? 5'h0 : _GEN_37554; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_37556 = 5'h1f == _T_3781 ? 5'h0 : _GEN_37555; // @[FanCtrl.scala 160:{37,37}]
  wire  _T_3782 = _GEN_37524 == _GEN_37556; // @[FanCtrl.scala 160:37]
  wire [5:0] _T_3788 = {{1'd0}, _T_3776}; // @[FanCtrl.scala 166:30]
  wire [4:0] _GEN_37653 = 5'h3 == _T_3788[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_37654 = 5'h4 == _T_3788[4:0] ? w_vn_4 : _GEN_37653; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_37655 = 5'h5 == _T_3788[4:0] ? 5'h0 : _GEN_37654; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_37656 = 5'h6 == _T_3788[4:0] ? 5'h0 : _GEN_37655; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_37657 = 5'h7 == _T_3788[4:0] ? w_vn_7 : _GEN_37656; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_37658 = 5'h8 == _T_3788[4:0] ? w_vn_8 : _GEN_37657; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_37659 = 5'h9 == _T_3788[4:0] ? 5'h0 : _GEN_37658; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_37660 = 5'ha == _T_3788[4:0] ? 5'h0 : _GEN_37659; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_37661 = 5'hb == _T_3788[4:0] ? w_vn_11 : _GEN_37660; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_37662 = 5'hc == _T_3788[4:0] ? w_vn_12 : _GEN_37661; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_37663 = 5'hd == _T_3788[4:0] ? w_vn_13 : _GEN_37662; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_37664 = 5'he == _T_3788[4:0] ? 5'h0 : _GEN_37663; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_37665 = 5'hf == _T_3788[4:0] ? w_vn_15 : _GEN_37664; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_37666 = 5'h10 == _T_3788[4:0] ? w_vn_16 : _GEN_37665; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_37667 = 5'h11 == _T_3788[4:0] ? 5'h0 : _GEN_37666; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_37668 = 5'h12 == _T_3788[4:0] ? w_vn_18 : _GEN_37667; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_37669 = 5'h13 == _T_3788[4:0] ? 5'h0 : _GEN_37668; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_37670 = 5'h14 == _T_3788[4:0] ? 5'h0 : _GEN_37669; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_37671 = 5'h15 == _T_3788[4:0] ? 5'h0 : _GEN_37670; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_37672 = 5'h16 == _T_3788[4:0] ? 5'h0 : _GEN_37671; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_37673 = 5'h17 == _T_3788[4:0] ? w_vn_23 : _GEN_37672; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_37674 = 5'h18 == _T_3788[4:0] ? w_vn_24 : _GEN_37673; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_37675 = 5'h19 == _T_3788[4:0] ? 5'h0 : _GEN_37674; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_37676 = 5'h1a == _T_3788[4:0] ? 5'h0 : _GEN_37675; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_37677 = 5'h1b == _T_3788[4:0] ? 5'h0 : _GEN_37676; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_37678 = 5'h1c == _T_3788[4:0] ? 5'h0 : _GEN_37677; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_37679 = 5'h1d == _T_3788[4:0] ? 5'h0 : _GEN_37678; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_37680 = 5'h1e == _T_3788[4:0] ? 5'h0 : _GEN_37679; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_37681 = 5'h1f == _T_3788[4:0] ? 5'h0 : _GEN_37680; // @[FanCtrl.scala 166:{38,38}]
  wire  _T_3793 = _GEN_37681 == _GEN_37524; // @[FanCtrl.scala 166:38]
  wire [4:0] _T_3799 = _T_3776 + 5'h3; // @[FanCtrl.scala 167:55]
  wire [4:0] _GEN_37749 = 5'h3 == _T_3799 ? w_vn_3 : 5'h0; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_37750 = 5'h4 == _T_3799 ? w_vn_4 : _GEN_37749; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_37751 = 5'h5 == _T_3799 ? 5'h0 : _GEN_37750; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_37752 = 5'h6 == _T_3799 ? 5'h0 : _GEN_37751; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_37753 = 5'h7 == _T_3799 ? w_vn_7 : _GEN_37752; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_37754 = 5'h8 == _T_3799 ? w_vn_8 : _GEN_37753; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_37755 = 5'h9 == _T_3799 ? 5'h0 : _GEN_37754; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_37756 = 5'ha == _T_3799 ? 5'h0 : _GEN_37755; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_37757 = 5'hb == _T_3799 ? w_vn_11 : _GEN_37756; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_37758 = 5'hc == _T_3799 ? w_vn_12 : _GEN_37757; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_37759 = 5'hd == _T_3799 ? w_vn_13 : _GEN_37758; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_37760 = 5'he == _T_3799 ? 5'h0 : _GEN_37759; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_37761 = 5'hf == _T_3799 ? w_vn_15 : _GEN_37760; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_37762 = 5'h10 == _T_3799 ? w_vn_16 : _GEN_37761; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_37763 = 5'h11 == _T_3799 ? 5'h0 : _GEN_37762; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_37764 = 5'h12 == _T_3799 ? w_vn_18 : _GEN_37763; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_37765 = 5'h13 == _T_3799 ? 5'h0 : _GEN_37764; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_37766 = 5'h14 == _T_3799 ? 5'h0 : _GEN_37765; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_37767 = 5'h15 == _T_3799 ? 5'h0 : _GEN_37766; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_37768 = 5'h16 == _T_3799 ? 5'h0 : _GEN_37767; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_37769 = 5'h17 == _T_3799 ? w_vn_23 : _GEN_37768; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_37770 = 5'h18 == _T_3799 ? w_vn_24 : _GEN_37769; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_37771 = 5'h19 == _T_3799 ? 5'h0 : _GEN_37770; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_37772 = 5'h1a == _T_3799 ? 5'h0 : _GEN_37771; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_37773 = 5'h1b == _T_3799 ? 5'h0 : _GEN_37772; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_37774 = 5'h1c == _T_3799 ? 5'h0 : _GEN_37773; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_37775 = 5'h1d == _T_3799 ? 5'h0 : _GEN_37774; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_37776 = 5'h1e == _T_3799 ? 5'h0 : _GEN_37775; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_37777 = 5'h1f == _T_3799 ? 5'h0 : _GEN_37776; // @[FanCtrl.scala 167:{36,36}]
  wire  _T_3800 = _GEN_37556 == _GEN_37777; // @[FanCtrl.scala 167:36]
  wire  _T_3801 = _GEN_37681 == _GEN_37524 & _T_3800; // @[FanCtrl.scala 166:65]
  wire [4:0] _T_3804 = _T_3776 + 5'h4; // @[FanCtrl.scala 168:29]
  wire [4:0] _GEN_37781 = 5'h3 == _T_3804 ? w_vn_3 : 5'h0; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_37782 = 5'h4 == _T_3804 ? w_vn_4 : _GEN_37781; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_37783 = 5'h5 == _T_3804 ? 5'h0 : _GEN_37782; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_37784 = 5'h6 == _T_3804 ? 5'h0 : _GEN_37783; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_37785 = 5'h7 == _T_3804 ? w_vn_7 : _GEN_37784; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_37786 = 5'h8 == _T_3804 ? w_vn_8 : _GEN_37785; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_37787 = 5'h9 == _T_3804 ? 5'h0 : _GEN_37786; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_37788 = 5'ha == _T_3804 ? 5'h0 : _GEN_37787; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_37789 = 5'hb == _T_3804 ? w_vn_11 : _GEN_37788; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_37790 = 5'hc == _T_3804 ? w_vn_12 : _GEN_37789; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_37791 = 5'hd == _T_3804 ? w_vn_13 : _GEN_37790; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_37792 = 5'he == _T_3804 ? 5'h0 : _GEN_37791; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_37793 = 5'hf == _T_3804 ? w_vn_15 : _GEN_37792; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_37794 = 5'h10 == _T_3804 ? w_vn_16 : _GEN_37793; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_37795 = 5'h11 == _T_3804 ? 5'h0 : _GEN_37794; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_37796 = 5'h12 == _T_3804 ? w_vn_18 : _GEN_37795; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_37797 = 5'h13 == _T_3804 ? 5'h0 : _GEN_37796; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_37798 = 5'h14 == _T_3804 ? 5'h0 : _GEN_37797; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_37799 = 5'h15 == _T_3804 ? 5'h0 : _GEN_37798; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_37800 = 5'h16 == _T_3804 ? 5'h0 : _GEN_37799; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_37801 = 5'h17 == _T_3804 ? w_vn_23 : _GEN_37800; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_37802 = 5'h18 == _T_3804 ? w_vn_24 : _GEN_37801; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_37803 = 5'h19 == _T_3804 ? 5'h0 : _GEN_37802; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_37804 = 5'h1a == _T_3804 ? 5'h0 : _GEN_37803; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_37805 = 5'h1b == _T_3804 ? 5'h0 : _GEN_37804; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_37806 = 5'h1c == _T_3804 ? 5'h0 : _GEN_37805; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_37807 = 5'h1d == _T_3804 ? 5'h0 : _GEN_37806; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_37808 = 5'h1e == _T_3804 ? 5'h0 : _GEN_37807; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_37809 = 5'h1f == _T_3804 ? 5'h0 : _GEN_37808; // @[FanCtrl.scala 168:{37,37}]
  wire  _T_3808 = _GEN_37809 != _GEN_37777; // @[FanCtrl.scala 168:37]
  wire  _T_3816 = _GEN_37524 != _GEN_37556; // @[FanCtrl.scala 169:37]
  wire  _T_3834 = _T_3800 & _T_3808; // @[FanCtrl.scala 173:71]
  wire  _T_3842 = _T_3834 & _T_3816; // @[FanCtrl.scala 174:71]
  wire  _GEN_38523 = r_valid_1 & _T_3782; // @[FanCtrl.scala 159:32]
  wire [4:0] _T_3905 = _T_3776 - 5'h1; // @[FanCtrl.scala 203:56]
  wire [4:0] _GEN_38949 = 5'h3 == _T_3905 ? w_vn_3 : 5'h0; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_38950 = 5'h4 == _T_3905 ? w_vn_4 : _GEN_38949; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_38951 = 5'h5 == _T_3905 ? 5'h0 : _GEN_38950; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_38952 = 5'h6 == _T_3905 ? 5'h0 : _GEN_38951; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_38953 = 5'h7 == _T_3905 ? w_vn_7 : _GEN_38952; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_38954 = 5'h8 == _T_3905 ? w_vn_8 : _GEN_38953; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_38955 = 5'h9 == _T_3905 ? 5'h0 : _GEN_38954; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_38956 = 5'ha == _T_3905 ? 5'h0 : _GEN_38955; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_38957 = 5'hb == _T_3905 ? w_vn_11 : _GEN_38956; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_38958 = 5'hc == _T_3905 ? w_vn_12 : _GEN_38957; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_38959 = 5'hd == _T_3905 ? w_vn_13 : _GEN_38958; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_38960 = 5'he == _T_3905 ? 5'h0 : _GEN_38959; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_38961 = 5'hf == _T_3905 ? w_vn_15 : _GEN_38960; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_38962 = 5'h10 == _T_3905 ? w_vn_16 : _GEN_38961; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_38963 = 5'h11 == _T_3905 ? 5'h0 : _GEN_38962; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_38964 = 5'h12 == _T_3905 ? w_vn_18 : _GEN_38963; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_38965 = 5'h13 == _T_3905 ? 5'h0 : _GEN_38964; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_38966 = 5'h14 == _T_3905 ? 5'h0 : _GEN_38965; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_38967 = 5'h15 == _T_3905 ? 5'h0 : _GEN_38966; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_38968 = 5'h16 == _T_3905 ? 5'h0 : _GEN_38967; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_38969 = 5'h17 == _T_3905 ? w_vn_23 : _GEN_38968; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_38970 = 5'h18 == _T_3905 ? w_vn_24 : _GEN_38969; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_38971 = 5'h19 == _T_3905 ? 5'h0 : _GEN_38970; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_38972 = 5'h1a == _T_3905 ? 5'h0 : _GEN_38971; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_38973 = 5'h1b == _T_3905 ? 5'h0 : _GEN_38972; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_38974 = 5'h1c == _T_3905 ? 5'h0 : _GEN_38973; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_38975 = 5'h1d == _T_3905 ? 5'h0 : _GEN_38974; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_38976 = 5'h1e == _T_3905 ? 5'h0 : _GEN_38975; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_38977 = 5'h1f == _T_3905 ? 5'h0 : _GEN_38976; // @[FanCtrl.scala 203:{37,37}]
  wire  _T_3906 = _GEN_37681 != _GEN_38977; // @[FanCtrl.scala 203:37]
  wire  _T_3907 = _T_3801 & _T_3906; // @[FanCtrl.scala 202:65]
  wire  _T_3932 = _T_3793 & _T_3906; // @[FanCtrl.scala 208:71]
  wire  _T_3940 = _T_3932 & _T_3816; // @[FanCtrl.scala 209:70]
  wire  _T_4012 = _T_3907 & _T_3808; // @[FanCtrl.scala 239:64]
  wire  _T_4020 = _T_4012 & _T_3816; // @[FanCtrl.scala 240:62]
  wire [2:0] _GEN_40768 = _T_3940 ? 3'h3 : 3'h0; // @[FanCtrl.scala 253:70]
  wire [2:0] _GEN_40799 = _T_3842 ? 3'h4 : _GEN_40768; // @[FanCtrl.scala 247:70]
  wire [2:0] _GEN_40830 = _T_4020 ? 3'h5 : _GEN_40799; // @[FanCtrl.scala 241:64]
  wire [2:0] _GEN_40954 = r_valid_1 ? _GEN_40830 : 3'h0; // @[FanCtrl.scala 230:30]
  wire [4:0] _T_4085 = 3'h4 * 2'h3; // @[FanCtrl.scala 160:23]
  wire [4:0] _T_4087 = _T_4085 + 5'h1; // @[FanCtrl.scala 160:29]
  wire [4:0] _T_4090 = _T_4085 + 5'h2; // @[FanCtrl.scala 160:56]
  wire [4:0] _GEN_41156 = 5'h3 == _T_4087 ? w_vn_3 : 5'h0; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_41157 = 5'h4 == _T_4087 ? w_vn_4 : _GEN_41156; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_41158 = 5'h5 == _T_4087 ? 5'h0 : _GEN_41157; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_41159 = 5'h6 == _T_4087 ? 5'h0 : _GEN_41158; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_41160 = 5'h7 == _T_4087 ? w_vn_7 : _GEN_41159; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_41161 = 5'h8 == _T_4087 ? w_vn_8 : _GEN_41160; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_41162 = 5'h9 == _T_4087 ? 5'h0 : _GEN_41161; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_41163 = 5'ha == _T_4087 ? 5'h0 : _GEN_41162; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_41164 = 5'hb == _T_4087 ? w_vn_11 : _GEN_41163; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_41165 = 5'hc == _T_4087 ? w_vn_12 : _GEN_41164; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_41166 = 5'hd == _T_4087 ? w_vn_13 : _GEN_41165; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_41167 = 5'he == _T_4087 ? 5'h0 : _GEN_41166; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_41168 = 5'hf == _T_4087 ? w_vn_15 : _GEN_41167; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_41169 = 5'h10 == _T_4087 ? w_vn_16 : _GEN_41168; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_41170 = 5'h11 == _T_4087 ? 5'h0 : _GEN_41169; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_41171 = 5'h12 == _T_4087 ? w_vn_18 : _GEN_41170; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_41172 = 5'h13 == _T_4087 ? 5'h0 : _GEN_41171; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_41173 = 5'h14 == _T_4087 ? 5'h0 : _GEN_41172; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_41174 = 5'h15 == _T_4087 ? 5'h0 : _GEN_41173; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_41175 = 5'h16 == _T_4087 ? 5'h0 : _GEN_41174; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_41176 = 5'h17 == _T_4087 ? w_vn_23 : _GEN_41175; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_41177 = 5'h18 == _T_4087 ? w_vn_24 : _GEN_41176; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_41178 = 5'h19 == _T_4087 ? 5'h0 : _GEN_41177; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_41179 = 5'h1a == _T_4087 ? 5'h0 : _GEN_41178; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_41180 = 5'h1b == _T_4087 ? 5'h0 : _GEN_41179; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_41181 = 5'h1c == _T_4087 ? 5'h0 : _GEN_41180; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_41182 = 5'h1d == _T_4087 ? 5'h0 : _GEN_41181; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_41183 = 5'h1e == _T_4087 ? 5'h0 : _GEN_41182; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_41184 = 5'h1f == _T_4087 ? 5'h0 : _GEN_41183; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_41188 = 5'h3 == _T_4090 ? w_vn_3 : 5'h0; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_41189 = 5'h4 == _T_4090 ? w_vn_4 : _GEN_41188; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_41190 = 5'h5 == _T_4090 ? 5'h0 : _GEN_41189; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_41191 = 5'h6 == _T_4090 ? 5'h0 : _GEN_41190; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_41192 = 5'h7 == _T_4090 ? w_vn_7 : _GEN_41191; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_41193 = 5'h8 == _T_4090 ? w_vn_8 : _GEN_41192; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_41194 = 5'h9 == _T_4090 ? 5'h0 : _GEN_41193; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_41195 = 5'ha == _T_4090 ? 5'h0 : _GEN_41194; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_41196 = 5'hb == _T_4090 ? w_vn_11 : _GEN_41195; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_41197 = 5'hc == _T_4090 ? w_vn_12 : _GEN_41196; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_41198 = 5'hd == _T_4090 ? w_vn_13 : _GEN_41197; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_41199 = 5'he == _T_4090 ? 5'h0 : _GEN_41198; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_41200 = 5'hf == _T_4090 ? w_vn_15 : _GEN_41199; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_41201 = 5'h10 == _T_4090 ? w_vn_16 : _GEN_41200; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_41202 = 5'h11 == _T_4090 ? 5'h0 : _GEN_41201; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_41203 = 5'h12 == _T_4090 ? w_vn_18 : _GEN_41202; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_41204 = 5'h13 == _T_4090 ? 5'h0 : _GEN_41203; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_41205 = 5'h14 == _T_4090 ? 5'h0 : _GEN_41204; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_41206 = 5'h15 == _T_4090 ? 5'h0 : _GEN_41205; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_41207 = 5'h16 == _T_4090 ? 5'h0 : _GEN_41206; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_41208 = 5'h17 == _T_4090 ? w_vn_23 : _GEN_41207; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_41209 = 5'h18 == _T_4090 ? w_vn_24 : _GEN_41208; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_41210 = 5'h19 == _T_4090 ? 5'h0 : _GEN_41209; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_41211 = 5'h1a == _T_4090 ? 5'h0 : _GEN_41210; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_41212 = 5'h1b == _T_4090 ? 5'h0 : _GEN_41211; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_41213 = 5'h1c == _T_4090 ? 5'h0 : _GEN_41212; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_41214 = 5'h1d == _T_4090 ? 5'h0 : _GEN_41213; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_41215 = 5'h1e == _T_4090 ? 5'h0 : _GEN_41214; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_41216 = 5'h1f == _T_4090 ? 5'h0 : _GEN_41215; // @[FanCtrl.scala 160:{37,37}]
  wire  _T_4091 = _GEN_41184 == _GEN_41216; // @[FanCtrl.scala 160:37]
  wire [5:0] _T_4097 = {{1'd0}, _T_4085}; // @[FanCtrl.scala 166:30]
  wire [4:0] _GEN_41313 = 5'h3 == _T_4097[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_41314 = 5'h4 == _T_4097[4:0] ? w_vn_4 : _GEN_41313; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_41315 = 5'h5 == _T_4097[4:0] ? 5'h0 : _GEN_41314; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_41316 = 5'h6 == _T_4097[4:0] ? 5'h0 : _GEN_41315; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_41317 = 5'h7 == _T_4097[4:0] ? w_vn_7 : _GEN_41316; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_41318 = 5'h8 == _T_4097[4:0] ? w_vn_8 : _GEN_41317; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_41319 = 5'h9 == _T_4097[4:0] ? 5'h0 : _GEN_41318; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_41320 = 5'ha == _T_4097[4:0] ? 5'h0 : _GEN_41319; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_41321 = 5'hb == _T_4097[4:0] ? w_vn_11 : _GEN_41320; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_41322 = 5'hc == _T_4097[4:0] ? w_vn_12 : _GEN_41321; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_41323 = 5'hd == _T_4097[4:0] ? w_vn_13 : _GEN_41322; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_41324 = 5'he == _T_4097[4:0] ? 5'h0 : _GEN_41323; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_41325 = 5'hf == _T_4097[4:0] ? w_vn_15 : _GEN_41324; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_41326 = 5'h10 == _T_4097[4:0] ? w_vn_16 : _GEN_41325; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_41327 = 5'h11 == _T_4097[4:0] ? 5'h0 : _GEN_41326; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_41328 = 5'h12 == _T_4097[4:0] ? w_vn_18 : _GEN_41327; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_41329 = 5'h13 == _T_4097[4:0] ? 5'h0 : _GEN_41328; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_41330 = 5'h14 == _T_4097[4:0] ? 5'h0 : _GEN_41329; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_41331 = 5'h15 == _T_4097[4:0] ? 5'h0 : _GEN_41330; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_41332 = 5'h16 == _T_4097[4:0] ? 5'h0 : _GEN_41331; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_41333 = 5'h17 == _T_4097[4:0] ? w_vn_23 : _GEN_41332; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_41334 = 5'h18 == _T_4097[4:0] ? w_vn_24 : _GEN_41333; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_41335 = 5'h19 == _T_4097[4:0] ? 5'h0 : _GEN_41334; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_41336 = 5'h1a == _T_4097[4:0] ? 5'h0 : _GEN_41335; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_41337 = 5'h1b == _T_4097[4:0] ? 5'h0 : _GEN_41336; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_41338 = 5'h1c == _T_4097[4:0] ? 5'h0 : _GEN_41337; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_41339 = 5'h1d == _T_4097[4:0] ? 5'h0 : _GEN_41338; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_41340 = 5'h1e == _T_4097[4:0] ? 5'h0 : _GEN_41339; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_41341 = 5'h1f == _T_4097[4:0] ? 5'h0 : _GEN_41340; // @[FanCtrl.scala 166:{38,38}]
  wire  _T_4102 = _GEN_41341 == _GEN_41184; // @[FanCtrl.scala 166:38]
  wire [4:0] _T_4108 = _T_4085 + 5'h3; // @[FanCtrl.scala 167:55]
  wire [4:0] _GEN_41409 = 5'h3 == _T_4108 ? w_vn_3 : 5'h0; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_41410 = 5'h4 == _T_4108 ? w_vn_4 : _GEN_41409; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_41411 = 5'h5 == _T_4108 ? 5'h0 : _GEN_41410; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_41412 = 5'h6 == _T_4108 ? 5'h0 : _GEN_41411; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_41413 = 5'h7 == _T_4108 ? w_vn_7 : _GEN_41412; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_41414 = 5'h8 == _T_4108 ? w_vn_8 : _GEN_41413; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_41415 = 5'h9 == _T_4108 ? 5'h0 : _GEN_41414; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_41416 = 5'ha == _T_4108 ? 5'h0 : _GEN_41415; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_41417 = 5'hb == _T_4108 ? w_vn_11 : _GEN_41416; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_41418 = 5'hc == _T_4108 ? w_vn_12 : _GEN_41417; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_41419 = 5'hd == _T_4108 ? w_vn_13 : _GEN_41418; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_41420 = 5'he == _T_4108 ? 5'h0 : _GEN_41419; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_41421 = 5'hf == _T_4108 ? w_vn_15 : _GEN_41420; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_41422 = 5'h10 == _T_4108 ? w_vn_16 : _GEN_41421; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_41423 = 5'h11 == _T_4108 ? 5'h0 : _GEN_41422; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_41424 = 5'h12 == _T_4108 ? w_vn_18 : _GEN_41423; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_41425 = 5'h13 == _T_4108 ? 5'h0 : _GEN_41424; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_41426 = 5'h14 == _T_4108 ? 5'h0 : _GEN_41425; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_41427 = 5'h15 == _T_4108 ? 5'h0 : _GEN_41426; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_41428 = 5'h16 == _T_4108 ? 5'h0 : _GEN_41427; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_41429 = 5'h17 == _T_4108 ? w_vn_23 : _GEN_41428; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_41430 = 5'h18 == _T_4108 ? w_vn_24 : _GEN_41429; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_41431 = 5'h19 == _T_4108 ? 5'h0 : _GEN_41430; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_41432 = 5'h1a == _T_4108 ? 5'h0 : _GEN_41431; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_41433 = 5'h1b == _T_4108 ? 5'h0 : _GEN_41432; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_41434 = 5'h1c == _T_4108 ? 5'h0 : _GEN_41433; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_41435 = 5'h1d == _T_4108 ? 5'h0 : _GEN_41434; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_41436 = 5'h1e == _T_4108 ? 5'h0 : _GEN_41435; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_41437 = 5'h1f == _T_4108 ? 5'h0 : _GEN_41436; // @[FanCtrl.scala 167:{36,36}]
  wire  _T_4109 = _GEN_41216 == _GEN_41437; // @[FanCtrl.scala 167:36]
  wire  _T_4110 = _GEN_41341 == _GEN_41184 & _T_4109; // @[FanCtrl.scala 166:65]
  wire [4:0] _T_4113 = _T_4085 + 5'h4; // @[FanCtrl.scala 168:29]
  wire [4:0] _GEN_41441 = 5'h3 == _T_4113 ? w_vn_3 : 5'h0; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_41442 = 5'h4 == _T_4113 ? w_vn_4 : _GEN_41441; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_41443 = 5'h5 == _T_4113 ? 5'h0 : _GEN_41442; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_41444 = 5'h6 == _T_4113 ? 5'h0 : _GEN_41443; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_41445 = 5'h7 == _T_4113 ? w_vn_7 : _GEN_41444; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_41446 = 5'h8 == _T_4113 ? w_vn_8 : _GEN_41445; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_41447 = 5'h9 == _T_4113 ? 5'h0 : _GEN_41446; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_41448 = 5'ha == _T_4113 ? 5'h0 : _GEN_41447; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_41449 = 5'hb == _T_4113 ? w_vn_11 : _GEN_41448; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_41450 = 5'hc == _T_4113 ? w_vn_12 : _GEN_41449; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_41451 = 5'hd == _T_4113 ? w_vn_13 : _GEN_41450; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_41452 = 5'he == _T_4113 ? 5'h0 : _GEN_41451; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_41453 = 5'hf == _T_4113 ? w_vn_15 : _GEN_41452; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_41454 = 5'h10 == _T_4113 ? w_vn_16 : _GEN_41453; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_41455 = 5'h11 == _T_4113 ? 5'h0 : _GEN_41454; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_41456 = 5'h12 == _T_4113 ? w_vn_18 : _GEN_41455; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_41457 = 5'h13 == _T_4113 ? 5'h0 : _GEN_41456; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_41458 = 5'h14 == _T_4113 ? 5'h0 : _GEN_41457; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_41459 = 5'h15 == _T_4113 ? 5'h0 : _GEN_41458; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_41460 = 5'h16 == _T_4113 ? 5'h0 : _GEN_41459; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_41461 = 5'h17 == _T_4113 ? w_vn_23 : _GEN_41460; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_41462 = 5'h18 == _T_4113 ? w_vn_24 : _GEN_41461; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_41463 = 5'h19 == _T_4113 ? 5'h0 : _GEN_41462; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_41464 = 5'h1a == _T_4113 ? 5'h0 : _GEN_41463; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_41465 = 5'h1b == _T_4113 ? 5'h0 : _GEN_41464; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_41466 = 5'h1c == _T_4113 ? 5'h0 : _GEN_41465; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_41467 = 5'h1d == _T_4113 ? 5'h0 : _GEN_41466; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_41468 = 5'h1e == _T_4113 ? 5'h0 : _GEN_41467; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_41469 = 5'h1f == _T_4113 ? 5'h0 : _GEN_41468; // @[FanCtrl.scala 168:{37,37}]
  wire  _T_4117 = _GEN_41469 != _GEN_41437; // @[FanCtrl.scala 168:37]
  wire  _T_4125 = _GEN_41184 != _GEN_41216; // @[FanCtrl.scala 169:37]
  wire  _T_4143 = _T_4109 & _T_4117; // @[FanCtrl.scala 173:71]
  wire  _T_4151 = _T_4143 & _T_4125; // @[FanCtrl.scala 174:71]
  wire  _GEN_42184 = r_valid_1 & _T_4091; // @[FanCtrl.scala 159:32]
  wire [4:0] _T_4214 = _T_4085 - 5'h1; // @[FanCtrl.scala 203:56]
  wire [4:0] _GEN_42609 = 5'h3 == _T_4214 ? w_vn_3 : 5'h0; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_42610 = 5'h4 == _T_4214 ? w_vn_4 : _GEN_42609; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_42611 = 5'h5 == _T_4214 ? 5'h0 : _GEN_42610; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_42612 = 5'h6 == _T_4214 ? 5'h0 : _GEN_42611; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_42613 = 5'h7 == _T_4214 ? w_vn_7 : _GEN_42612; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_42614 = 5'h8 == _T_4214 ? w_vn_8 : _GEN_42613; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_42615 = 5'h9 == _T_4214 ? 5'h0 : _GEN_42614; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_42616 = 5'ha == _T_4214 ? 5'h0 : _GEN_42615; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_42617 = 5'hb == _T_4214 ? w_vn_11 : _GEN_42616; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_42618 = 5'hc == _T_4214 ? w_vn_12 : _GEN_42617; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_42619 = 5'hd == _T_4214 ? w_vn_13 : _GEN_42618; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_42620 = 5'he == _T_4214 ? 5'h0 : _GEN_42619; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_42621 = 5'hf == _T_4214 ? w_vn_15 : _GEN_42620; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_42622 = 5'h10 == _T_4214 ? w_vn_16 : _GEN_42621; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_42623 = 5'h11 == _T_4214 ? 5'h0 : _GEN_42622; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_42624 = 5'h12 == _T_4214 ? w_vn_18 : _GEN_42623; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_42625 = 5'h13 == _T_4214 ? 5'h0 : _GEN_42624; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_42626 = 5'h14 == _T_4214 ? 5'h0 : _GEN_42625; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_42627 = 5'h15 == _T_4214 ? 5'h0 : _GEN_42626; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_42628 = 5'h16 == _T_4214 ? 5'h0 : _GEN_42627; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_42629 = 5'h17 == _T_4214 ? w_vn_23 : _GEN_42628; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_42630 = 5'h18 == _T_4214 ? w_vn_24 : _GEN_42629; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_42631 = 5'h19 == _T_4214 ? 5'h0 : _GEN_42630; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_42632 = 5'h1a == _T_4214 ? 5'h0 : _GEN_42631; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_42633 = 5'h1b == _T_4214 ? 5'h0 : _GEN_42632; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_42634 = 5'h1c == _T_4214 ? 5'h0 : _GEN_42633; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_42635 = 5'h1d == _T_4214 ? 5'h0 : _GEN_42634; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_42636 = 5'h1e == _T_4214 ? 5'h0 : _GEN_42635; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_42637 = 5'h1f == _T_4214 ? 5'h0 : _GEN_42636; // @[FanCtrl.scala 203:{37,37}]
  wire  _T_4215 = _GEN_41341 != _GEN_42637; // @[FanCtrl.scala 203:37]
  wire  _T_4216 = _T_4110 & _T_4215; // @[FanCtrl.scala 202:65]
  wire  _T_4241 = _T_4102 & _T_4215; // @[FanCtrl.scala 208:71]
  wire  _T_4249 = _T_4241 & _T_4125; // @[FanCtrl.scala 209:70]
  wire  _T_4321 = _T_4216 & _T_4117; // @[FanCtrl.scala 239:64]
  wire  _T_4329 = _T_4321 & _T_4125; // @[FanCtrl.scala 240:62]
  wire [2:0] _GEN_44429 = _T_4249 ? 3'h3 : 3'h0; // @[FanCtrl.scala 253:70]
  wire [2:0] _GEN_44460 = _T_4151 ? 3'h4 : _GEN_44429; // @[FanCtrl.scala 247:70]
  wire [2:0] _GEN_44491 = _T_4329 ? 3'h5 : _GEN_44460; // @[FanCtrl.scala 241:64]
  wire [2:0] _GEN_44615 = r_valid_1 ? _GEN_44491 : 3'h0; // @[FanCtrl.scala 230:30]
  wire [5:0] _T_4394 = 3'h4 * 3'h4; // @[FanCtrl.scala 160:23]
  wire [5:0] _T_4396 = _T_4394 + 6'h1; // @[FanCtrl.scala 160:29]
  wire [5:0] _T_4400 = _T_4394 + 6'h2; // @[FanCtrl.scala 160:56]
  wire [4:0] _GEN_44816 = 5'h3 == _T_4396[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_44817 = 5'h4 == _T_4396[4:0] ? w_vn_4 : _GEN_44816; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_44818 = 5'h5 == _T_4396[4:0] ? 5'h0 : _GEN_44817; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_44819 = 5'h6 == _T_4396[4:0] ? 5'h0 : _GEN_44818; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_44820 = 5'h7 == _T_4396[4:0] ? w_vn_7 : _GEN_44819; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_44821 = 5'h8 == _T_4396[4:0] ? w_vn_8 : _GEN_44820; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_44822 = 5'h9 == _T_4396[4:0] ? 5'h0 : _GEN_44821; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_44823 = 5'ha == _T_4396[4:0] ? 5'h0 : _GEN_44822; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_44824 = 5'hb == _T_4396[4:0] ? w_vn_11 : _GEN_44823; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_44825 = 5'hc == _T_4396[4:0] ? w_vn_12 : _GEN_44824; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_44826 = 5'hd == _T_4396[4:0] ? w_vn_13 : _GEN_44825; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_44827 = 5'he == _T_4396[4:0] ? 5'h0 : _GEN_44826; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_44828 = 5'hf == _T_4396[4:0] ? w_vn_15 : _GEN_44827; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_44829 = 5'h10 == _T_4396[4:0] ? w_vn_16 : _GEN_44828; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_44830 = 5'h11 == _T_4396[4:0] ? 5'h0 : _GEN_44829; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_44831 = 5'h12 == _T_4396[4:0] ? w_vn_18 : _GEN_44830; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_44832 = 5'h13 == _T_4396[4:0] ? 5'h0 : _GEN_44831; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_44833 = 5'h14 == _T_4396[4:0] ? 5'h0 : _GEN_44832; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_44834 = 5'h15 == _T_4396[4:0] ? 5'h0 : _GEN_44833; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_44835 = 5'h16 == _T_4396[4:0] ? 5'h0 : _GEN_44834; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_44836 = 5'h17 == _T_4396[4:0] ? w_vn_23 : _GEN_44835; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_44837 = 5'h18 == _T_4396[4:0] ? w_vn_24 : _GEN_44836; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_44838 = 5'h19 == _T_4396[4:0] ? 5'h0 : _GEN_44837; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_44839 = 5'h1a == _T_4396[4:0] ? 5'h0 : _GEN_44838; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_44840 = 5'h1b == _T_4396[4:0] ? 5'h0 : _GEN_44839; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_44841 = 5'h1c == _T_4396[4:0] ? 5'h0 : _GEN_44840; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_44842 = 5'h1d == _T_4396[4:0] ? 5'h0 : _GEN_44841; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_44843 = 5'h1e == _T_4396[4:0] ? 5'h0 : _GEN_44842; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_44844 = 5'h1f == _T_4396[4:0] ? 5'h0 : _GEN_44843; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_44848 = 5'h3 == _T_4400[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_44849 = 5'h4 == _T_4400[4:0] ? w_vn_4 : _GEN_44848; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_44850 = 5'h5 == _T_4400[4:0] ? 5'h0 : _GEN_44849; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_44851 = 5'h6 == _T_4400[4:0] ? 5'h0 : _GEN_44850; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_44852 = 5'h7 == _T_4400[4:0] ? w_vn_7 : _GEN_44851; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_44853 = 5'h8 == _T_4400[4:0] ? w_vn_8 : _GEN_44852; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_44854 = 5'h9 == _T_4400[4:0] ? 5'h0 : _GEN_44853; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_44855 = 5'ha == _T_4400[4:0] ? 5'h0 : _GEN_44854; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_44856 = 5'hb == _T_4400[4:0] ? w_vn_11 : _GEN_44855; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_44857 = 5'hc == _T_4400[4:0] ? w_vn_12 : _GEN_44856; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_44858 = 5'hd == _T_4400[4:0] ? w_vn_13 : _GEN_44857; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_44859 = 5'he == _T_4400[4:0] ? 5'h0 : _GEN_44858; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_44860 = 5'hf == _T_4400[4:0] ? w_vn_15 : _GEN_44859; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_44861 = 5'h10 == _T_4400[4:0] ? w_vn_16 : _GEN_44860; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_44862 = 5'h11 == _T_4400[4:0] ? 5'h0 : _GEN_44861; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_44863 = 5'h12 == _T_4400[4:0] ? w_vn_18 : _GEN_44862; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_44864 = 5'h13 == _T_4400[4:0] ? 5'h0 : _GEN_44863; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_44865 = 5'h14 == _T_4400[4:0] ? 5'h0 : _GEN_44864; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_44866 = 5'h15 == _T_4400[4:0] ? 5'h0 : _GEN_44865; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_44867 = 5'h16 == _T_4400[4:0] ? 5'h0 : _GEN_44866; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_44868 = 5'h17 == _T_4400[4:0] ? w_vn_23 : _GEN_44867; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_44869 = 5'h18 == _T_4400[4:0] ? w_vn_24 : _GEN_44868; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_44870 = 5'h19 == _T_4400[4:0] ? 5'h0 : _GEN_44869; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_44871 = 5'h1a == _T_4400[4:0] ? 5'h0 : _GEN_44870; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_44872 = 5'h1b == _T_4400[4:0] ? 5'h0 : _GEN_44871; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_44873 = 5'h1c == _T_4400[4:0] ? 5'h0 : _GEN_44872; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_44874 = 5'h1d == _T_4400[4:0] ? 5'h0 : _GEN_44873; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_44875 = 5'h1e == _T_4400[4:0] ? 5'h0 : _GEN_44874; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_44876 = 5'h1f == _T_4400[4:0] ? 5'h0 : _GEN_44875; // @[FanCtrl.scala 160:{37,37}]
  wire  _T_4402 = _GEN_44844 == _GEN_44876; // @[FanCtrl.scala 160:37]
  wire [6:0] _T_4408 = {{1'd0}, _T_4394}; // @[FanCtrl.scala 166:30]
  wire [4:0] _GEN_44973 = 5'h3 == _T_4408[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_44974 = 5'h4 == _T_4408[4:0] ? w_vn_4 : _GEN_44973; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_44975 = 5'h5 == _T_4408[4:0] ? 5'h0 : _GEN_44974; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_44976 = 5'h6 == _T_4408[4:0] ? 5'h0 : _GEN_44975; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_44977 = 5'h7 == _T_4408[4:0] ? w_vn_7 : _GEN_44976; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_44978 = 5'h8 == _T_4408[4:0] ? w_vn_8 : _GEN_44977; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_44979 = 5'h9 == _T_4408[4:0] ? 5'h0 : _GEN_44978; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_44980 = 5'ha == _T_4408[4:0] ? 5'h0 : _GEN_44979; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_44981 = 5'hb == _T_4408[4:0] ? w_vn_11 : _GEN_44980; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_44982 = 5'hc == _T_4408[4:0] ? w_vn_12 : _GEN_44981; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_44983 = 5'hd == _T_4408[4:0] ? w_vn_13 : _GEN_44982; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_44984 = 5'he == _T_4408[4:0] ? 5'h0 : _GEN_44983; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_44985 = 5'hf == _T_4408[4:0] ? w_vn_15 : _GEN_44984; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_44986 = 5'h10 == _T_4408[4:0] ? w_vn_16 : _GEN_44985; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_44987 = 5'h11 == _T_4408[4:0] ? 5'h0 : _GEN_44986; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_44988 = 5'h12 == _T_4408[4:0] ? w_vn_18 : _GEN_44987; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_44989 = 5'h13 == _T_4408[4:0] ? 5'h0 : _GEN_44988; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_44990 = 5'h14 == _T_4408[4:0] ? 5'h0 : _GEN_44989; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_44991 = 5'h15 == _T_4408[4:0] ? 5'h0 : _GEN_44990; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_44992 = 5'h16 == _T_4408[4:0] ? 5'h0 : _GEN_44991; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_44993 = 5'h17 == _T_4408[4:0] ? w_vn_23 : _GEN_44992; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_44994 = 5'h18 == _T_4408[4:0] ? w_vn_24 : _GEN_44993; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_44995 = 5'h19 == _T_4408[4:0] ? 5'h0 : _GEN_44994; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_44996 = 5'h1a == _T_4408[4:0] ? 5'h0 : _GEN_44995; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_44997 = 5'h1b == _T_4408[4:0] ? 5'h0 : _GEN_44996; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_44998 = 5'h1c == _T_4408[4:0] ? 5'h0 : _GEN_44997; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_44999 = 5'h1d == _T_4408[4:0] ? 5'h0 : _GEN_44998; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_45000 = 5'h1e == _T_4408[4:0] ? 5'h0 : _GEN_44999; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_45001 = 5'h1f == _T_4408[4:0] ? 5'h0 : _GEN_45000; // @[FanCtrl.scala 166:{38,38}]
  wire  _T_4415 = _GEN_45001 == _GEN_44844; // @[FanCtrl.scala 166:38]
  wire [5:0] _T_4422 = _T_4394 + 6'h3; // @[FanCtrl.scala 167:55]
  wire [4:0] _GEN_45069 = 5'h3 == _T_4422[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_45070 = 5'h4 == _T_4422[4:0] ? w_vn_4 : _GEN_45069; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_45071 = 5'h5 == _T_4422[4:0] ? 5'h0 : _GEN_45070; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_45072 = 5'h6 == _T_4422[4:0] ? 5'h0 : _GEN_45071; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_45073 = 5'h7 == _T_4422[4:0] ? w_vn_7 : _GEN_45072; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_45074 = 5'h8 == _T_4422[4:0] ? w_vn_8 : _GEN_45073; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_45075 = 5'h9 == _T_4422[4:0] ? 5'h0 : _GEN_45074; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_45076 = 5'ha == _T_4422[4:0] ? 5'h0 : _GEN_45075; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_45077 = 5'hb == _T_4422[4:0] ? w_vn_11 : _GEN_45076; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_45078 = 5'hc == _T_4422[4:0] ? w_vn_12 : _GEN_45077; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_45079 = 5'hd == _T_4422[4:0] ? w_vn_13 : _GEN_45078; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_45080 = 5'he == _T_4422[4:0] ? 5'h0 : _GEN_45079; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_45081 = 5'hf == _T_4422[4:0] ? w_vn_15 : _GEN_45080; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_45082 = 5'h10 == _T_4422[4:0] ? w_vn_16 : _GEN_45081; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_45083 = 5'h11 == _T_4422[4:0] ? 5'h0 : _GEN_45082; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_45084 = 5'h12 == _T_4422[4:0] ? w_vn_18 : _GEN_45083; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_45085 = 5'h13 == _T_4422[4:0] ? 5'h0 : _GEN_45084; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_45086 = 5'h14 == _T_4422[4:0] ? 5'h0 : _GEN_45085; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_45087 = 5'h15 == _T_4422[4:0] ? 5'h0 : _GEN_45086; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_45088 = 5'h16 == _T_4422[4:0] ? 5'h0 : _GEN_45087; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_45089 = 5'h17 == _T_4422[4:0] ? w_vn_23 : _GEN_45088; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_45090 = 5'h18 == _T_4422[4:0] ? w_vn_24 : _GEN_45089; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_45091 = 5'h19 == _T_4422[4:0] ? 5'h0 : _GEN_45090; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_45092 = 5'h1a == _T_4422[4:0] ? 5'h0 : _GEN_45091; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_45093 = 5'h1b == _T_4422[4:0] ? 5'h0 : _GEN_45092; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_45094 = 5'h1c == _T_4422[4:0] ? 5'h0 : _GEN_45093; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_45095 = 5'h1d == _T_4422[4:0] ? 5'h0 : _GEN_45094; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_45096 = 5'h1e == _T_4422[4:0] ? 5'h0 : _GEN_45095; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_45097 = 5'h1f == _T_4422[4:0] ? 5'h0 : _GEN_45096; // @[FanCtrl.scala 167:{36,36}]
  wire  _T_4424 = _GEN_44876 == _GEN_45097; // @[FanCtrl.scala 167:36]
  wire  _T_4425 = _GEN_45001 == _GEN_44844 & _T_4424; // @[FanCtrl.scala 166:65]
  wire [5:0] _T_4428 = _T_4394 + 6'h4; // @[FanCtrl.scala 168:29]
  wire [4:0] _GEN_45101 = 5'h3 == _T_4428[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_45102 = 5'h4 == _T_4428[4:0] ? w_vn_4 : _GEN_45101; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_45103 = 5'h5 == _T_4428[4:0] ? 5'h0 : _GEN_45102; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_45104 = 5'h6 == _T_4428[4:0] ? 5'h0 : _GEN_45103; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_45105 = 5'h7 == _T_4428[4:0] ? w_vn_7 : _GEN_45104; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_45106 = 5'h8 == _T_4428[4:0] ? w_vn_8 : _GEN_45105; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_45107 = 5'h9 == _T_4428[4:0] ? 5'h0 : _GEN_45106; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_45108 = 5'ha == _T_4428[4:0] ? 5'h0 : _GEN_45107; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_45109 = 5'hb == _T_4428[4:0] ? w_vn_11 : _GEN_45108; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_45110 = 5'hc == _T_4428[4:0] ? w_vn_12 : _GEN_45109; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_45111 = 5'hd == _T_4428[4:0] ? w_vn_13 : _GEN_45110; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_45112 = 5'he == _T_4428[4:0] ? 5'h0 : _GEN_45111; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_45113 = 5'hf == _T_4428[4:0] ? w_vn_15 : _GEN_45112; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_45114 = 5'h10 == _T_4428[4:0] ? w_vn_16 : _GEN_45113; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_45115 = 5'h11 == _T_4428[4:0] ? 5'h0 : _GEN_45114; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_45116 = 5'h12 == _T_4428[4:0] ? w_vn_18 : _GEN_45115; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_45117 = 5'h13 == _T_4428[4:0] ? 5'h0 : _GEN_45116; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_45118 = 5'h14 == _T_4428[4:0] ? 5'h0 : _GEN_45117; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_45119 = 5'h15 == _T_4428[4:0] ? 5'h0 : _GEN_45118; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_45120 = 5'h16 == _T_4428[4:0] ? 5'h0 : _GEN_45119; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_45121 = 5'h17 == _T_4428[4:0] ? w_vn_23 : _GEN_45120; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_45122 = 5'h18 == _T_4428[4:0] ? w_vn_24 : _GEN_45121; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_45123 = 5'h19 == _T_4428[4:0] ? 5'h0 : _GEN_45122; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_45124 = 5'h1a == _T_4428[4:0] ? 5'h0 : _GEN_45123; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_45125 = 5'h1b == _T_4428[4:0] ? 5'h0 : _GEN_45124; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_45126 = 5'h1c == _T_4428[4:0] ? 5'h0 : _GEN_45125; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_45127 = 5'h1d == _T_4428[4:0] ? 5'h0 : _GEN_45126; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_45128 = 5'h1e == _T_4428[4:0] ? 5'h0 : _GEN_45127; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_45129 = 5'h1f == _T_4428[4:0] ? 5'h0 : _GEN_45128; // @[FanCtrl.scala 168:{37,37}]
  wire  _T_4434 = _GEN_45129 != _GEN_45097; // @[FanCtrl.scala 168:37]
  wire  _T_4444 = _GEN_44844 != _GEN_44876; // @[FanCtrl.scala 169:37]
  wire  _T_4466 = _T_4424 & _T_4434; // @[FanCtrl.scala 173:71]
  wire  _T_4476 = _T_4466 & _T_4444; // @[FanCtrl.scala 174:71]
  wire  _GEN_45845 = r_valid_1 & _T_4402; // @[FanCtrl.scala 159:32]
  wire [5:0] _T_4550 = _T_4394 - 6'h1; // @[FanCtrl.scala 203:56]
  wire [4:0] _GEN_46269 = 5'h3 == _T_4550[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_46270 = 5'h4 == _T_4550[4:0] ? w_vn_4 : _GEN_46269; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_46271 = 5'h5 == _T_4550[4:0] ? 5'h0 : _GEN_46270; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_46272 = 5'h6 == _T_4550[4:0] ? 5'h0 : _GEN_46271; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_46273 = 5'h7 == _T_4550[4:0] ? w_vn_7 : _GEN_46272; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_46274 = 5'h8 == _T_4550[4:0] ? w_vn_8 : _GEN_46273; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_46275 = 5'h9 == _T_4550[4:0] ? 5'h0 : _GEN_46274; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_46276 = 5'ha == _T_4550[4:0] ? 5'h0 : _GEN_46275; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_46277 = 5'hb == _T_4550[4:0] ? w_vn_11 : _GEN_46276; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_46278 = 5'hc == _T_4550[4:0] ? w_vn_12 : _GEN_46277; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_46279 = 5'hd == _T_4550[4:0] ? w_vn_13 : _GEN_46278; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_46280 = 5'he == _T_4550[4:0] ? 5'h0 : _GEN_46279; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_46281 = 5'hf == _T_4550[4:0] ? w_vn_15 : _GEN_46280; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_46282 = 5'h10 == _T_4550[4:0] ? w_vn_16 : _GEN_46281; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_46283 = 5'h11 == _T_4550[4:0] ? 5'h0 : _GEN_46282; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_46284 = 5'h12 == _T_4550[4:0] ? w_vn_18 : _GEN_46283; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_46285 = 5'h13 == _T_4550[4:0] ? 5'h0 : _GEN_46284; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_46286 = 5'h14 == _T_4550[4:0] ? 5'h0 : _GEN_46285; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_46287 = 5'h15 == _T_4550[4:0] ? 5'h0 : _GEN_46286; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_46288 = 5'h16 == _T_4550[4:0] ? 5'h0 : _GEN_46287; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_46289 = 5'h17 == _T_4550[4:0] ? w_vn_23 : _GEN_46288; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_46290 = 5'h18 == _T_4550[4:0] ? w_vn_24 : _GEN_46289; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_46291 = 5'h19 == _T_4550[4:0] ? 5'h0 : _GEN_46290; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_46292 = 5'h1a == _T_4550[4:0] ? 5'h0 : _GEN_46291; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_46293 = 5'h1b == _T_4550[4:0] ? 5'h0 : _GEN_46292; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_46294 = 5'h1c == _T_4550[4:0] ? 5'h0 : _GEN_46293; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_46295 = 5'h1d == _T_4550[4:0] ? 5'h0 : _GEN_46294; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_46296 = 5'h1e == _T_4550[4:0] ? 5'h0 : _GEN_46295; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_46297 = 5'h1f == _T_4550[4:0] ? 5'h0 : _GEN_46296; // @[FanCtrl.scala 203:{37,37}]
  wire  _T_4552 = _GEN_45001 != _GEN_46297; // @[FanCtrl.scala 203:37]
  wire  _T_4553 = _T_4425 & _T_4552; // @[FanCtrl.scala 202:65]
  wire  _T_4584 = _T_4415 & _T_4552; // @[FanCtrl.scala 208:71]
  wire  _T_4594 = _T_4584 & _T_4444; // @[FanCtrl.scala 209:70]
  wire  _T_4680 = _T_4553 & _T_4434; // @[FanCtrl.scala 239:64]
  wire  _T_4690 = _T_4680 & _T_4444; // @[FanCtrl.scala 240:62]
  wire [2:0] _GEN_48090 = _T_4594 ? 3'h3 : 3'h0; // @[FanCtrl.scala 253:70]
  wire [2:0] _GEN_48121 = _T_4476 ? 3'h4 : _GEN_48090; // @[FanCtrl.scala 247:70]
  wire [2:0] _GEN_48152 = _T_4690 ? 3'h5 : _GEN_48121; // @[FanCtrl.scala 241:64]
  wire [2:0] _GEN_48276 = r_valid_1 ? _GEN_48152 : 3'h0; // @[FanCtrl.scala 230:30]
  wire [5:0] _T_4767 = 3'h4 * 3'h5; // @[FanCtrl.scala 160:23]
  wire [5:0] _T_4769 = _T_4767 + 6'h1; // @[FanCtrl.scala 160:29]
  wire [5:0] _T_4773 = _T_4767 + 6'h2; // @[FanCtrl.scala 160:56]
  wire [4:0] _GEN_48476 = 5'h3 == _T_4769[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_48477 = 5'h4 == _T_4769[4:0] ? w_vn_4 : _GEN_48476; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_48478 = 5'h5 == _T_4769[4:0] ? 5'h0 : _GEN_48477; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_48479 = 5'h6 == _T_4769[4:0] ? 5'h0 : _GEN_48478; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_48480 = 5'h7 == _T_4769[4:0] ? w_vn_7 : _GEN_48479; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_48481 = 5'h8 == _T_4769[4:0] ? w_vn_8 : _GEN_48480; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_48482 = 5'h9 == _T_4769[4:0] ? 5'h0 : _GEN_48481; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_48483 = 5'ha == _T_4769[4:0] ? 5'h0 : _GEN_48482; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_48484 = 5'hb == _T_4769[4:0] ? w_vn_11 : _GEN_48483; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_48485 = 5'hc == _T_4769[4:0] ? w_vn_12 : _GEN_48484; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_48486 = 5'hd == _T_4769[4:0] ? w_vn_13 : _GEN_48485; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_48487 = 5'he == _T_4769[4:0] ? 5'h0 : _GEN_48486; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_48488 = 5'hf == _T_4769[4:0] ? w_vn_15 : _GEN_48487; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_48489 = 5'h10 == _T_4769[4:0] ? w_vn_16 : _GEN_48488; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_48490 = 5'h11 == _T_4769[4:0] ? 5'h0 : _GEN_48489; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_48491 = 5'h12 == _T_4769[4:0] ? w_vn_18 : _GEN_48490; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_48492 = 5'h13 == _T_4769[4:0] ? 5'h0 : _GEN_48491; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_48493 = 5'h14 == _T_4769[4:0] ? 5'h0 : _GEN_48492; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_48494 = 5'h15 == _T_4769[4:0] ? 5'h0 : _GEN_48493; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_48495 = 5'h16 == _T_4769[4:0] ? 5'h0 : _GEN_48494; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_48496 = 5'h17 == _T_4769[4:0] ? w_vn_23 : _GEN_48495; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_48497 = 5'h18 == _T_4769[4:0] ? w_vn_24 : _GEN_48496; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_48498 = 5'h19 == _T_4769[4:0] ? 5'h0 : _GEN_48497; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_48499 = 5'h1a == _T_4769[4:0] ? 5'h0 : _GEN_48498; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_48500 = 5'h1b == _T_4769[4:0] ? 5'h0 : _GEN_48499; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_48501 = 5'h1c == _T_4769[4:0] ? 5'h0 : _GEN_48500; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_48502 = 5'h1d == _T_4769[4:0] ? 5'h0 : _GEN_48501; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_48503 = 5'h1e == _T_4769[4:0] ? 5'h0 : _GEN_48502; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_48504 = 5'h1f == _T_4769[4:0] ? 5'h0 : _GEN_48503; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_48508 = 5'h3 == _T_4773[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_48509 = 5'h4 == _T_4773[4:0] ? w_vn_4 : _GEN_48508; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_48510 = 5'h5 == _T_4773[4:0] ? 5'h0 : _GEN_48509; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_48511 = 5'h6 == _T_4773[4:0] ? 5'h0 : _GEN_48510; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_48512 = 5'h7 == _T_4773[4:0] ? w_vn_7 : _GEN_48511; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_48513 = 5'h8 == _T_4773[4:0] ? w_vn_8 : _GEN_48512; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_48514 = 5'h9 == _T_4773[4:0] ? 5'h0 : _GEN_48513; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_48515 = 5'ha == _T_4773[4:0] ? 5'h0 : _GEN_48514; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_48516 = 5'hb == _T_4773[4:0] ? w_vn_11 : _GEN_48515; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_48517 = 5'hc == _T_4773[4:0] ? w_vn_12 : _GEN_48516; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_48518 = 5'hd == _T_4773[4:0] ? w_vn_13 : _GEN_48517; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_48519 = 5'he == _T_4773[4:0] ? 5'h0 : _GEN_48518; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_48520 = 5'hf == _T_4773[4:0] ? w_vn_15 : _GEN_48519; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_48521 = 5'h10 == _T_4773[4:0] ? w_vn_16 : _GEN_48520; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_48522 = 5'h11 == _T_4773[4:0] ? 5'h0 : _GEN_48521; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_48523 = 5'h12 == _T_4773[4:0] ? w_vn_18 : _GEN_48522; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_48524 = 5'h13 == _T_4773[4:0] ? 5'h0 : _GEN_48523; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_48525 = 5'h14 == _T_4773[4:0] ? 5'h0 : _GEN_48524; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_48526 = 5'h15 == _T_4773[4:0] ? 5'h0 : _GEN_48525; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_48527 = 5'h16 == _T_4773[4:0] ? 5'h0 : _GEN_48526; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_48528 = 5'h17 == _T_4773[4:0] ? w_vn_23 : _GEN_48527; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_48529 = 5'h18 == _T_4773[4:0] ? w_vn_24 : _GEN_48528; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_48530 = 5'h19 == _T_4773[4:0] ? 5'h0 : _GEN_48529; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_48531 = 5'h1a == _T_4773[4:0] ? 5'h0 : _GEN_48530; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_48532 = 5'h1b == _T_4773[4:0] ? 5'h0 : _GEN_48531; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_48533 = 5'h1c == _T_4773[4:0] ? 5'h0 : _GEN_48532; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_48534 = 5'h1d == _T_4773[4:0] ? 5'h0 : _GEN_48533; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_48535 = 5'h1e == _T_4773[4:0] ? 5'h0 : _GEN_48534; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_48536 = 5'h1f == _T_4773[4:0] ? 5'h0 : _GEN_48535; // @[FanCtrl.scala 160:{37,37}]
  wire  _T_4775 = _GEN_48504 == _GEN_48536; // @[FanCtrl.scala 160:37]
  wire [6:0] _T_4781 = {{1'd0}, _T_4767}; // @[FanCtrl.scala 166:30]
  wire [4:0] _GEN_48633 = 5'h3 == _T_4781[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_48634 = 5'h4 == _T_4781[4:0] ? w_vn_4 : _GEN_48633; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_48635 = 5'h5 == _T_4781[4:0] ? 5'h0 : _GEN_48634; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_48636 = 5'h6 == _T_4781[4:0] ? 5'h0 : _GEN_48635; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_48637 = 5'h7 == _T_4781[4:0] ? w_vn_7 : _GEN_48636; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_48638 = 5'h8 == _T_4781[4:0] ? w_vn_8 : _GEN_48637; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_48639 = 5'h9 == _T_4781[4:0] ? 5'h0 : _GEN_48638; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_48640 = 5'ha == _T_4781[4:0] ? 5'h0 : _GEN_48639; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_48641 = 5'hb == _T_4781[4:0] ? w_vn_11 : _GEN_48640; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_48642 = 5'hc == _T_4781[4:0] ? w_vn_12 : _GEN_48641; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_48643 = 5'hd == _T_4781[4:0] ? w_vn_13 : _GEN_48642; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_48644 = 5'he == _T_4781[4:0] ? 5'h0 : _GEN_48643; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_48645 = 5'hf == _T_4781[4:0] ? w_vn_15 : _GEN_48644; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_48646 = 5'h10 == _T_4781[4:0] ? w_vn_16 : _GEN_48645; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_48647 = 5'h11 == _T_4781[4:0] ? 5'h0 : _GEN_48646; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_48648 = 5'h12 == _T_4781[4:0] ? w_vn_18 : _GEN_48647; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_48649 = 5'h13 == _T_4781[4:0] ? 5'h0 : _GEN_48648; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_48650 = 5'h14 == _T_4781[4:0] ? 5'h0 : _GEN_48649; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_48651 = 5'h15 == _T_4781[4:0] ? 5'h0 : _GEN_48650; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_48652 = 5'h16 == _T_4781[4:0] ? 5'h0 : _GEN_48651; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_48653 = 5'h17 == _T_4781[4:0] ? w_vn_23 : _GEN_48652; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_48654 = 5'h18 == _T_4781[4:0] ? w_vn_24 : _GEN_48653; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_48655 = 5'h19 == _T_4781[4:0] ? 5'h0 : _GEN_48654; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_48656 = 5'h1a == _T_4781[4:0] ? 5'h0 : _GEN_48655; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_48657 = 5'h1b == _T_4781[4:0] ? 5'h0 : _GEN_48656; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_48658 = 5'h1c == _T_4781[4:0] ? 5'h0 : _GEN_48657; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_48659 = 5'h1d == _T_4781[4:0] ? 5'h0 : _GEN_48658; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_48660 = 5'h1e == _T_4781[4:0] ? 5'h0 : _GEN_48659; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_48661 = 5'h1f == _T_4781[4:0] ? 5'h0 : _GEN_48660; // @[FanCtrl.scala 166:{38,38}]
  wire  _T_4788 = _GEN_48661 == _GEN_48504; // @[FanCtrl.scala 166:38]
  wire [5:0] _T_4795 = _T_4767 + 6'h3; // @[FanCtrl.scala 167:55]
  wire [4:0] _GEN_48729 = 5'h3 == _T_4795[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_48730 = 5'h4 == _T_4795[4:0] ? w_vn_4 : _GEN_48729; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_48731 = 5'h5 == _T_4795[4:0] ? 5'h0 : _GEN_48730; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_48732 = 5'h6 == _T_4795[4:0] ? 5'h0 : _GEN_48731; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_48733 = 5'h7 == _T_4795[4:0] ? w_vn_7 : _GEN_48732; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_48734 = 5'h8 == _T_4795[4:0] ? w_vn_8 : _GEN_48733; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_48735 = 5'h9 == _T_4795[4:0] ? 5'h0 : _GEN_48734; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_48736 = 5'ha == _T_4795[4:0] ? 5'h0 : _GEN_48735; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_48737 = 5'hb == _T_4795[4:0] ? w_vn_11 : _GEN_48736; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_48738 = 5'hc == _T_4795[4:0] ? w_vn_12 : _GEN_48737; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_48739 = 5'hd == _T_4795[4:0] ? w_vn_13 : _GEN_48738; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_48740 = 5'he == _T_4795[4:0] ? 5'h0 : _GEN_48739; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_48741 = 5'hf == _T_4795[4:0] ? w_vn_15 : _GEN_48740; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_48742 = 5'h10 == _T_4795[4:0] ? w_vn_16 : _GEN_48741; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_48743 = 5'h11 == _T_4795[4:0] ? 5'h0 : _GEN_48742; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_48744 = 5'h12 == _T_4795[4:0] ? w_vn_18 : _GEN_48743; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_48745 = 5'h13 == _T_4795[4:0] ? 5'h0 : _GEN_48744; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_48746 = 5'h14 == _T_4795[4:0] ? 5'h0 : _GEN_48745; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_48747 = 5'h15 == _T_4795[4:0] ? 5'h0 : _GEN_48746; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_48748 = 5'h16 == _T_4795[4:0] ? 5'h0 : _GEN_48747; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_48749 = 5'h17 == _T_4795[4:0] ? w_vn_23 : _GEN_48748; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_48750 = 5'h18 == _T_4795[4:0] ? w_vn_24 : _GEN_48749; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_48751 = 5'h19 == _T_4795[4:0] ? 5'h0 : _GEN_48750; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_48752 = 5'h1a == _T_4795[4:0] ? 5'h0 : _GEN_48751; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_48753 = 5'h1b == _T_4795[4:0] ? 5'h0 : _GEN_48752; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_48754 = 5'h1c == _T_4795[4:0] ? 5'h0 : _GEN_48753; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_48755 = 5'h1d == _T_4795[4:0] ? 5'h0 : _GEN_48754; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_48756 = 5'h1e == _T_4795[4:0] ? 5'h0 : _GEN_48755; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_48757 = 5'h1f == _T_4795[4:0] ? 5'h0 : _GEN_48756; // @[FanCtrl.scala 167:{36,36}]
  wire  _T_4797 = _GEN_48536 == _GEN_48757; // @[FanCtrl.scala 167:36]
  wire  _T_4798 = _GEN_48661 == _GEN_48504 & _T_4797; // @[FanCtrl.scala 166:65]
  wire [5:0] _T_4801 = _T_4767 + 6'h4; // @[FanCtrl.scala 168:29]
  wire [4:0] _GEN_48761 = 5'h3 == _T_4801[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_48762 = 5'h4 == _T_4801[4:0] ? w_vn_4 : _GEN_48761; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_48763 = 5'h5 == _T_4801[4:0] ? 5'h0 : _GEN_48762; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_48764 = 5'h6 == _T_4801[4:0] ? 5'h0 : _GEN_48763; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_48765 = 5'h7 == _T_4801[4:0] ? w_vn_7 : _GEN_48764; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_48766 = 5'h8 == _T_4801[4:0] ? w_vn_8 : _GEN_48765; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_48767 = 5'h9 == _T_4801[4:0] ? 5'h0 : _GEN_48766; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_48768 = 5'ha == _T_4801[4:0] ? 5'h0 : _GEN_48767; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_48769 = 5'hb == _T_4801[4:0] ? w_vn_11 : _GEN_48768; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_48770 = 5'hc == _T_4801[4:0] ? w_vn_12 : _GEN_48769; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_48771 = 5'hd == _T_4801[4:0] ? w_vn_13 : _GEN_48770; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_48772 = 5'he == _T_4801[4:0] ? 5'h0 : _GEN_48771; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_48773 = 5'hf == _T_4801[4:0] ? w_vn_15 : _GEN_48772; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_48774 = 5'h10 == _T_4801[4:0] ? w_vn_16 : _GEN_48773; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_48775 = 5'h11 == _T_4801[4:0] ? 5'h0 : _GEN_48774; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_48776 = 5'h12 == _T_4801[4:0] ? w_vn_18 : _GEN_48775; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_48777 = 5'h13 == _T_4801[4:0] ? 5'h0 : _GEN_48776; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_48778 = 5'h14 == _T_4801[4:0] ? 5'h0 : _GEN_48777; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_48779 = 5'h15 == _T_4801[4:0] ? 5'h0 : _GEN_48778; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_48780 = 5'h16 == _T_4801[4:0] ? 5'h0 : _GEN_48779; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_48781 = 5'h17 == _T_4801[4:0] ? w_vn_23 : _GEN_48780; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_48782 = 5'h18 == _T_4801[4:0] ? w_vn_24 : _GEN_48781; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_48783 = 5'h19 == _T_4801[4:0] ? 5'h0 : _GEN_48782; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_48784 = 5'h1a == _T_4801[4:0] ? 5'h0 : _GEN_48783; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_48785 = 5'h1b == _T_4801[4:0] ? 5'h0 : _GEN_48784; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_48786 = 5'h1c == _T_4801[4:0] ? 5'h0 : _GEN_48785; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_48787 = 5'h1d == _T_4801[4:0] ? 5'h0 : _GEN_48786; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_48788 = 5'h1e == _T_4801[4:0] ? 5'h0 : _GEN_48787; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_48789 = 5'h1f == _T_4801[4:0] ? 5'h0 : _GEN_48788; // @[FanCtrl.scala 168:{37,37}]
  wire  _T_4807 = _GEN_48789 != _GEN_48757; // @[FanCtrl.scala 168:37]
  wire  _T_4817 = _GEN_48504 != _GEN_48536; // @[FanCtrl.scala 169:37]
  wire  _T_4839 = _T_4797 & _T_4807; // @[FanCtrl.scala 173:71]
  wire  _T_4849 = _T_4839 & _T_4817; // @[FanCtrl.scala 174:71]
  wire  _GEN_49506 = r_valid_1 & _T_4775; // @[FanCtrl.scala 159:32]
  wire [5:0] _T_4923 = _T_4767 - 6'h1; // @[FanCtrl.scala 203:56]
  wire [4:0] _GEN_49929 = 5'h3 == _T_4923[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_49930 = 5'h4 == _T_4923[4:0] ? w_vn_4 : _GEN_49929; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_49931 = 5'h5 == _T_4923[4:0] ? 5'h0 : _GEN_49930; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_49932 = 5'h6 == _T_4923[4:0] ? 5'h0 : _GEN_49931; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_49933 = 5'h7 == _T_4923[4:0] ? w_vn_7 : _GEN_49932; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_49934 = 5'h8 == _T_4923[4:0] ? w_vn_8 : _GEN_49933; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_49935 = 5'h9 == _T_4923[4:0] ? 5'h0 : _GEN_49934; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_49936 = 5'ha == _T_4923[4:0] ? 5'h0 : _GEN_49935; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_49937 = 5'hb == _T_4923[4:0] ? w_vn_11 : _GEN_49936; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_49938 = 5'hc == _T_4923[4:0] ? w_vn_12 : _GEN_49937; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_49939 = 5'hd == _T_4923[4:0] ? w_vn_13 : _GEN_49938; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_49940 = 5'he == _T_4923[4:0] ? 5'h0 : _GEN_49939; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_49941 = 5'hf == _T_4923[4:0] ? w_vn_15 : _GEN_49940; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_49942 = 5'h10 == _T_4923[4:0] ? w_vn_16 : _GEN_49941; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_49943 = 5'h11 == _T_4923[4:0] ? 5'h0 : _GEN_49942; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_49944 = 5'h12 == _T_4923[4:0] ? w_vn_18 : _GEN_49943; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_49945 = 5'h13 == _T_4923[4:0] ? 5'h0 : _GEN_49944; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_49946 = 5'h14 == _T_4923[4:0] ? 5'h0 : _GEN_49945; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_49947 = 5'h15 == _T_4923[4:0] ? 5'h0 : _GEN_49946; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_49948 = 5'h16 == _T_4923[4:0] ? 5'h0 : _GEN_49947; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_49949 = 5'h17 == _T_4923[4:0] ? w_vn_23 : _GEN_49948; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_49950 = 5'h18 == _T_4923[4:0] ? w_vn_24 : _GEN_49949; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_49951 = 5'h19 == _T_4923[4:0] ? 5'h0 : _GEN_49950; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_49952 = 5'h1a == _T_4923[4:0] ? 5'h0 : _GEN_49951; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_49953 = 5'h1b == _T_4923[4:0] ? 5'h0 : _GEN_49952; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_49954 = 5'h1c == _T_4923[4:0] ? 5'h0 : _GEN_49953; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_49955 = 5'h1d == _T_4923[4:0] ? 5'h0 : _GEN_49954; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_49956 = 5'h1e == _T_4923[4:0] ? 5'h0 : _GEN_49955; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_49957 = 5'h1f == _T_4923[4:0] ? 5'h0 : _GEN_49956; // @[FanCtrl.scala 203:{37,37}]
  wire  _T_4925 = _GEN_48661 != _GEN_49957; // @[FanCtrl.scala 203:37]
  wire  _T_4926 = _T_4798 & _T_4925; // @[FanCtrl.scala 202:65]
  wire  _T_4957 = _T_4788 & _T_4925; // @[FanCtrl.scala 208:71]
  wire  _T_4967 = _T_4957 & _T_4817; // @[FanCtrl.scala 209:70]
  wire  _T_5053 = _T_4926 & _T_4807; // @[FanCtrl.scala 239:64]
  wire  _T_5063 = _T_5053 & _T_4817; // @[FanCtrl.scala 240:62]
  wire [2:0] _GEN_51751 = _T_4967 ? 3'h3 : 3'h0; // @[FanCtrl.scala 253:70]
  wire [2:0] _GEN_51782 = _T_4849 ? 3'h4 : _GEN_51751; // @[FanCtrl.scala 247:70]
  wire [2:0] _GEN_51813 = _T_5063 ? 3'h5 : _GEN_51782; // @[FanCtrl.scala 241:64]
  wire [2:0] _GEN_51937 = r_valid_1 ? _GEN_51813 : 3'h0; // @[FanCtrl.scala 230:30]
  wire [5:0] _T_5140 = 3'h4 * 3'h6; // @[FanCtrl.scala 160:23]
  wire [5:0] _T_5142 = _T_5140 + 6'h1; // @[FanCtrl.scala 160:29]
  wire [5:0] _T_5146 = _T_5140 + 6'h2; // @[FanCtrl.scala 160:56]
  wire [4:0] _GEN_52136 = 5'h3 == _T_5142[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_52137 = 5'h4 == _T_5142[4:0] ? w_vn_4 : _GEN_52136; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_52138 = 5'h5 == _T_5142[4:0] ? 5'h0 : _GEN_52137; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_52139 = 5'h6 == _T_5142[4:0] ? 5'h0 : _GEN_52138; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_52140 = 5'h7 == _T_5142[4:0] ? w_vn_7 : _GEN_52139; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_52141 = 5'h8 == _T_5142[4:0] ? w_vn_8 : _GEN_52140; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_52142 = 5'h9 == _T_5142[4:0] ? 5'h0 : _GEN_52141; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_52143 = 5'ha == _T_5142[4:0] ? 5'h0 : _GEN_52142; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_52144 = 5'hb == _T_5142[4:0] ? w_vn_11 : _GEN_52143; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_52145 = 5'hc == _T_5142[4:0] ? w_vn_12 : _GEN_52144; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_52146 = 5'hd == _T_5142[4:0] ? w_vn_13 : _GEN_52145; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_52147 = 5'he == _T_5142[4:0] ? 5'h0 : _GEN_52146; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_52148 = 5'hf == _T_5142[4:0] ? w_vn_15 : _GEN_52147; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_52149 = 5'h10 == _T_5142[4:0] ? w_vn_16 : _GEN_52148; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_52150 = 5'h11 == _T_5142[4:0] ? 5'h0 : _GEN_52149; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_52151 = 5'h12 == _T_5142[4:0] ? w_vn_18 : _GEN_52150; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_52152 = 5'h13 == _T_5142[4:0] ? 5'h0 : _GEN_52151; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_52153 = 5'h14 == _T_5142[4:0] ? 5'h0 : _GEN_52152; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_52154 = 5'h15 == _T_5142[4:0] ? 5'h0 : _GEN_52153; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_52155 = 5'h16 == _T_5142[4:0] ? 5'h0 : _GEN_52154; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_52156 = 5'h17 == _T_5142[4:0] ? w_vn_23 : _GEN_52155; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_52157 = 5'h18 == _T_5142[4:0] ? w_vn_24 : _GEN_52156; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_52158 = 5'h19 == _T_5142[4:0] ? 5'h0 : _GEN_52157; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_52159 = 5'h1a == _T_5142[4:0] ? 5'h0 : _GEN_52158; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_52160 = 5'h1b == _T_5142[4:0] ? 5'h0 : _GEN_52159; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_52161 = 5'h1c == _T_5142[4:0] ? 5'h0 : _GEN_52160; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_52162 = 5'h1d == _T_5142[4:0] ? 5'h0 : _GEN_52161; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_52163 = 5'h1e == _T_5142[4:0] ? 5'h0 : _GEN_52162; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_52164 = 5'h1f == _T_5142[4:0] ? 5'h0 : _GEN_52163; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_52168 = 5'h3 == _T_5146[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_52169 = 5'h4 == _T_5146[4:0] ? w_vn_4 : _GEN_52168; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_52170 = 5'h5 == _T_5146[4:0] ? 5'h0 : _GEN_52169; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_52171 = 5'h6 == _T_5146[4:0] ? 5'h0 : _GEN_52170; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_52172 = 5'h7 == _T_5146[4:0] ? w_vn_7 : _GEN_52171; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_52173 = 5'h8 == _T_5146[4:0] ? w_vn_8 : _GEN_52172; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_52174 = 5'h9 == _T_5146[4:0] ? 5'h0 : _GEN_52173; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_52175 = 5'ha == _T_5146[4:0] ? 5'h0 : _GEN_52174; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_52176 = 5'hb == _T_5146[4:0] ? w_vn_11 : _GEN_52175; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_52177 = 5'hc == _T_5146[4:0] ? w_vn_12 : _GEN_52176; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_52178 = 5'hd == _T_5146[4:0] ? w_vn_13 : _GEN_52177; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_52179 = 5'he == _T_5146[4:0] ? 5'h0 : _GEN_52178; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_52180 = 5'hf == _T_5146[4:0] ? w_vn_15 : _GEN_52179; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_52181 = 5'h10 == _T_5146[4:0] ? w_vn_16 : _GEN_52180; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_52182 = 5'h11 == _T_5146[4:0] ? 5'h0 : _GEN_52181; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_52183 = 5'h12 == _T_5146[4:0] ? w_vn_18 : _GEN_52182; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_52184 = 5'h13 == _T_5146[4:0] ? 5'h0 : _GEN_52183; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_52185 = 5'h14 == _T_5146[4:0] ? 5'h0 : _GEN_52184; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_52186 = 5'h15 == _T_5146[4:0] ? 5'h0 : _GEN_52185; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_52187 = 5'h16 == _T_5146[4:0] ? 5'h0 : _GEN_52186; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_52188 = 5'h17 == _T_5146[4:0] ? w_vn_23 : _GEN_52187; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_52189 = 5'h18 == _T_5146[4:0] ? w_vn_24 : _GEN_52188; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_52190 = 5'h19 == _T_5146[4:0] ? 5'h0 : _GEN_52189; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_52191 = 5'h1a == _T_5146[4:0] ? 5'h0 : _GEN_52190; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_52192 = 5'h1b == _T_5146[4:0] ? 5'h0 : _GEN_52191; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_52193 = 5'h1c == _T_5146[4:0] ? 5'h0 : _GEN_52192; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_52194 = 5'h1d == _T_5146[4:0] ? 5'h0 : _GEN_52193; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_52195 = 5'h1e == _T_5146[4:0] ? 5'h0 : _GEN_52194; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_52196 = 5'h1f == _T_5146[4:0] ? 5'h0 : _GEN_52195; // @[FanCtrl.scala 160:{37,37}]
  wire  _T_5148 = _GEN_52164 == _GEN_52196; // @[FanCtrl.scala 160:37]
  wire [6:0] _T_5154 = {{1'd0}, _T_5140}; // @[FanCtrl.scala 166:30]
  wire [4:0] _GEN_52293 = 5'h3 == _T_5154[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_52294 = 5'h4 == _T_5154[4:0] ? w_vn_4 : _GEN_52293; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_52295 = 5'h5 == _T_5154[4:0] ? 5'h0 : _GEN_52294; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_52296 = 5'h6 == _T_5154[4:0] ? 5'h0 : _GEN_52295; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_52297 = 5'h7 == _T_5154[4:0] ? w_vn_7 : _GEN_52296; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_52298 = 5'h8 == _T_5154[4:0] ? w_vn_8 : _GEN_52297; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_52299 = 5'h9 == _T_5154[4:0] ? 5'h0 : _GEN_52298; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_52300 = 5'ha == _T_5154[4:0] ? 5'h0 : _GEN_52299; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_52301 = 5'hb == _T_5154[4:0] ? w_vn_11 : _GEN_52300; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_52302 = 5'hc == _T_5154[4:0] ? w_vn_12 : _GEN_52301; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_52303 = 5'hd == _T_5154[4:0] ? w_vn_13 : _GEN_52302; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_52304 = 5'he == _T_5154[4:0] ? 5'h0 : _GEN_52303; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_52305 = 5'hf == _T_5154[4:0] ? w_vn_15 : _GEN_52304; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_52306 = 5'h10 == _T_5154[4:0] ? w_vn_16 : _GEN_52305; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_52307 = 5'h11 == _T_5154[4:0] ? 5'h0 : _GEN_52306; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_52308 = 5'h12 == _T_5154[4:0] ? w_vn_18 : _GEN_52307; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_52309 = 5'h13 == _T_5154[4:0] ? 5'h0 : _GEN_52308; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_52310 = 5'h14 == _T_5154[4:0] ? 5'h0 : _GEN_52309; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_52311 = 5'h15 == _T_5154[4:0] ? 5'h0 : _GEN_52310; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_52312 = 5'h16 == _T_5154[4:0] ? 5'h0 : _GEN_52311; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_52313 = 5'h17 == _T_5154[4:0] ? w_vn_23 : _GEN_52312; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_52314 = 5'h18 == _T_5154[4:0] ? w_vn_24 : _GEN_52313; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_52315 = 5'h19 == _T_5154[4:0] ? 5'h0 : _GEN_52314; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_52316 = 5'h1a == _T_5154[4:0] ? 5'h0 : _GEN_52315; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_52317 = 5'h1b == _T_5154[4:0] ? 5'h0 : _GEN_52316; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_52318 = 5'h1c == _T_5154[4:0] ? 5'h0 : _GEN_52317; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_52319 = 5'h1d == _T_5154[4:0] ? 5'h0 : _GEN_52318; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_52320 = 5'h1e == _T_5154[4:0] ? 5'h0 : _GEN_52319; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_52321 = 5'h1f == _T_5154[4:0] ? 5'h0 : _GEN_52320; // @[FanCtrl.scala 166:{38,38}]
  wire  _T_5161 = _GEN_52321 == _GEN_52164; // @[FanCtrl.scala 166:38]
  wire [5:0] _T_5168 = _T_5140 + 6'h3; // @[FanCtrl.scala 167:55]
  wire [4:0] _GEN_52389 = 5'h3 == _T_5168[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_52390 = 5'h4 == _T_5168[4:0] ? w_vn_4 : _GEN_52389; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_52391 = 5'h5 == _T_5168[4:0] ? 5'h0 : _GEN_52390; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_52392 = 5'h6 == _T_5168[4:0] ? 5'h0 : _GEN_52391; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_52393 = 5'h7 == _T_5168[4:0] ? w_vn_7 : _GEN_52392; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_52394 = 5'h8 == _T_5168[4:0] ? w_vn_8 : _GEN_52393; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_52395 = 5'h9 == _T_5168[4:0] ? 5'h0 : _GEN_52394; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_52396 = 5'ha == _T_5168[4:0] ? 5'h0 : _GEN_52395; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_52397 = 5'hb == _T_5168[4:0] ? w_vn_11 : _GEN_52396; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_52398 = 5'hc == _T_5168[4:0] ? w_vn_12 : _GEN_52397; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_52399 = 5'hd == _T_5168[4:0] ? w_vn_13 : _GEN_52398; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_52400 = 5'he == _T_5168[4:0] ? 5'h0 : _GEN_52399; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_52401 = 5'hf == _T_5168[4:0] ? w_vn_15 : _GEN_52400; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_52402 = 5'h10 == _T_5168[4:0] ? w_vn_16 : _GEN_52401; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_52403 = 5'h11 == _T_5168[4:0] ? 5'h0 : _GEN_52402; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_52404 = 5'h12 == _T_5168[4:0] ? w_vn_18 : _GEN_52403; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_52405 = 5'h13 == _T_5168[4:0] ? 5'h0 : _GEN_52404; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_52406 = 5'h14 == _T_5168[4:0] ? 5'h0 : _GEN_52405; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_52407 = 5'h15 == _T_5168[4:0] ? 5'h0 : _GEN_52406; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_52408 = 5'h16 == _T_5168[4:0] ? 5'h0 : _GEN_52407; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_52409 = 5'h17 == _T_5168[4:0] ? w_vn_23 : _GEN_52408; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_52410 = 5'h18 == _T_5168[4:0] ? w_vn_24 : _GEN_52409; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_52411 = 5'h19 == _T_5168[4:0] ? 5'h0 : _GEN_52410; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_52412 = 5'h1a == _T_5168[4:0] ? 5'h0 : _GEN_52411; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_52413 = 5'h1b == _T_5168[4:0] ? 5'h0 : _GEN_52412; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_52414 = 5'h1c == _T_5168[4:0] ? 5'h0 : _GEN_52413; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_52415 = 5'h1d == _T_5168[4:0] ? 5'h0 : _GEN_52414; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_52416 = 5'h1e == _T_5168[4:0] ? 5'h0 : _GEN_52415; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_52417 = 5'h1f == _T_5168[4:0] ? 5'h0 : _GEN_52416; // @[FanCtrl.scala 167:{36,36}]
  wire  _T_5170 = _GEN_52196 == _GEN_52417; // @[FanCtrl.scala 167:36]
  wire  _T_5171 = _GEN_52321 == _GEN_52164 & _T_5170; // @[FanCtrl.scala 166:65]
  wire [5:0] _T_5174 = _T_5140 + 6'h4; // @[FanCtrl.scala 168:29]
  wire [4:0] _GEN_52421 = 5'h3 == _T_5174[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_52422 = 5'h4 == _T_5174[4:0] ? w_vn_4 : _GEN_52421; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_52423 = 5'h5 == _T_5174[4:0] ? 5'h0 : _GEN_52422; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_52424 = 5'h6 == _T_5174[4:0] ? 5'h0 : _GEN_52423; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_52425 = 5'h7 == _T_5174[4:0] ? w_vn_7 : _GEN_52424; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_52426 = 5'h8 == _T_5174[4:0] ? w_vn_8 : _GEN_52425; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_52427 = 5'h9 == _T_5174[4:0] ? 5'h0 : _GEN_52426; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_52428 = 5'ha == _T_5174[4:0] ? 5'h0 : _GEN_52427; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_52429 = 5'hb == _T_5174[4:0] ? w_vn_11 : _GEN_52428; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_52430 = 5'hc == _T_5174[4:0] ? w_vn_12 : _GEN_52429; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_52431 = 5'hd == _T_5174[4:0] ? w_vn_13 : _GEN_52430; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_52432 = 5'he == _T_5174[4:0] ? 5'h0 : _GEN_52431; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_52433 = 5'hf == _T_5174[4:0] ? w_vn_15 : _GEN_52432; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_52434 = 5'h10 == _T_5174[4:0] ? w_vn_16 : _GEN_52433; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_52435 = 5'h11 == _T_5174[4:0] ? 5'h0 : _GEN_52434; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_52436 = 5'h12 == _T_5174[4:0] ? w_vn_18 : _GEN_52435; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_52437 = 5'h13 == _T_5174[4:0] ? 5'h0 : _GEN_52436; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_52438 = 5'h14 == _T_5174[4:0] ? 5'h0 : _GEN_52437; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_52439 = 5'h15 == _T_5174[4:0] ? 5'h0 : _GEN_52438; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_52440 = 5'h16 == _T_5174[4:0] ? 5'h0 : _GEN_52439; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_52441 = 5'h17 == _T_5174[4:0] ? w_vn_23 : _GEN_52440; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_52442 = 5'h18 == _T_5174[4:0] ? w_vn_24 : _GEN_52441; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_52443 = 5'h19 == _T_5174[4:0] ? 5'h0 : _GEN_52442; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_52444 = 5'h1a == _T_5174[4:0] ? 5'h0 : _GEN_52443; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_52445 = 5'h1b == _T_5174[4:0] ? 5'h0 : _GEN_52444; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_52446 = 5'h1c == _T_5174[4:0] ? 5'h0 : _GEN_52445; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_52447 = 5'h1d == _T_5174[4:0] ? 5'h0 : _GEN_52446; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_52448 = 5'h1e == _T_5174[4:0] ? 5'h0 : _GEN_52447; // @[FanCtrl.scala 168:{37,37}]
  wire [4:0] _GEN_52449 = 5'h1f == _T_5174[4:0] ? 5'h0 : _GEN_52448; // @[FanCtrl.scala 168:{37,37}]
  wire  _T_5180 = _GEN_52449 != _GEN_52417; // @[FanCtrl.scala 168:37]
  wire  _T_5190 = _GEN_52164 != _GEN_52196; // @[FanCtrl.scala 169:37]
  wire  _T_5212 = _T_5170 & _T_5180; // @[FanCtrl.scala 173:71]
  wire  _T_5222 = _T_5212 & _T_5190; // @[FanCtrl.scala 174:71]
  wire  _GEN_53167 = r_valid_1 & _T_5148; // @[FanCtrl.scala 159:32]
  wire [5:0] _T_5296 = _T_5140 - 6'h1; // @[FanCtrl.scala 203:56]
  wire [4:0] _GEN_53589 = 5'h3 == _T_5296[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_53590 = 5'h4 == _T_5296[4:0] ? w_vn_4 : _GEN_53589; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_53591 = 5'h5 == _T_5296[4:0] ? 5'h0 : _GEN_53590; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_53592 = 5'h6 == _T_5296[4:0] ? 5'h0 : _GEN_53591; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_53593 = 5'h7 == _T_5296[4:0] ? w_vn_7 : _GEN_53592; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_53594 = 5'h8 == _T_5296[4:0] ? w_vn_8 : _GEN_53593; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_53595 = 5'h9 == _T_5296[4:0] ? 5'h0 : _GEN_53594; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_53596 = 5'ha == _T_5296[4:0] ? 5'h0 : _GEN_53595; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_53597 = 5'hb == _T_5296[4:0] ? w_vn_11 : _GEN_53596; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_53598 = 5'hc == _T_5296[4:0] ? w_vn_12 : _GEN_53597; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_53599 = 5'hd == _T_5296[4:0] ? w_vn_13 : _GEN_53598; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_53600 = 5'he == _T_5296[4:0] ? 5'h0 : _GEN_53599; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_53601 = 5'hf == _T_5296[4:0] ? w_vn_15 : _GEN_53600; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_53602 = 5'h10 == _T_5296[4:0] ? w_vn_16 : _GEN_53601; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_53603 = 5'h11 == _T_5296[4:0] ? 5'h0 : _GEN_53602; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_53604 = 5'h12 == _T_5296[4:0] ? w_vn_18 : _GEN_53603; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_53605 = 5'h13 == _T_5296[4:0] ? 5'h0 : _GEN_53604; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_53606 = 5'h14 == _T_5296[4:0] ? 5'h0 : _GEN_53605; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_53607 = 5'h15 == _T_5296[4:0] ? 5'h0 : _GEN_53606; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_53608 = 5'h16 == _T_5296[4:0] ? 5'h0 : _GEN_53607; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_53609 = 5'h17 == _T_5296[4:0] ? w_vn_23 : _GEN_53608; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_53610 = 5'h18 == _T_5296[4:0] ? w_vn_24 : _GEN_53609; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_53611 = 5'h19 == _T_5296[4:0] ? 5'h0 : _GEN_53610; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_53612 = 5'h1a == _T_5296[4:0] ? 5'h0 : _GEN_53611; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_53613 = 5'h1b == _T_5296[4:0] ? 5'h0 : _GEN_53612; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_53614 = 5'h1c == _T_5296[4:0] ? 5'h0 : _GEN_53613; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_53615 = 5'h1d == _T_5296[4:0] ? 5'h0 : _GEN_53614; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_53616 = 5'h1e == _T_5296[4:0] ? 5'h0 : _GEN_53615; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_53617 = 5'h1f == _T_5296[4:0] ? 5'h0 : _GEN_53616; // @[FanCtrl.scala 203:{37,37}]
  wire  _T_5298 = _GEN_52321 != _GEN_53617; // @[FanCtrl.scala 203:37]
  wire  _T_5299 = _T_5171 & _T_5298; // @[FanCtrl.scala 202:65]
  wire  _T_5330 = _T_5161 & _T_5298; // @[FanCtrl.scala 208:71]
  wire  _T_5340 = _T_5330 & _T_5190; // @[FanCtrl.scala 209:70]
  wire  _T_5426 = _T_5299 & _T_5180; // @[FanCtrl.scala 239:64]
  wire  _T_5436 = _T_5426 & _T_5190; // @[FanCtrl.scala 240:62]
  wire [2:0] _GEN_55412 = _T_5340 ? 3'h3 : 3'h0; // @[FanCtrl.scala 253:70]
  wire [2:0] _GEN_55443 = _T_5222 ? 3'h4 : _GEN_55412; // @[FanCtrl.scala 247:70]
  wire [2:0] _GEN_55474 = _T_5436 ? 3'h5 : _GEN_55443; // @[FanCtrl.scala 241:64]
  wire [2:0] _GEN_55598 = r_valid_1 ? _GEN_55474 : 3'h0; // @[FanCtrl.scala 230:30]
  wire [5:0] _T_5513 = 3'h4 * 3'h7; // @[FanCtrl.scala 160:23]
  wire [5:0] _T_5515 = _T_5513 + 6'h1; // @[FanCtrl.scala 160:29]
  wire [5:0] _T_5519 = _T_5513 + 6'h2; // @[FanCtrl.scala 160:56]
  wire [4:0] _GEN_55796 = 5'h3 == _T_5515[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_55797 = 5'h4 == _T_5515[4:0] ? w_vn_4 : _GEN_55796; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_55798 = 5'h5 == _T_5515[4:0] ? 5'h0 : _GEN_55797; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_55799 = 5'h6 == _T_5515[4:0] ? 5'h0 : _GEN_55798; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_55800 = 5'h7 == _T_5515[4:0] ? w_vn_7 : _GEN_55799; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_55801 = 5'h8 == _T_5515[4:0] ? w_vn_8 : _GEN_55800; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_55802 = 5'h9 == _T_5515[4:0] ? 5'h0 : _GEN_55801; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_55803 = 5'ha == _T_5515[4:0] ? 5'h0 : _GEN_55802; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_55804 = 5'hb == _T_5515[4:0] ? w_vn_11 : _GEN_55803; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_55805 = 5'hc == _T_5515[4:0] ? w_vn_12 : _GEN_55804; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_55806 = 5'hd == _T_5515[4:0] ? w_vn_13 : _GEN_55805; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_55807 = 5'he == _T_5515[4:0] ? 5'h0 : _GEN_55806; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_55808 = 5'hf == _T_5515[4:0] ? w_vn_15 : _GEN_55807; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_55809 = 5'h10 == _T_5515[4:0] ? w_vn_16 : _GEN_55808; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_55810 = 5'h11 == _T_5515[4:0] ? 5'h0 : _GEN_55809; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_55811 = 5'h12 == _T_5515[4:0] ? w_vn_18 : _GEN_55810; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_55812 = 5'h13 == _T_5515[4:0] ? 5'h0 : _GEN_55811; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_55813 = 5'h14 == _T_5515[4:0] ? 5'h0 : _GEN_55812; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_55814 = 5'h15 == _T_5515[4:0] ? 5'h0 : _GEN_55813; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_55815 = 5'h16 == _T_5515[4:0] ? 5'h0 : _GEN_55814; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_55816 = 5'h17 == _T_5515[4:0] ? w_vn_23 : _GEN_55815; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_55817 = 5'h18 == _T_5515[4:0] ? w_vn_24 : _GEN_55816; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_55818 = 5'h19 == _T_5515[4:0] ? 5'h0 : _GEN_55817; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_55819 = 5'h1a == _T_5515[4:0] ? 5'h0 : _GEN_55818; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_55820 = 5'h1b == _T_5515[4:0] ? 5'h0 : _GEN_55819; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_55821 = 5'h1c == _T_5515[4:0] ? 5'h0 : _GEN_55820; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_55822 = 5'h1d == _T_5515[4:0] ? 5'h0 : _GEN_55821; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_55823 = 5'h1e == _T_5515[4:0] ? 5'h0 : _GEN_55822; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_55824 = 5'h1f == _T_5515[4:0] ? 5'h0 : _GEN_55823; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_55828 = 5'h3 == _T_5519[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_55829 = 5'h4 == _T_5519[4:0] ? w_vn_4 : _GEN_55828; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_55830 = 5'h5 == _T_5519[4:0] ? 5'h0 : _GEN_55829; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_55831 = 5'h6 == _T_5519[4:0] ? 5'h0 : _GEN_55830; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_55832 = 5'h7 == _T_5519[4:0] ? w_vn_7 : _GEN_55831; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_55833 = 5'h8 == _T_5519[4:0] ? w_vn_8 : _GEN_55832; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_55834 = 5'h9 == _T_5519[4:0] ? 5'h0 : _GEN_55833; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_55835 = 5'ha == _T_5519[4:0] ? 5'h0 : _GEN_55834; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_55836 = 5'hb == _T_5519[4:0] ? w_vn_11 : _GEN_55835; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_55837 = 5'hc == _T_5519[4:0] ? w_vn_12 : _GEN_55836; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_55838 = 5'hd == _T_5519[4:0] ? w_vn_13 : _GEN_55837; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_55839 = 5'he == _T_5519[4:0] ? 5'h0 : _GEN_55838; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_55840 = 5'hf == _T_5519[4:0] ? w_vn_15 : _GEN_55839; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_55841 = 5'h10 == _T_5519[4:0] ? w_vn_16 : _GEN_55840; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_55842 = 5'h11 == _T_5519[4:0] ? 5'h0 : _GEN_55841; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_55843 = 5'h12 == _T_5519[4:0] ? w_vn_18 : _GEN_55842; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_55844 = 5'h13 == _T_5519[4:0] ? 5'h0 : _GEN_55843; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_55845 = 5'h14 == _T_5519[4:0] ? 5'h0 : _GEN_55844; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_55846 = 5'h15 == _T_5519[4:0] ? 5'h0 : _GEN_55845; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_55847 = 5'h16 == _T_5519[4:0] ? 5'h0 : _GEN_55846; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_55848 = 5'h17 == _T_5519[4:0] ? w_vn_23 : _GEN_55847; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_55849 = 5'h18 == _T_5519[4:0] ? w_vn_24 : _GEN_55848; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_55850 = 5'h19 == _T_5519[4:0] ? 5'h0 : _GEN_55849; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_55851 = 5'h1a == _T_5519[4:0] ? 5'h0 : _GEN_55850; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_55852 = 5'h1b == _T_5519[4:0] ? 5'h0 : _GEN_55851; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_55853 = 5'h1c == _T_5519[4:0] ? 5'h0 : _GEN_55852; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_55854 = 5'h1d == _T_5519[4:0] ? 5'h0 : _GEN_55853; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_55855 = 5'h1e == _T_5519[4:0] ? 5'h0 : _GEN_55854; // @[FanCtrl.scala 160:{37,37}]
  wire [4:0] _GEN_55856 = 5'h1f == _T_5519[4:0] ? 5'h0 : _GEN_55855; // @[FanCtrl.scala 160:{37,37}]
  wire  _T_5521 = _GEN_55824 == _GEN_55856; // @[FanCtrl.scala 160:37]
  wire [6:0] _T_5527 = {{1'd0}, _T_5513}; // @[FanCtrl.scala 166:30]
  wire [4:0] _GEN_55953 = 5'h3 == _T_5527[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_55954 = 5'h4 == _T_5527[4:0] ? w_vn_4 : _GEN_55953; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_55955 = 5'h5 == _T_5527[4:0] ? 5'h0 : _GEN_55954; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_55956 = 5'h6 == _T_5527[4:0] ? 5'h0 : _GEN_55955; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_55957 = 5'h7 == _T_5527[4:0] ? w_vn_7 : _GEN_55956; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_55958 = 5'h8 == _T_5527[4:0] ? w_vn_8 : _GEN_55957; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_55959 = 5'h9 == _T_5527[4:0] ? 5'h0 : _GEN_55958; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_55960 = 5'ha == _T_5527[4:0] ? 5'h0 : _GEN_55959; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_55961 = 5'hb == _T_5527[4:0] ? w_vn_11 : _GEN_55960; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_55962 = 5'hc == _T_5527[4:0] ? w_vn_12 : _GEN_55961; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_55963 = 5'hd == _T_5527[4:0] ? w_vn_13 : _GEN_55962; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_55964 = 5'he == _T_5527[4:0] ? 5'h0 : _GEN_55963; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_55965 = 5'hf == _T_5527[4:0] ? w_vn_15 : _GEN_55964; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_55966 = 5'h10 == _T_5527[4:0] ? w_vn_16 : _GEN_55965; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_55967 = 5'h11 == _T_5527[4:0] ? 5'h0 : _GEN_55966; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_55968 = 5'h12 == _T_5527[4:0] ? w_vn_18 : _GEN_55967; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_55969 = 5'h13 == _T_5527[4:0] ? 5'h0 : _GEN_55968; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_55970 = 5'h14 == _T_5527[4:0] ? 5'h0 : _GEN_55969; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_55971 = 5'h15 == _T_5527[4:0] ? 5'h0 : _GEN_55970; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_55972 = 5'h16 == _T_5527[4:0] ? 5'h0 : _GEN_55971; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_55973 = 5'h17 == _T_5527[4:0] ? w_vn_23 : _GEN_55972; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_55974 = 5'h18 == _T_5527[4:0] ? w_vn_24 : _GEN_55973; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_55975 = 5'h19 == _T_5527[4:0] ? 5'h0 : _GEN_55974; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_55976 = 5'h1a == _T_5527[4:0] ? 5'h0 : _GEN_55975; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_55977 = 5'h1b == _T_5527[4:0] ? 5'h0 : _GEN_55976; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_55978 = 5'h1c == _T_5527[4:0] ? 5'h0 : _GEN_55977; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_55979 = 5'h1d == _T_5527[4:0] ? 5'h0 : _GEN_55978; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_55980 = 5'h1e == _T_5527[4:0] ? 5'h0 : _GEN_55979; // @[FanCtrl.scala 166:{38,38}]
  wire [4:0] _GEN_55981 = 5'h1f == _T_5527[4:0] ? 5'h0 : _GEN_55980; // @[FanCtrl.scala 166:{38,38}]
  wire  _T_5534 = _GEN_55981 == _GEN_55824; // @[FanCtrl.scala 166:38]
  wire [5:0] _T_5541 = _T_5513 + 6'h3; // @[FanCtrl.scala 167:55]
  wire [4:0] _GEN_56049 = 5'h3 == _T_5541[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_56050 = 5'h4 == _T_5541[4:0] ? w_vn_4 : _GEN_56049; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_56051 = 5'h5 == _T_5541[4:0] ? 5'h0 : _GEN_56050; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_56052 = 5'h6 == _T_5541[4:0] ? 5'h0 : _GEN_56051; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_56053 = 5'h7 == _T_5541[4:0] ? w_vn_7 : _GEN_56052; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_56054 = 5'h8 == _T_5541[4:0] ? w_vn_8 : _GEN_56053; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_56055 = 5'h9 == _T_5541[4:0] ? 5'h0 : _GEN_56054; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_56056 = 5'ha == _T_5541[4:0] ? 5'h0 : _GEN_56055; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_56057 = 5'hb == _T_5541[4:0] ? w_vn_11 : _GEN_56056; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_56058 = 5'hc == _T_5541[4:0] ? w_vn_12 : _GEN_56057; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_56059 = 5'hd == _T_5541[4:0] ? w_vn_13 : _GEN_56058; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_56060 = 5'he == _T_5541[4:0] ? 5'h0 : _GEN_56059; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_56061 = 5'hf == _T_5541[4:0] ? w_vn_15 : _GEN_56060; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_56062 = 5'h10 == _T_5541[4:0] ? w_vn_16 : _GEN_56061; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_56063 = 5'h11 == _T_5541[4:0] ? 5'h0 : _GEN_56062; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_56064 = 5'h12 == _T_5541[4:0] ? w_vn_18 : _GEN_56063; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_56065 = 5'h13 == _T_5541[4:0] ? 5'h0 : _GEN_56064; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_56066 = 5'h14 == _T_5541[4:0] ? 5'h0 : _GEN_56065; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_56067 = 5'h15 == _T_5541[4:0] ? 5'h0 : _GEN_56066; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_56068 = 5'h16 == _T_5541[4:0] ? 5'h0 : _GEN_56067; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_56069 = 5'h17 == _T_5541[4:0] ? w_vn_23 : _GEN_56068; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_56070 = 5'h18 == _T_5541[4:0] ? w_vn_24 : _GEN_56069; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_56071 = 5'h19 == _T_5541[4:0] ? 5'h0 : _GEN_56070; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_56072 = 5'h1a == _T_5541[4:0] ? 5'h0 : _GEN_56071; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_56073 = 5'h1b == _T_5541[4:0] ? 5'h0 : _GEN_56072; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_56074 = 5'h1c == _T_5541[4:0] ? 5'h0 : _GEN_56073; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_56075 = 5'h1d == _T_5541[4:0] ? 5'h0 : _GEN_56074; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_56076 = 5'h1e == _T_5541[4:0] ? 5'h0 : _GEN_56075; // @[FanCtrl.scala 167:{36,36}]
  wire [4:0] _GEN_56077 = 5'h1f == _T_5541[4:0] ? 5'h0 : _GEN_56076; // @[FanCtrl.scala 167:{36,36}]
  wire  _T_5543 = _GEN_55856 == _GEN_56077; // @[FanCtrl.scala 167:36]
  wire  _T_5544 = _GEN_55981 == _GEN_55824 & _T_5543; // @[FanCtrl.scala 166:65]
  wire  _T_5563 = _GEN_55824 != _GEN_55856; // @[FanCtrl.scala 169:37]
  wire  _GEN_56828 = r_valid_1 & _T_5521; // @[FanCtrl.scala 159:32]
  wire [5:0] _T_5669 = _T_5513 - 6'h1; // @[FanCtrl.scala 203:56]
  wire [4:0] _GEN_57249 = 5'h3 == _T_5669[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_57250 = 5'h4 == _T_5669[4:0] ? w_vn_4 : _GEN_57249; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_57251 = 5'h5 == _T_5669[4:0] ? 5'h0 : _GEN_57250; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_57252 = 5'h6 == _T_5669[4:0] ? 5'h0 : _GEN_57251; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_57253 = 5'h7 == _T_5669[4:0] ? w_vn_7 : _GEN_57252; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_57254 = 5'h8 == _T_5669[4:0] ? w_vn_8 : _GEN_57253; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_57255 = 5'h9 == _T_5669[4:0] ? 5'h0 : _GEN_57254; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_57256 = 5'ha == _T_5669[4:0] ? 5'h0 : _GEN_57255; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_57257 = 5'hb == _T_5669[4:0] ? w_vn_11 : _GEN_57256; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_57258 = 5'hc == _T_5669[4:0] ? w_vn_12 : _GEN_57257; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_57259 = 5'hd == _T_5669[4:0] ? w_vn_13 : _GEN_57258; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_57260 = 5'he == _T_5669[4:0] ? 5'h0 : _GEN_57259; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_57261 = 5'hf == _T_5669[4:0] ? w_vn_15 : _GEN_57260; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_57262 = 5'h10 == _T_5669[4:0] ? w_vn_16 : _GEN_57261; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_57263 = 5'h11 == _T_5669[4:0] ? 5'h0 : _GEN_57262; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_57264 = 5'h12 == _T_5669[4:0] ? w_vn_18 : _GEN_57263; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_57265 = 5'h13 == _T_5669[4:0] ? 5'h0 : _GEN_57264; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_57266 = 5'h14 == _T_5669[4:0] ? 5'h0 : _GEN_57265; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_57267 = 5'h15 == _T_5669[4:0] ? 5'h0 : _GEN_57266; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_57268 = 5'h16 == _T_5669[4:0] ? 5'h0 : _GEN_57267; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_57269 = 5'h17 == _T_5669[4:0] ? w_vn_23 : _GEN_57268; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_57270 = 5'h18 == _T_5669[4:0] ? w_vn_24 : _GEN_57269; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_57271 = 5'h19 == _T_5669[4:0] ? 5'h0 : _GEN_57270; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_57272 = 5'h1a == _T_5669[4:0] ? 5'h0 : _GEN_57271; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_57273 = 5'h1b == _T_5669[4:0] ? 5'h0 : _GEN_57272; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_57274 = 5'h1c == _T_5669[4:0] ? 5'h0 : _GEN_57273; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_57275 = 5'h1d == _T_5669[4:0] ? 5'h0 : _GEN_57274; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_57276 = 5'h1e == _T_5669[4:0] ? 5'h0 : _GEN_57275; // @[FanCtrl.scala 203:{37,37}]
  wire [4:0] _GEN_57277 = 5'h1f == _T_5669[4:0] ? 5'h0 : _GEN_57276; // @[FanCtrl.scala 203:{37,37}]
  wire  _T_5671 = _GEN_55981 != _GEN_57277; // @[FanCtrl.scala 203:37]
  wire  _T_5672 = _T_5544 & _T_5671; // @[FanCtrl.scala 202:65]
  wire  _T_5682 = _T_5672 & _T_5563; // @[FanCtrl.scala 203:65]
  wire  _T_5703 = _T_5534 & _T_5671; // @[FanCtrl.scala 208:71]
  wire  _T_5713 = _T_5703 & _T_5563; // @[FanCtrl.scala 209:70]
  wire  _T_5734 = _T_5543 & _T_5563; // @[FanCtrl.scala 214:71]
  wire [2:0] _GEN_57809 = _T_5734 ? 3'h4 : 3'h0; // @[FanCtrl.scala 215:72]
  wire [2:0] _GEN_57840 = _T_5713 ? 3'h3 : _GEN_57809; // @[FanCtrl.scala 210:71]
  wire [2:0] _GEN_57871 = _T_5682 ? 3'h5 : _GEN_57840; // @[FanCtrl.scala 204:65]
  wire [2:0] _GEN_57995 = r_valid_1 ? _GEN_57871 : 3'h0; // @[FanCtrl.scala 194:35]
  wire [4:0] _T_5888 = 4'h8 * 1'h0; // @[FanCtrl.scala 276:23]
  wire [4:0] _T_5890 = _T_5888 + 5'h3; // @[FanCtrl.scala 276:29]
  wire [4:0] _T_5893 = _T_5888 + 5'h4; // @[FanCtrl.scala 276:56]
  wire [4:0] _GEN_59476 = 5'h3 == _T_5890 ? w_vn_3 : 5'h0; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_59477 = 5'h4 == _T_5890 ? w_vn_4 : _GEN_59476; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_59478 = 5'h5 == _T_5890 ? 5'h0 : _GEN_59477; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_59479 = 5'h6 == _T_5890 ? 5'h0 : _GEN_59478; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_59480 = 5'h7 == _T_5890 ? w_vn_7 : _GEN_59479; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_59481 = 5'h8 == _T_5890 ? w_vn_8 : _GEN_59480; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_59482 = 5'h9 == _T_5890 ? 5'h0 : _GEN_59481; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_59483 = 5'ha == _T_5890 ? 5'h0 : _GEN_59482; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_59484 = 5'hb == _T_5890 ? w_vn_11 : _GEN_59483; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_59485 = 5'hc == _T_5890 ? w_vn_12 : _GEN_59484; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_59486 = 5'hd == _T_5890 ? w_vn_13 : _GEN_59485; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_59487 = 5'he == _T_5890 ? 5'h0 : _GEN_59486; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_59488 = 5'hf == _T_5890 ? w_vn_15 : _GEN_59487; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_59489 = 5'h10 == _T_5890 ? w_vn_16 : _GEN_59488; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_59490 = 5'h11 == _T_5890 ? 5'h0 : _GEN_59489; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_59491 = 5'h12 == _T_5890 ? w_vn_18 : _GEN_59490; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_59492 = 5'h13 == _T_5890 ? 5'h0 : _GEN_59491; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_59493 = 5'h14 == _T_5890 ? 5'h0 : _GEN_59492; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_59494 = 5'h15 == _T_5890 ? 5'h0 : _GEN_59493; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_59495 = 5'h16 == _T_5890 ? 5'h0 : _GEN_59494; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_59496 = 5'h17 == _T_5890 ? w_vn_23 : _GEN_59495; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_59497 = 5'h18 == _T_5890 ? w_vn_24 : _GEN_59496; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_59498 = 5'h19 == _T_5890 ? 5'h0 : _GEN_59497; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_59499 = 5'h1a == _T_5890 ? 5'h0 : _GEN_59498; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_59500 = 5'h1b == _T_5890 ? 5'h0 : _GEN_59499; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_59501 = 5'h1c == _T_5890 ? 5'h0 : _GEN_59500; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_59502 = 5'h1d == _T_5890 ? 5'h0 : _GEN_59501; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_59503 = 5'h1e == _T_5890 ? 5'h0 : _GEN_59502; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_59504 = 5'h1f == _T_5890 ? 5'h0 : _GEN_59503; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_59508 = 5'h3 == _T_5893 ? w_vn_3 : 5'h0; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_59509 = 5'h4 == _T_5893 ? w_vn_4 : _GEN_59508; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_59510 = 5'h5 == _T_5893 ? 5'h0 : _GEN_59509; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_59511 = 5'h6 == _T_5893 ? 5'h0 : _GEN_59510; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_59512 = 5'h7 == _T_5893 ? w_vn_7 : _GEN_59511; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_59513 = 5'h8 == _T_5893 ? w_vn_8 : _GEN_59512; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_59514 = 5'h9 == _T_5893 ? 5'h0 : _GEN_59513; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_59515 = 5'ha == _T_5893 ? 5'h0 : _GEN_59514; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_59516 = 5'hb == _T_5893 ? w_vn_11 : _GEN_59515; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_59517 = 5'hc == _T_5893 ? w_vn_12 : _GEN_59516; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_59518 = 5'hd == _T_5893 ? w_vn_13 : _GEN_59517; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_59519 = 5'he == _T_5893 ? 5'h0 : _GEN_59518; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_59520 = 5'hf == _T_5893 ? w_vn_15 : _GEN_59519; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_59521 = 5'h10 == _T_5893 ? w_vn_16 : _GEN_59520; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_59522 = 5'h11 == _T_5893 ? 5'h0 : _GEN_59521; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_59523 = 5'h12 == _T_5893 ? w_vn_18 : _GEN_59522; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_59524 = 5'h13 == _T_5893 ? 5'h0 : _GEN_59523; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_59525 = 5'h14 == _T_5893 ? 5'h0 : _GEN_59524; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_59526 = 5'h15 == _T_5893 ? 5'h0 : _GEN_59525; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_59527 = 5'h16 == _T_5893 ? 5'h0 : _GEN_59526; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_59528 = 5'h17 == _T_5893 ? w_vn_23 : _GEN_59527; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_59529 = 5'h18 == _T_5893 ? w_vn_24 : _GEN_59528; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_59530 = 5'h19 == _T_5893 ? 5'h0 : _GEN_59529; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_59531 = 5'h1a == _T_5893 ? 5'h0 : _GEN_59530; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_59532 = 5'h1b == _T_5893 ? 5'h0 : _GEN_59531; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_59533 = 5'h1c == _T_5893 ? 5'h0 : _GEN_59532; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_59534 = 5'h1d == _T_5893 ? 5'h0 : _GEN_59533; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_59535 = 5'h1e == _T_5893 ? 5'h0 : _GEN_59534; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_59536 = 5'h1f == _T_5893 ? 5'h0 : _GEN_59535; // @[FanCtrl.scala 276:{37,37}]
  wire  _T_5894 = _GEN_59504 == _GEN_59536; // @[FanCtrl.scala 276:37]
  wire [4:0] _T_5901 = _T_5888 + 5'h1; // @[FanCtrl.scala 282:30]
  wire [4:0] _T_5904 = _T_5888 + 5'h2; // @[FanCtrl.scala 282:56]
  wire [4:0] _GEN_59633 = 5'h3 == _T_5901 ? w_vn_3 : 5'h0; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_59634 = 5'h4 == _T_5901 ? w_vn_4 : _GEN_59633; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_59635 = 5'h5 == _T_5901 ? 5'h0 : _GEN_59634; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_59636 = 5'h6 == _T_5901 ? 5'h0 : _GEN_59635; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_59637 = 5'h7 == _T_5901 ? w_vn_7 : _GEN_59636; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_59638 = 5'h8 == _T_5901 ? w_vn_8 : _GEN_59637; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_59639 = 5'h9 == _T_5901 ? 5'h0 : _GEN_59638; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_59640 = 5'ha == _T_5901 ? 5'h0 : _GEN_59639; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_59641 = 5'hb == _T_5901 ? w_vn_11 : _GEN_59640; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_59642 = 5'hc == _T_5901 ? w_vn_12 : _GEN_59641; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_59643 = 5'hd == _T_5901 ? w_vn_13 : _GEN_59642; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_59644 = 5'he == _T_5901 ? 5'h0 : _GEN_59643; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_59645 = 5'hf == _T_5901 ? w_vn_15 : _GEN_59644; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_59646 = 5'h10 == _T_5901 ? w_vn_16 : _GEN_59645; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_59647 = 5'h11 == _T_5901 ? 5'h0 : _GEN_59646; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_59648 = 5'h12 == _T_5901 ? w_vn_18 : _GEN_59647; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_59649 = 5'h13 == _T_5901 ? 5'h0 : _GEN_59648; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_59650 = 5'h14 == _T_5901 ? 5'h0 : _GEN_59649; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_59651 = 5'h15 == _T_5901 ? 5'h0 : _GEN_59650; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_59652 = 5'h16 == _T_5901 ? 5'h0 : _GEN_59651; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_59653 = 5'h17 == _T_5901 ? w_vn_23 : _GEN_59652; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_59654 = 5'h18 == _T_5901 ? w_vn_24 : _GEN_59653; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_59655 = 5'h19 == _T_5901 ? 5'h0 : _GEN_59654; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_59656 = 5'h1a == _T_5901 ? 5'h0 : _GEN_59655; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_59657 = 5'h1b == _T_5901 ? 5'h0 : _GEN_59656; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_59658 = 5'h1c == _T_5901 ? 5'h0 : _GEN_59657; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_59659 = 5'h1d == _T_5901 ? 5'h0 : _GEN_59658; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_59660 = 5'h1e == _T_5901 ? 5'h0 : _GEN_59659; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_59661 = 5'h1f == _T_5901 ? 5'h0 : _GEN_59660; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_59665 = 5'h3 == _T_5904 ? w_vn_3 : 5'h0; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_59666 = 5'h4 == _T_5904 ? w_vn_4 : _GEN_59665; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_59667 = 5'h5 == _T_5904 ? 5'h0 : _GEN_59666; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_59668 = 5'h6 == _T_5904 ? 5'h0 : _GEN_59667; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_59669 = 5'h7 == _T_5904 ? w_vn_7 : _GEN_59668; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_59670 = 5'h8 == _T_5904 ? w_vn_8 : _GEN_59669; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_59671 = 5'h9 == _T_5904 ? 5'h0 : _GEN_59670; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_59672 = 5'ha == _T_5904 ? 5'h0 : _GEN_59671; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_59673 = 5'hb == _T_5904 ? w_vn_11 : _GEN_59672; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_59674 = 5'hc == _T_5904 ? w_vn_12 : _GEN_59673; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_59675 = 5'hd == _T_5904 ? w_vn_13 : _GEN_59674; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_59676 = 5'he == _T_5904 ? 5'h0 : _GEN_59675; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_59677 = 5'hf == _T_5904 ? w_vn_15 : _GEN_59676; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_59678 = 5'h10 == _T_5904 ? w_vn_16 : _GEN_59677; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_59679 = 5'h11 == _T_5904 ? 5'h0 : _GEN_59678; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_59680 = 5'h12 == _T_5904 ? w_vn_18 : _GEN_59679; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_59681 = 5'h13 == _T_5904 ? 5'h0 : _GEN_59680; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_59682 = 5'h14 == _T_5904 ? 5'h0 : _GEN_59681; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_59683 = 5'h15 == _T_5904 ? 5'h0 : _GEN_59682; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_59684 = 5'h16 == _T_5904 ? 5'h0 : _GEN_59683; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_59685 = 5'h17 == _T_5904 ? w_vn_23 : _GEN_59684; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_59686 = 5'h18 == _T_5904 ? w_vn_24 : _GEN_59685; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_59687 = 5'h19 == _T_5904 ? 5'h0 : _GEN_59686; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_59688 = 5'h1a == _T_5904 ? 5'h0 : _GEN_59687; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_59689 = 5'h1b == _T_5904 ? 5'h0 : _GEN_59688; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_59690 = 5'h1c == _T_5904 ? 5'h0 : _GEN_59689; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_59691 = 5'h1d == _T_5904 ? 5'h0 : _GEN_59690; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_59692 = 5'h1e == _T_5904 ? 5'h0 : _GEN_59691; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_59693 = 5'h1f == _T_5904 ? 5'h0 : _GEN_59692; // @[FanCtrl.scala 282:{37,37}]
  wire  _T_5905 = _GEN_59661 == _GEN_59693; // @[FanCtrl.scala 282:37]
  wire [4:0] _T_5908 = _T_5888 + 5'h5; // @[FanCtrl.scala 283:29]
  wire [4:0] _T_5911 = _T_5888 + 5'h6; // @[FanCtrl.scala 283:56]
  wire [4:0] _GEN_59697 = 5'h3 == _T_5908 ? w_vn_3 : 5'h0; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_59698 = 5'h4 == _T_5908 ? w_vn_4 : _GEN_59697; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_59699 = 5'h5 == _T_5908 ? 5'h0 : _GEN_59698; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_59700 = 5'h6 == _T_5908 ? 5'h0 : _GEN_59699; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_59701 = 5'h7 == _T_5908 ? w_vn_7 : _GEN_59700; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_59702 = 5'h8 == _T_5908 ? w_vn_8 : _GEN_59701; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_59703 = 5'h9 == _T_5908 ? 5'h0 : _GEN_59702; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_59704 = 5'ha == _T_5908 ? 5'h0 : _GEN_59703; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_59705 = 5'hb == _T_5908 ? w_vn_11 : _GEN_59704; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_59706 = 5'hc == _T_5908 ? w_vn_12 : _GEN_59705; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_59707 = 5'hd == _T_5908 ? w_vn_13 : _GEN_59706; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_59708 = 5'he == _T_5908 ? 5'h0 : _GEN_59707; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_59709 = 5'hf == _T_5908 ? w_vn_15 : _GEN_59708; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_59710 = 5'h10 == _T_5908 ? w_vn_16 : _GEN_59709; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_59711 = 5'h11 == _T_5908 ? 5'h0 : _GEN_59710; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_59712 = 5'h12 == _T_5908 ? w_vn_18 : _GEN_59711; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_59713 = 5'h13 == _T_5908 ? 5'h0 : _GEN_59712; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_59714 = 5'h14 == _T_5908 ? 5'h0 : _GEN_59713; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_59715 = 5'h15 == _T_5908 ? 5'h0 : _GEN_59714; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_59716 = 5'h16 == _T_5908 ? 5'h0 : _GEN_59715; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_59717 = 5'h17 == _T_5908 ? w_vn_23 : _GEN_59716; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_59718 = 5'h18 == _T_5908 ? w_vn_24 : _GEN_59717; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_59719 = 5'h19 == _T_5908 ? 5'h0 : _GEN_59718; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_59720 = 5'h1a == _T_5908 ? 5'h0 : _GEN_59719; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_59721 = 5'h1b == _T_5908 ? 5'h0 : _GEN_59720; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_59722 = 5'h1c == _T_5908 ? 5'h0 : _GEN_59721; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_59723 = 5'h1d == _T_5908 ? 5'h0 : _GEN_59722; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_59724 = 5'h1e == _T_5908 ? 5'h0 : _GEN_59723; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_59725 = 5'h1f == _T_5908 ? 5'h0 : _GEN_59724; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_59729 = 5'h3 == _T_5911 ? w_vn_3 : 5'h0; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_59730 = 5'h4 == _T_5911 ? w_vn_4 : _GEN_59729; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_59731 = 5'h5 == _T_5911 ? 5'h0 : _GEN_59730; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_59732 = 5'h6 == _T_5911 ? 5'h0 : _GEN_59731; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_59733 = 5'h7 == _T_5911 ? w_vn_7 : _GEN_59732; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_59734 = 5'h8 == _T_5911 ? w_vn_8 : _GEN_59733; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_59735 = 5'h9 == _T_5911 ? 5'h0 : _GEN_59734; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_59736 = 5'ha == _T_5911 ? 5'h0 : _GEN_59735; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_59737 = 5'hb == _T_5911 ? w_vn_11 : _GEN_59736; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_59738 = 5'hc == _T_5911 ? w_vn_12 : _GEN_59737; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_59739 = 5'hd == _T_5911 ? w_vn_13 : _GEN_59738; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_59740 = 5'he == _T_5911 ? 5'h0 : _GEN_59739; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_59741 = 5'hf == _T_5911 ? w_vn_15 : _GEN_59740; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_59742 = 5'h10 == _T_5911 ? w_vn_16 : _GEN_59741; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_59743 = 5'h11 == _T_5911 ? 5'h0 : _GEN_59742; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_59744 = 5'h12 == _T_5911 ? w_vn_18 : _GEN_59743; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_59745 = 5'h13 == _T_5911 ? 5'h0 : _GEN_59744; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_59746 = 5'h14 == _T_5911 ? 5'h0 : _GEN_59745; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_59747 = 5'h15 == _T_5911 ? 5'h0 : _GEN_59746; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_59748 = 5'h16 == _T_5911 ? 5'h0 : _GEN_59747; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_59749 = 5'h17 == _T_5911 ? w_vn_23 : _GEN_59748; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_59750 = 5'h18 == _T_5911 ? w_vn_24 : _GEN_59749; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_59751 = 5'h19 == _T_5911 ? 5'h0 : _GEN_59750; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_59752 = 5'h1a == _T_5911 ? 5'h0 : _GEN_59751; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_59753 = 5'h1b == _T_5911 ? 5'h0 : _GEN_59752; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_59754 = 5'h1c == _T_5911 ? 5'h0 : _GEN_59753; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_59755 = 5'h1d == _T_5911 ? 5'h0 : _GEN_59754; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_59756 = 5'h1e == _T_5911 ? 5'h0 : _GEN_59755; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_59757 = 5'h1f == _T_5911 ? 5'h0 : _GEN_59756; // @[FanCtrl.scala 283:{37,37}]
  wire  _T_5912 = _GEN_59725 == _GEN_59757; // @[FanCtrl.scala 283:37]
  wire  _T_5913 = _GEN_59661 == _GEN_59693 & _T_5912; // @[FanCtrl.scala 282:64]
  wire [4:0] _T_5916 = _T_5888 + 5'h8; // @[FanCtrl.scala 284:29]
  wire [4:0] _GEN_59761 = 5'h3 == _T_5916 ? w_vn_3 : 5'h0; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_59762 = 5'h4 == _T_5916 ? w_vn_4 : _GEN_59761; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_59763 = 5'h5 == _T_5916 ? 5'h0 : _GEN_59762; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_59764 = 5'h6 == _T_5916 ? 5'h0 : _GEN_59763; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_59765 = 5'h7 == _T_5916 ? w_vn_7 : _GEN_59764; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_59766 = 5'h8 == _T_5916 ? w_vn_8 : _GEN_59765; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_59767 = 5'h9 == _T_5916 ? 5'h0 : _GEN_59766; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_59768 = 5'ha == _T_5916 ? 5'h0 : _GEN_59767; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_59769 = 5'hb == _T_5916 ? w_vn_11 : _GEN_59768; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_59770 = 5'hc == _T_5916 ? w_vn_12 : _GEN_59769; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_59771 = 5'hd == _T_5916 ? w_vn_13 : _GEN_59770; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_59772 = 5'he == _T_5916 ? 5'h0 : _GEN_59771; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_59773 = 5'hf == _T_5916 ? w_vn_15 : _GEN_59772; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_59774 = 5'h10 == _T_5916 ? w_vn_16 : _GEN_59773; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_59775 = 5'h11 == _T_5916 ? 5'h0 : _GEN_59774; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_59776 = 5'h12 == _T_5916 ? w_vn_18 : _GEN_59775; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_59777 = 5'h13 == _T_5916 ? 5'h0 : _GEN_59776; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_59778 = 5'h14 == _T_5916 ? 5'h0 : _GEN_59777; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_59779 = 5'h15 == _T_5916 ? 5'h0 : _GEN_59778; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_59780 = 5'h16 == _T_5916 ? 5'h0 : _GEN_59779; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_59781 = 5'h17 == _T_5916 ? w_vn_23 : _GEN_59780; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_59782 = 5'h18 == _T_5916 ? w_vn_24 : _GEN_59781; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_59783 = 5'h19 == _T_5916 ? 5'h0 : _GEN_59782; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_59784 = 5'h1a == _T_5916 ? 5'h0 : _GEN_59783; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_59785 = 5'h1b == _T_5916 ? 5'h0 : _GEN_59784; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_59786 = 5'h1c == _T_5916 ? 5'h0 : _GEN_59785; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_59787 = 5'h1d == _T_5916 ? 5'h0 : _GEN_59786; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_59788 = 5'h1e == _T_5916 ? 5'h0 : _GEN_59787; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_59789 = 5'h1f == _T_5916 ? 5'h0 : _GEN_59788; // @[FanCtrl.scala 284:{36,36}]
  wire  _T_5920 = _GEN_59789 != _GEN_59757; // @[FanCtrl.scala 284:36]
  wire  _T_5921 = _T_5913 & _T_5920; // @[FanCtrl.scala 283:64]
  wire  _T_5928 = _GEN_59693 != _GEN_59536; // @[FanCtrl.scala 285:36]
  wire  _T_5929 = _T_5921 & _T_5928; // @[FanCtrl.scala 284:64]
  wire  _T_5936 = _GEN_59725 != _GEN_59504; // @[FanCtrl.scala 286:37]
  wire  _T_5937 = _T_5929 & _T_5936; // @[FanCtrl.scala 285:64]
  wire  _T_5954 = _T_5912 & _T_5920; // @[FanCtrl.scala 290:71]
  wire  _T_5962 = _T_5954 & _T_5936; // @[FanCtrl.scala 291:70]
  wire  _T_5979 = _T_5905 & _T_5928; // @[FanCtrl.scala 296:72]
  wire [2:0] _GEN_60418 = _T_5979 ? 3'h3 : 3'h0; // @[FanCtrl.scala 297:71]
  wire [2:0] _GEN_60449 = _T_5962 ? 3'h4 : _GEN_60418; // @[FanCtrl.scala 292:72]
  wire [2:0] _GEN_60480 = _T_5937 ? 3'h5 : _GEN_60449; // @[FanCtrl.scala 286:65]
  wire  _GEN_60573 = r_valid_1 & _T_5894; // @[FanCtrl.scala 274:32]
  wire [2:0] _GEN_60604 = r_valid_1 ? _GEN_60480 : 3'h0; // @[FanCtrl.scala 274:32]
  wire [1:0] _GEN_60715 = _GEN_59504 == _GEN_59661 ? 2'h0 : 2'h1; // @[FanCtrl.scala 313:69]
  wire [1:0] _GEN_60755 = r_valid_1 ? _GEN_60715 : 2'h0; // @[FanCtrl.scala 312:32]
  wire [1:0] _GEN_60880 = _GEN_59536 == _GEN_59757 ? 2'h1 : 2'h0; // @[FanCtrl.scala 325:67]
  wire [1:0] _GEN_60919 = r_valid_1 ? _GEN_60755 : 2'h0; // @[FanCtrl.scala 324:32]
  wire [1:0] _GEN_60920 = r_valid_1 ? _GEN_60880 : r_reduction_sel_1; // @[FanCtrl.scala 324:32]
  wire [4:0] _T_6325 = 4'h8 * 1'h1; // @[FanCtrl.scala 276:23]
  wire [4:0] _T_6327 = _T_6325 + 5'h3; // @[FanCtrl.scala 276:29]
  wire [4:0] _T_6330 = _T_6325 + 5'h4; // @[FanCtrl.scala 276:56]
  wire [4:0] _GEN_64412 = 5'h3 == _T_6327 ? w_vn_3 : 5'h0; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_64413 = 5'h4 == _T_6327 ? w_vn_4 : _GEN_64412; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_64414 = 5'h5 == _T_6327 ? 5'h0 : _GEN_64413; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_64415 = 5'h6 == _T_6327 ? 5'h0 : _GEN_64414; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_64416 = 5'h7 == _T_6327 ? w_vn_7 : _GEN_64415; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_64417 = 5'h8 == _T_6327 ? w_vn_8 : _GEN_64416; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_64418 = 5'h9 == _T_6327 ? 5'h0 : _GEN_64417; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_64419 = 5'ha == _T_6327 ? 5'h0 : _GEN_64418; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_64420 = 5'hb == _T_6327 ? w_vn_11 : _GEN_64419; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_64421 = 5'hc == _T_6327 ? w_vn_12 : _GEN_64420; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_64422 = 5'hd == _T_6327 ? w_vn_13 : _GEN_64421; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_64423 = 5'he == _T_6327 ? 5'h0 : _GEN_64422; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_64424 = 5'hf == _T_6327 ? w_vn_15 : _GEN_64423; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_64425 = 5'h10 == _T_6327 ? w_vn_16 : _GEN_64424; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_64426 = 5'h11 == _T_6327 ? 5'h0 : _GEN_64425; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_64427 = 5'h12 == _T_6327 ? w_vn_18 : _GEN_64426; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_64428 = 5'h13 == _T_6327 ? 5'h0 : _GEN_64427; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_64429 = 5'h14 == _T_6327 ? 5'h0 : _GEN_64428; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_64430 = 5'h15 == _T_6327 ? 5'h0 : _GEN_64429; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_64431 = 5'h16 == _T_6327 ? 5'h0 : _GEN_64430; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_64432 = 5'h17 == _T_6327 ? w_vn_23 : _GEN_64431; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_64433 = 5'h18 == _T_6327 ? w_vn_24 : _GEN_64432; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_64434 = 5'h19 == _T_6327 ? 5'h0 : _GEN_64433; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_64435 = 5'h1a == _T_6327 ? 5'h0 : _GEN_64434; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_64436 = 5'h1b == _T_6327 ? 5'h0 : _GEN_64435; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_64437 = 5'h1c == _T_6327 ? 5'h0 : _GEN_64436; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_64438 = 5'h1d == _T_6327 ? 5'h0 : _GEN_64437; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_64439 = 5'h1e == _T_6327 ? 5'h0 : _GEN_64438; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_64440 = 5'h1f == _T_6327 ? 5'h0 : _GEN_64439; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_64444 = 5'h3 == _T_6330 ? w_vn_3 : 5'h0; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_64445 = 5'h4 == _T_6330 ? w_vn_4 : _GEN_64444; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_64446 = 5'h5 == _T_6330 ? 5'h0 : _GEN_64445; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_64447 = 5'h6 == _T_6330 ? 5'h0 : _GEN_64446; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_64448 = 5'h7 == _T_6330 ? w_vn_7 : _GEN_64447; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_64449 = 5'h8 == _T_6330 ? w_vn_8 : _GEN_64448; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_64450 = 5'h9 == _T_6330 ? 5'h0 : _GEN_64449; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_64451 = 5'ha == _T_6330 ? 5'h0 : _GEN_64450; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_64452 = 5'hb == _T_6330 ? w_vn_11 : _GEN_64451; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_64453 = 5'hc == _T_6330 ? w_vn_12 : _GEN_64452; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_64454 = 5'hd == _T_6330 ? w_vn_13 : _GEN_64453; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_64455 = 5'he == _T_6330 ? 5'h0 : _GEN_64454; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_64456 = 5'hf == _T_6330 ? w_vn_15 : _GEN_64455; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_64457 = 5'h10 == _T_6330 ? w_vn_16 : _GEN_64456; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_64458 = 5'h11 == _T_6330 ? 5'h0 : _GEN_64457; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_64459 = 5'h12 == _T_6330 ? w_vn_18 : _GEN_64458; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_64460 = 5'h13 == _T_6330 ? 5'h0 : _GEN_64459; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_64461 = 5'h14 == _T_6330 ? 5'h0 : _GEN_64460; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_64462 = 5'h15 == _T_6330 ? 5'h0 : _GEN_64461; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_64463 = 5'h16 == _T_6330 ? 5'h0 : _GEN_64462; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_64464 = 5'h17 == _T_6330 ? w_vn_23 : _GEN_64463; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_64465 = 5'h18 == _T_6330 ? w_vn_24 : _GEN_64464; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_64466 = 5'h19 == _T_6330 ? 5'h0 : _GEN_64465; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_64467 = 5'h1a == _T_6330 ? 5'h0 : _GEN_64466; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_64468 = 5'h1b == _T_6330 ? 5'h0 : _GEN_64467; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_64469 = 5'h1c == _T_6330 ? 5'h0 : _GEN_64468; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_64470 = 5'h1d == _T_6330 ? 5'h0 : _GEN_64469; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_64471 = 5'h1e == _T_6330 ? 5'h0 : _GEN_64470; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_64472 = 5'h1f == _T_6330 ? 5'h0 : _GEN_64471; // @[FanCtrl.scala 276:{37,37}]
  wire  _T_6331 = _GEN_64440 == _GEN_64472; // @[FanCtrl.scala 276:37]
  wire [4:0] _T_6338 = _T_6325 + 5'h1; // @[FanCtrl.scala 282:30]
  wire [4:0] _T_6341 = _T_6325 + 5'h2; // @[FanCtrl.scala 282:56]
  wire [4:0] _GEN_64569 = 5'h3 == _T_6338 ? w_vn_3 : 5'h0; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_64570 = 5'h4 == _T_6338 ? w_vn_4 : _GEN_64569; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_64571 = 5'h5 == _T_6338 ? 5'h0 : _GEN_64570; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_64572 = 5'h6 == _T_6338 ? 5'h0 : _GEN_64571; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_64573 = 5'h7 == _T_6338 ? w_vn_7 : _GEN_64572; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_64574 = 5'h8 == _T_6338 ? w_vn_8 : _GEN_64573; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_64575 = 5'h9 == _T_6338 ? 5'h0 : _GEN_64574; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_64576 = 5'ha == _T_6338 ? 5'h0 : _GEN_64575; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_64577 = 5'hb == _T_6338 ? w_vn_11 : _GEN_64576; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_64578 = 5'hc == _T_6338 ? w_vn_12 : _GEN_64577; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_64579 = 5'hd == _T_6338 ? w_vn_13 : _GEN_64578; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_64580 = 5'he == _T_6338 ? 5'h0 : _GEN_64579; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_64581 = 5'hf == _T_6338 ? w_vn_15 : _GEN_64580; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_64582 = 5'h10 == _T_6338 ? w_vn_16 : _GEN_64581; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_64583 = 5'h11 == _T_6338 ? 5'h0 : _GEN_64582; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_64584 = 5'h12 == _T_6338 ? w_vn_18 : _GEN_64583; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_64585 = 5'h13 == _T_6338 ? 5'h0 : _GEN_64584; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_64586 = 5'h14 == _T_6338 ? 5'h0 : _GEN_64585; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_64587 = 5'h15 == _T_6338 ? 5'h0 : _GEN_64586; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_64588 = 5'h16 == _T_6338 ? 5'h0 : _GEN_64587; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_64589 = 5'h17 == _T_6338 ? w_vn_23 : _GEN_64588; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_64590 = 5'h18 == _T_6338 ? w_vn_24 : _GEN_64589; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_64591 = 5'h19 == _T_6338 ? 5'h0 : _GEN_64590; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_64592 = 5'h1a == _T_6338 ? 5'h0 : _GEN_64591; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_64593 = 5'h1b == _T_6338 ? 5'h0 : _GEN_64592; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_64594 = 5'h1c == _T_6338 ? 5'h0 : _GEN_64593; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_64595 = 5'h1d == _T_6338 ? 5'h0 : _GEN_64594; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_64596 = 5'h1e == _T_6338 ? 5'h0 : _GEN_64595; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_64597 = 5'h1f == _T_6338 ? 5'h0 : _GEN_64596; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_64601 = 5'h3 == _T_6341 ? w_vn_3 : 5'h0; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_64602 = 5'h4 == _T_6341 ? w_vn_4 : _GEN_64601; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_64603 = 5'h5 == _T_6341 ? 5'h0 : _GEN_64602; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_64604 = 5'h6 == _T_6341 ? 5'h0 : _GEN_64603; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_64605 = 5'h7 == _T_6341 ? w_vn_7 : _GEN_64604; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_64606 = 5'h8 == _T_6341 ? w_vn_8 : _GEN_64605; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_64607 = 5'h9 == _T_6341 ? 5'h0 : _GEN_64606; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_64608 = 5'ha == _T_6341 ? 5'h0 : _GEN_64607; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_64609 = 5'hb == _T_6341 ? w_vn_11 : _GEN_64608; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_64610 = 5'hc == _T_6341 ? w_vn_12 : _GEN_64609; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_64611 = 5'hd == _T_6341 ? w_vn_13 : _GEN_64610; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_64612 = 5'he == _T_6341 ? 5'h0 : _GEN_64611; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_64613 = 5'hf == _T_6341 ? w_vn_15 : _GEN_64612; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_64614 = 5'h10 == _T_6341 ? w_vn_16 : _GEN_64613; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_64615 = 5'h11 == _T_6341 ? 5'h0 : _GEN_64614; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_64616 = 5'h12 == _T_6341 ? w_vn_18 : _GEN_64615; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_64617 = 5'h13 == _T_6341 ? 5'h0 : _GEN_64616; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_64618 = 5'h14 == _T_6341 ? 5'h0 : _GEN_64617; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_64619 = 5'h15 == _T_6341 ? 5'h0 : _GEN_64618; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_64620 = 5'h16 == _T_6341 ? 5'h0 : _GEN_64619; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_64621 = 5'h17 == _T_6341 ? w_vn_23 : _GEN_64620; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_64622 = 5'h18 == _T_6341 ? w_vn_24 : _GEN_64621; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_64623 = 5'h19 == _T_6341 ? 5'h0 : _GEN_64622; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_64624 = 5'h1a == _T_6341 ? 5'h0 : _GEN_64623; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_64625 = 5'h1b == _T_6341 ? 5'h0 : _GEN_64624; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_64626 = 5'h1c == _T_6341 ? 5'h0 : _GEN_64625; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_64627 = 5'h1d == _T_6341 ? 5'h0 : _GEN_64626; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_64628 = 5'h1e == _T_6341 ? 5'h0 : _GEN_64627; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_64629 = 5'h1f == _T_6341 ? 5'h0 : _GEN_64628; // @[FanCtrl.scala 282:{37,37}]
  wire  _T_6342 = _GEN_64597 == _GEN_64629; // @[FanCtrl.scala 282:37]
  wire [4:0] _T_6345 = _T_6325 + 5'h5; // @[FanCtrl.scala 283:29]
  wire [4:0] _T_6348 = _T_6325 + 5'h6; // @[FanCtrl.scala 283:56]
  wire [4:0] _GEN_64633 = 5'h3 == _T_6345 ? w_vn_3 : 5'h0; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_64634 = 5'h4 == _T_6345 ? w_vn_4 : _GEN_64633; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_64635 = 5'h5 == _T_6345 ? 5'h0 : _GEN_64634; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_64636 = 5'h6 == _T_6345 ? 5'h0 : _GEN_64635; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_64637 = 5'h7 == _T_6345 ? w_vn_7 : _GEN_64636; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_64638 = 5'h8 == _T_6345 ? w_vn_8 : _GEN_64637; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_64639 = 5'h9 == _T_6345 ? 5'h0 : _GEN_64638; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_64640 = 5'ha == _T_6345 ? 5'h0 : _GEN_64639; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_64641 = 5'hb == _T_6345 ? w_vn_11 : _GEN_64640; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_64642 = 5'hc == _T_6345 ? w_vn_12 : _GEN_64641; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_64643 = 5'hd == _T_6345 ? w_vn_13 : _GEN_64642; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_64644 = 5'he == _T_6345 ? 5'h0 : _GEN_64643; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_64645 = 5'hf == _T_6345 ? w_vn_15 : _GEN_64644; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_64646 = 5'h10 == _T_6345 ? w_vn_16 : _GEN_64645; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_64647 = 5'h11 == _T_6345 ? 5'h0 : _GEN_64646; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_64648 = 5'h12 == _T_6345 ? w_vn_18 : _GEN_64647; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_64649 = 5'h13 == _T_6345 ? 5'h0 : _GEN_64648; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_64650 = 5'h14 == _T_6345 ? 5'h0 : _GEN_64649; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_64651 = 5'h15 == _T_6345 ? 5'h0 : _GEN_64650; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_64652 = 5'h16 == _T_6345 ? 5'h0 : _GEN_64651; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_64653 = 5'h17 == _T_6345 ? w_vn_23 : _GEN_64652; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_64654 = 5'h18 == _T_6345 ? w_vn_24 : _GEN_64653; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_64655 = 5'h19 == _T_6345 ? 5'h0 : _GEN_64654; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_64656 = 5'h1a == _T_6345 ? 5'h0 : _GEN_64655; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_64657 = 5'h1b == _T_6345 ? 5'h0 : _GEN_64656; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_64658 = 5'h1c == _T_6345 ? 5'h0 : _GEN_64657; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_64659 = 5'h1d == _T_6345 ? 5'h0 : _GEN_64658; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_64660 = 5'h1e == _T_6345 ? 5'h0 : _GEN_64659; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_64661 = 5'h1f == _T_6345 ? 5'h0 : _GEN_64660; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_64665 = 5'h3 == _T_6348 ? w_vn_3 : 5'h0; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_64666 = 5'h4 == _T_6348 ? w_vn_4 : _GEN_64665; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_64667 = 5'h5 == _T_6348 ? 5'h0 : _GEN_64666; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_64668 = 5'h6 == _T_6348 ? 5'h0 : _GEN_64667; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_64669 = 5'h7 == _T_6348 ? w_vn_7 : _GEN_64668; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_64670 = 5'h8 == _T_6348 ? w_vn_8 : _GEN_64669; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_64671 = 5'h9 == _T_6348 ? 5'h0 : _GEN_64670; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_64672 = 5'ha == _T_6348 ? 5'h0 : _GEN_64671; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_64673 = 5'hb == _T_6348 ? w_vn_11 : _GEN_64672; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_64674 = 5'hc == _T_6348 ? w_vn_12 : _GEN_64673; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_64675 = 5'hd == _T_6348 ? w_vn_13 : _GEN_64674; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_64676 = 5'he == _T_6348 ? 5'h0 : _GEN_64675; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_64677 = 5'hf == _T_6348 ? w_vn_15 : _GEN_64676; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_64678 = 5'h10 == _T_6348 ? w_vn_16 : _GEN_64677; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_64679 = 5'h11 == _T_6348 ? 5'h0 : _GEN_64678; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_64680 = 5'h12 == _T_6348 ? w_vn_18 : _GEN_64679; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_64681 = 5'h13 == _T_6348 ? 5'h0 : _GEN_64680; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_64682 = 5'h14 == _T_6348 ? 5'h0 : _GEN_64681; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_64683 = 5'h15 == _T_6348 ? 5'h0 : _GEN_64682; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_64684 = 5'h16 == _T_6348 ? 5'h0 : _GEN_64683; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_64685 = 5'h17 == _T_6348 ? w_vn_23 : _GEN_64684; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_64686 = 5'h18 == _T_6348 ? w_vn_24 : _GEN_64685; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_64687 = 5'h19 == _T_6348 ? 5'h0 : _GEN_64686; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_64688 = 5'h1a == _T_6348 ? 5'h0 : _GEN_64687; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_64689 = 5'h1b == _T_6348 ? 5'h0 : _GEN_64688; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_64690 = 5'h1c == _T_6348 ? 5'h0 : _GEN_64689; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_64691 = 5'h1d == _T_6348 ? 5'h0 : _GEN_64690; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_64692 = 5'h1e == _T_6348 ? 5'h0 : _GEN_64691; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_64693 = 5'h1f == _T_6348 ? 5'h0 : _GEN_64692; // @[FanCtrl.scala 283:{37,37}]
  wire  _T_6349 = _GEN_64661 == _GEN_64693; // @[FanCtrl.scala 283:37]
  wire  _T_6350 = _GEN_64597 == _GEN_64629 & _T_6349; // @[FanCtrl.scala 282:64]
  wire [4:0] _T_6353 = _T_6325 + 5'h8; // @[FanCtrl.scala 284:29]
  wire [4:0] _GEN_64697 = 5'h3 == _T_6353 ? w_vn_3 : 5'h0; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_64698 = 5'h4 == _T_6353 ? w_vn_4 : _GEN_64697; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_64699 = 5'h5 == _T_6353 ? 5'h0 : _GEN_64698; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_64700 = 5'h6 == _T_6353 ? 5'h0 : _GEN_64699; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_64701 = 5'h7 == _T_6353 ? w_vn_7 : _GEN_64700; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_64702 = 5'h8 == _T_6353 ? w_vn_8 : _GEN_64701; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_64703 = 5'h9 == _T_6353 ? 5'h0 : _GEN_64702; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_64704 = 5'ha == _T_6353 ? 5'h0 : _GEN_64703; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_64705 = 5'hb == _T_6353 ? w_vn_11 : _GEN_64704; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_64706 = 5'hc == _T_6353 ? w_vn_12 : _GEN_64705; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_64707 = 5'hd == _T_6353 ? w_vn_13 : _GEN_64706; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_64708 = 5'he == _T_6353 ? 5'h0 : _GEN_64707; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_64709 = 5'hf == _T_6353 ? w_vn_15 : _GEN_64708; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_64710 = 5'h10 == _T_6353 ? w_vn_16 : _GEN_64709; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_64711 = 5'h11 == _T_6353 ? 5'h0 : _GEN_64710; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_64712 = 5'h12 == _T_6353 ? w_vn_18 : _GEN_64711; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_64713 = 5'h13 == _T_6353 ? 5'h0 : _GEN_64712; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_64714 = 5'h14 == _T_6353 ? 5'h0 : _GEN_64713; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_64715 = 5'h15 == _T_6353 ? 5'h0 : _GEN_64714; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_64716 = 5'h16 == _T_6353 ? 5'h0 : _GEN_64715; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_64717 = 5'h17 == _T_6353 ? w_vn_23 : _GEN_64716; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_64718 = 5'h18 == _T_6353 ? w_vn_24 : _GEN_64717; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_64719 = 5'h19 == _T_6353 ? 5'h0 : _GEN_64718; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_64720 = 5'h1a == _T_6353 ? 5'h0 : _GEN_64719; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_64721 = 5'h1b == _T_6353 ? 5'h0 : _GEN_64720; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_64722 = 5'h1c == _T_6353 ? 5'h0 : _GEN_64721; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_64723 = 5'h1d == _T_6353 ? 5'h0 : _GEN_64722; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_64724 = 5'h1e == _T_6353 ? 5'h0 : _GEN_64723; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_64725 = 5'h1f == _T_6353 ? 5'h0 : _GEN_64724; // @[FanCtrl.scala 284:{36,36}]
  wire  _T_6357 = _GEN_64725 != _GEN_64693; // @[FanCtrl.scala 284:36]
  wire  _T_6365 = _GEN_64629 != _GEN_64472; // @[FanCtrl.scala 285:36]
  wire  _T_6373 = _GEN_64661 != _GEN_64440; // @[FanCtrl.scala 286:37]
  wire  _T_6391 = _T_6349 & _T_6357; // @[FanCtrl.scala 290:71]
  wire  _T_6399 = _T_6391 & _T_6373; // @[FanCtrl.scala 291:70]
  wire  _GEN_65510 = r_valid_1 & _T_6331; // @[FanCtrl.scala 274:32]
  wire  _T_6432 = _GEN_64440 == _GEN_64597; // @[FanCtrl.scala 313:39]
  wire  _T_6446 = _GEN_64472 == _GEN_64693; // @[FanCtrl.scala 325:39]
  wire [2:0] _T_6458 = 1'h1 * 2'h2; // @[FanCtrl.scala 338:28]
  wire [3:0] _T_6459 = {{1'd0}, _T_6458}; // @[FanCtrl.scala 338:35]
  wire [1:0] _GEN_65937 = 3'h0 == _T_6459[2:0] ? 2'h0 : _GEN_60919; // @[FanCtrl.scala 338:{42,42}]
  wire [1:0] _GEN_65938 = 3'h1 == _T_6459[2:0] ? 2'h0 : _GEN_60920; // @[FanCtrl.scala 338:{42,42}]
  wire [1:0] _GEN_65939 = 3'h2 == _T_6459[2:0] ? 2'h0 : r_reduction_sel_2; // @[FanCtrl.scala 338:{42,42}]
  wire [1:0] _GEN_65940 = 3'h3 == _T_6459[2:0] ? 2'h0 : r_reduction_sel_3; // @[FanCtrl.scala 338:{42,42}]
  wire [1:0] _GEN_65941 = 3'h4 == _T_6459[2:0] ? 2'h0 : r_reduction_sel_4; // @[FanCtrl.scala 338:{42,42}]
  wire [1:0] _GEN_65942 = 3'h5 == _T_6459[2:0] ? 2'h0 : r_reduction_sel_5; // @[FanCtrl.scala 338:{42,42}]
  wire [1:0] _GEN_65943 = 3'h6 == _T_6459[2:0] ? 2'h0 : r_reduction_sel_6; // @[FanCtrl.scala 338:{42,42}]
  wire [1:0] _GEN_65944 = 3'h7 == _T_6459[2:0] ? 2'h0 : r_reduction_sel_7; // @[FanCtrl.scala 338:{42,42}]
  wire [3:0] _GEN_97590 = {{1'd0}, _T_6459[2:0]}; // @[FanCtrl.scala 338:{42,42}]
  wire [1:0] _GEN_65945 = 4'h8 == _GEN_97590 ? 2'h0 : r_reduction_sel_8; // @[FanCtrl.scala 338:{42,42}]
  wire [1:0] _GEN_65946 = 4'h9 == _GEN_97590 ? 2'h0 : r_reduction_sel_9; // @[FanCtrl.scala 338:{42,42}]
  wire [1:0] _GEN_65947 = 4'ha == _GEN_97590 ? 2'h0 : r_reduction_sel_10; // @[FanCtrl.scala 338:{42,42}]
  wire [1:0] _GEN_65948 = 4'hb == _GEN_97590 ? 2'h0 : r_reduction_sel_11; // @[FanCtrl.scala 338:{42,42}]
  wire [1:0] _GEN_65949 = 4'hc == _GEN_97590 ? 2'h0 : r_reduction_sel_12; // @[FanCtrl.scala 338:{42,42}]
  wire [1:0] _GEN_65950 = 4'hd == _GEN_97590 ? 2'h0 : r_reduction_sel_13; // @[FanCtrl.scala 338:{42,42}]
  wire [1:0] _GEN_65951 = 4'he == _GEN_97590 ? 2'h0 : r_reduction_sel_14; // @[FanCtrl.scala 338:{42,42}]
  wire [1:0] _GEN_65952 = 4'hf == _GEN_97590 ? 2'h0 : r_reduction_sel_15; // @[FanCtrl.scala 338:{42,42}]
  wire [4:0] _GEN_97598 = {{2'd0}, _T_6459[2:0]}; // @[FanCtrl.scala 338:{42,42}]
  wire [1:0] _GEN_65953 = 5'h10 == _GEN_97598 ? 2'h0 : r_reduction_sel_16; // @[FanCtrl.scala 338:{42,42}]
  wire [1:0] _GEN_65954 = 5'h11 == _GEN_97598 ? 2'h0 : r_reduction_sel_17; // @[FanCtrl.scala 338:{42,42}]
  wire [1:0] _GEN_65955 = 5'h12 == _GEN_97598 ? 2'h0 : r_reduction_sel_18; // @[FanCtrl.scala 338:{42,42}]
  wire [1:0] _GEN_65956 = 5'h13 == _GEN_97598 ? 2'h0 : r_reduction_sel_19; // @[FanCtrl.scala 338:{42,42}]
  wire [4:0] _T_6493 = _T_6325 - 5'h1; // @[FanCtrl.scala 349:58]
  wire [4:0] _GEN_66277 = 5'h3 == _T_6493 ? w_vn_3 : 5'h0; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_66278 = 5'h4 == _T_6493 ? w_vn_4 : _GEN_66277; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_66279 = 5'h5 == _T_6493 ? 5'h0 : _GEN_66278; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_66280 = 5'h6 == _T_6493 ? 5'h0 : _GEN_66279; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_66281 = 5'h7 == _T_6493 ? w_vn_7 : _GEN_66280; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_66282 = 5'h8 == _T_6493 ? w_vn_8 : _GEN_66281; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_66283 = 5'h9 == _T_6493 ? 5'h0 : _GEN_66282; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_66284 = 5'ha == _T_6493 ? 5'h0 : _GEN_66283; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_66285 = 5'hb == _T_6493 ? w_vn_11 : _GEN_66284; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_66286 = 5'hc == _T_6493 ? w_vn_12 : _GEN_66285; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_66287 = 5'hd == _T_6493 ? w_vn_13 : _GEN_66286; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_66288 = 5'he == _T_6493 ? 5'h0 : _GEN_66287; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_66289 = 5'hf == _T_6493 ? w_vn_15 : _GEN_66288; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_66290 = 5'h10 == _T_6493 ? w_vn_16 : _GEN_66289; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_66291 = 5'h11 == _T_6493 ? 5'h0 : _GEN_66290; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_66292 = 5'h12 == _T_6493 ? w_vn_18 : _GEN_66291; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_66293 = 5'h13 == _T_6493 ? 5'h0 : _GEN_66292; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_66294 = 5'h14 == _T_6493 ? 5'h0 : _GEN_66293; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_66295 = 5'h15 == _T_6493 ? 5'h0 : _GEN_66294; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_66296 = 5'h16 == _T_6493 ? 5'h0 : _GEN_66295; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_66297 = 5'h17 == _T_6493 ? w_vn_23 : _GEN_66296; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_66298 = 5'h18 == _T_6493 ? w_vn_24 : _GEN_66297; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_66299 = 5'h19 == _T_6493 ? 5'h0 : _GEN_66298; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_66300 = 5'h1a == _T_6493 ? 5'h0 : _GEN_66299; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_66301 = 5'h1b == _T_6493 ? 5'h0 : _GEN_66300; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_66302 = 5'h1c == _T_6493 ? 5'h0 : _GEN_66301; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_66303 = 5'h1d == _T_6493 ? 5'h0 : _GEN_66302; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_66304 = 5'h1e == _T_6493 ? 5'h0 : _GEN_66303; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_66305 = 5'h1f == _T_6493 ? 5'h0 : _GEN_66304; // @[FanCtrl.scala 349:{39,39}]
  wire  _T_6494 = _GEN_64597 != _GEN_66305; // @[FanCtrl.scala 349:39]
  wire  _T_6495 = _T_6350 & _T_6494; // @[FanCtrl.scala 348:67]
  wire  _T_6528 = _T_6342 & _T_6494; // @[FanCtrl.scala 355:73]
  wire  _T_6535 = _GEN_64472 != _GEN_64629; // @[FanCtrl.scala 357:42]
  wire  _T_6536 = _T_6528 & _T_6535; // @[FanCtrl.scala 356:71]
  wire [1:0] _GEN_67159 = 3'h0 == _T_6459[2:0] ? 2'h0 : _GEN_65937; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_67160 = 3'h1 == _T_6459[2:0] ? 2'h0 : _GEN_65938; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_67161 = 3'h2 == _T_6459[2:0] ? 2'h0 : _GEN_65939; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_67162 = 3'h3 == _T_6459[2:0] ? 2'h0 : _GEN_65940; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_67163 = 3'h4 == _T_6459[2:0] ? 2'h0 : _GEN_65941; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_67164 = 3'h5 == _T_6459[2:0] ? 2'h0 : _GEN_65942; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_67165 = 3'h6 == _T_6459[2:0] ? 2'h0 : _GEN_65943; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_67166 = 3'h7 == _T_6459[2:0] ? 2'h0 : _GEN_65944; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_67167 = 4'h8 == _GEN_97590 ? 2'h0 : _GEN_65945; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_67168 = 4'h9 == _GEN_97590 ? 2'h0 : _GEN_65946; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_67169 = 4'ha == _GEN_97590 ? 2'h0 : _GEN_65947; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_67170 = 4'hb == _GEN_97590 ? 2'h0 : _GEN_65948; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_67171 = 4'hc == _GEN_97590 ? 2'h0 : _GEN_65949; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_67172 = 4'hd == _GEN_97590 ? 2'h0 : _GEN_65950; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_67173 = 4'he == _GEN_97590 ? 2'h0 : _GEN_65951; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_67174 = 4'hf == _GEN_97590 ? 2'h0 : _GEN_65952; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_67175 = 5'h10 == _GEN_97598 ? 2'h0 : _GEN_65953; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_67176 = 5'h11 == _GEN_97598 ? 2'h0 : _GEN_65954; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_67177 = 5'h12 == _GEN_97598 ? 2'h0 : _GEN_65955; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_67178 = 5'h13 == _GEN_97598 ? 2'h0 : _GEN_65956; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_67179 = 3'h0 == _T_6459[2:0] ? 2'h1 : _GEN_65937; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_67180 = 3'h1 == _T_6459[2:0] ? 2'h1 : _GEN_65938; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_67181 = 3'h2 == _T_6459[2:0] ? 2'h1 : _GEN_65939; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_67182 = 3'h3 == _T_6459[2:0] ? 2'h1 : _GEN_65940; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_67183 = 3'h4 == _T_6459[2:0] ? 2'h1 : _GEN_65941; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_67184 = 3'h5 == _T_6459[2:0] ? 2'h1 : _GEN_65942; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_67185 = 3'h6 == _T_6459[2:0] ? 2'h1 : _GEN_65943; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_67186 = 3'h7 == _T_6459[2:0] ? 2'h1 : _GEN_65944; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_67187 = 4'h8 == _GEN_97590 ? 2'h1 : _GEN_65945; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_67188 = 4'h9 == _GEN_97590 ? 2'h1 : _GEN_65946; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_67189 = 4'ha == _GEN_97590 ? 2'h1 : _GEN_65947; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_67190 = 4'hb == _GEN_97590 ? 2'h1 : _GEN_65948; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_67191 = 4'hc == _GEN_97590 ? 2'h1 : _GEN_65949; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_67192 = 4'hd == _GEN_97590 ? 2'h1 : _GEN_65950; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_67193 = 4'he == _GEN_97590 ? 2'h1 : _GEN_65951; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_67194 = 4'hf == _GEN_97590 ? 2'h1 : _GEN_65952; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_67195 = 5'h10 == _GEN_97598 ? 2'h1 : _GEN_65953; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_67196 = 5'h11 == _GEN_97598 ? 2'h1 : _GEN_65954; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_67197 = 5'h12 == _GEN_97598 ? 2'h1 : _GEN_65955; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_67198 = 5'h13 == _GEN_97598 ? 2'h1 : _GEN_65956; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_67199 = _T_6432 ? _GEN_67159 : _GEN_67179; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_67200 = _T_6432 ? _GEN_67160 : _GEN_67180; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_67201 = _T_6432 ? _GEN_67161 : _GEN_67181; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_67202 = _T_6432 ? _GEN_67162 : _GEN_67182; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_67203 = _T_6432 ? _GEN_67163 : _GEN_67183; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_67204 = _T_6432 ? _GEN_67164 : _GEN_67184; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_67205 = _T_6432 ? _GEN_67165 : _GEN_67185; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_67206 = _T_6432 ? _GEN_67166 : _GEN_67186; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_67207 = _T_6432 ? _GEN_67167 : _GEN_67187; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_67208 = _T_6432 ? _GEN_67168 : _GEN_67188; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_67209 = _T_6432 ? _GEN_67169 : _GEN_67189; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_67210 = _T_6432 ? _GEN_67170 : _GEN_67190; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_67211 = _T_6432 ? _GEN_67171 : _GEN_67191; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_67212 = _T_6432 ? _GEN_67172 : _GEN_67192; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_67213 = _T_6432 ? _GEN_67173 : _GEN_67193; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_67214 = _T_6432 ? _GEN_67174 : _GEN_67194; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_67215 = _T_6432 ? _GEN_67175 : _GEN_67195; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_67216 = _T_6432 ? _GEN_67176 : _GEN_67196; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_67217 = _T_6432 ? _GEN_67177 : _GEN_67197; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_67218 = _T_6432 ? _GEN_67178 : _GEN_67198; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_67239 = r_valid_1 ? _GEN_67199 : _GEN_67159; // @[FanCtrl.scala 376:33]
  wire [1:0] _GEN_67240 = r_valid_1 ? _GEN_67200 : _GEN_67160; // @[FanCtrl.scala 376:33]
  wire [1:0] _GEN_67241 = r_valid_1 ? _GEN_67201 : _GEN_67161; // @[FanCtrl.scala 376:33]
  wire [1:0] _GEN_67242 = r_valid_1 ? _GEN_67202 : _GEN_67162; // @[FanCtrl.scala 376:33]
  wire [1:0] _GEN_67243 = r_valid_1 ? _GEN_67203 : _GEN_67163; // @[FanCtrl.scala 376:33]
  wire [1:0] _GEN_67244 = r_valid_1 ? _GEN_67204 : _GEN_67164; // @[FanCtrl.scala 376:33]
  wire [1:0] _GEN_67245 = r_valid_1 ? _GEN_67205 : _GEN_67165; // @[FanCtrl.scala 376:33]
  wire [1:0] _GEN_67246 = r_valid_1 ? _GEN_67206 : _GEN_67166; // @[FanCtrl.scala 376:33]
  wire [1:0] _GEN_67247 = r_valid_1 ? _GEN_67207 : _GEN_67167; // @[FanCtrl.scala 376:33]
  wire [1:0] _GEN_67248 = r_valid_1 ? _GEN_67208 : _GEN_67168; // @[FanCtrl.scala 376:33]
  wire [1:0] _GEN_67249 = r_valid_1 ? _GEN_67209 : _GEN_67169; // @[FanCtrl.scala 376:33]
  wire [1:0] _GEN_67250 = r_valid_1 ? _GEN_67210 : _GEN_67170; // @[FanCtrl.scala 376:33]
  wire [1:0] _GEN_67251 = r_valid_1 ? _GEN_67211 : _GEN_67171; // @[FanCtrl.scala 376:33]
  wire [1:0] _GEN_67252 = r_valid_1 ? _GEN_67212 : _GEN_67172; // @[FanCtrl.scala 376:33]
  wire [1:0] _GEN_67253 = r_valid_1 ? _GEN_67213 : _GEN_67173; // @[FanCtrl.scala 376:33]
  wire [1:0] _GEN_67254 = r_valid_1 ? _GEN_67214 : _GEN_67174; // @[FanCtrl.scala 376:33]
  wire [1:0] _GEN_67255 = r_valid_1 ? _GEN_67215 : _GEN_67175; // @[FanCtrl.scala 376:33]
  wire [1:0] _GEN_67256 = r_valid_1 ? _GEN_67216 : _GEN_67176; // @[FanCtrl.scala 376:33]
  wire [1:0] _GEN_67257 = r_valid_1 ? _GEN_67217 : _GEN_67177; // @[FanCtrl.scala 376:33]
  wire [1:0] _GEN_67258 = r_valid_1 ? _GEN_67218 : _GEN_67178; // @[FanCtrl.scala 376:33]
  wire [2:0] _T_6589 = _T_6458 + 3'h1; // @[FanCtrl.scala 392:39]
  wire [1:0] _GEN_67323 = 3'h0 == _T_6589 ? 2'h1 : _GEN_67239; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_67324 = 3'h1 == _T_6589 ? 2'h1 : _GEN_67240; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_67325 = 3'h2 == _T_6589 ? 2'h1 : _GEN_67241; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_67326 = 3'h3 == _T_6589 ? 2'h1 : _GEN_67242; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_67327 = 3'h4 == _T_6589 ? 2'h1 : _GEN_67243; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_67328 = 3'h5 == _T_6589 ? 2'h1 : _GEN_67244; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_67329 = 3'h6 == _T_6589 ? 2'h1 : _GEN_67245; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_67330 = 3'h7 == _T_6589 ? 2'h1 : _GEN_67246; // @[FanCtrl.scala 392:{46,46}]
  wire [3:0] _GEN_97638 = {{1'd0}, _T_6589}; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_67331 = 4'h8 == _GEN_97638 ? 2'h1 : _GEN_67247; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_67332 = 4'h9 == _GEN_97638 ? 2'h1 : _GEN_67248; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_67333 = 4'ha == _GEN_97638 ? 2'h1 : _GEN_67249; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_67334 = 4'hb == _GEN_97638 ? 2'h1 : _GEN_67250; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_67335 = 4'hc == _GEN_97638 ? 2'h1 : _GEN_67251; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_67336 = 4'hd == _GEN_97638 ? 2'h1 : _GEN_67252; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_67337 = 4'he == _GEN_97638 ? 2'h1 : _GEN_67253; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_67338 = 4'hf == _GEN_97638 ? 2'h1 : _GEN_67254; // @[FanCtrl.scala 392:{46,46}]
  wire [4:0] _GEN_97646 = {{2'd0}, _T_6589}; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_67339 = 5'h10 == _GEN_97646 ? 2'h1 : _GEN_67255; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_67340 = 5'h11 == _GEN_97646 ? 2'h1 : _GEN_67256; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_67341 = 5'h12 == _GEN_97646 ? 2'h1 : _GEN_67257; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_67342 = 5'h13 == _GEN_97646 ? 2'h1 : _GEN_67258; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_67343 = 3'h0 == _T_6589 ? 2'h0 : _GEN_67239; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_67344 = 3'h1 == _T_6589 ? 2'h0 : _GEN_67240; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_67345 = 3'h2 == _T_6589 ? 2'h0 : _GEN_67241; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_67346 = 3'h3 == _T_6589 ? 2'h0 : _GEN_67242; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_67347 = 3'h4 == _T_6589 ? 2'h0 : _GEN_67243; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_67348 = 3'h5 == _T_6589 ? 2'h0 : _GEN_67244; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_67349 = 3'h6 == _T_6589 ? 2'h0 : _GEN_67245; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_67350 = 3'h7 == _T_6589 ? 2'h0 : _GEN_67246; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_67351 = 4'h8 == _GEN_97638 ? 2'h0 : _GEN_67247; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_67352 = 4'h9 == _GEN_97638 ? 2'h0 : _GEN_67248; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_67353 = 4'ha == _GEN_97638 ? 2'h0 : _GEN_67249; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_67354 = 4'hb == _GEN_97638 ? 2'h0 : _GEN_67250; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_67355 = 4'hc == _GEN_97638 ? 2'h0 : _GEN_67251; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_67356 = 4'hd == _GEN_97638 ? 2'h0 : _GEN_67252; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_67357 = 4'he == _GEN_97638 ? 2'h0 : _GEN_67253; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_67358 = 4'hf == _GEN_97638 ? 2'h0 : _GEN_67254; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_67359 = 5'h10 == _GEN_97646 ? 2'h0 : _GEN_67255; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_67360 = 5'h11 == _GEN_97646 ? 2'h0 : _GEN_67256; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_67361 = 5'h12 == _GEN_97646 ? 2'h0 : _GEN_67257; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_67362 = 5'h13 == _GEN_97646 ? 2'h0 : _GEN_67258; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_67363 = _T_6446 ? _GEN_67323 : _GEN_67343; // @[FanCtrl.scala 390:64]
  wire [1:0] _GEN_67364 = _T_6446 ? _GEN_67324 : _GEN_67344; // @[FanCtrl.scala 390:64]
  wire [1:0] _GEN_67365 = _T_6446 ? _GEN_67325 : _GEN_67345; // @[FanCtrl.scala 390:64]
  wire [1:0] _GEN_67366 = _T_6446 ? _GEN_67326 : _GEN_67346; // @[FanCtrl.scala 390:64]
  wire [1:0] _GEN_67367 = _T_6446 ? _GEN_67327 : _GEN_67347; // @[FanCtrl.scala 390:64]
  wire [1:0] _GEN_67368 = _T_6446 ? _GEN_67328 : _GEN_67348; // @[FanCtrl.scala 390:64]
  wire [1:0] _GEN_67369 = _T_6446 ? _GEN_67329 : _GEN_67349; // @[FanCtrl.scala 390:64]
  wire [1:0] _GEN_67370 = _T_6446 ? _GEN_67330 : _GEN_67350; // @[FanCtrl.scala 390:64]
  wire [1:0] _GEN_67371 = _T_6446 ? _GEN_67331 : _GEN_67351; // @[FanCtrl.scala 390:64]
  wire [1:0] _GEN_67372 = _T_6446 ? _GEN_67332 : _GEN_67352; // @[FanCtrl.scala 390:64]
  wire [1:0] _GEN_67373 = _T_6446 ? _GEN_67333 : _GEN_67353; // @[FanCtrl.scala 390:64]
  wire [1:0] _GEN_67374 = _T_6446 ? _GEN_67334 : _GEN_67354; // @[FanCtrl.scala 390:64]
  wire [1:0] _GEN_67375 = _T_6446 ? _GEN_67335 : _GEN_67355; // @[FanCtrl.scala 390:64]
  wire [1:0] _GEN_67376 = _T_6446 ? _GEN_67336 : _GEN_67356; // @[FanCtrl.scala 390:64]
  wire [1:0] _GEN_67377 = _T_6446 ? _GEN_67337 : _GEN_67357; // @[FanCtrl.scala 390:64]
  wire [1:0] _GEN_67378 = _T_6446 ? _GEN_67338 : _GEN_67358; // @[FanCtrl.scala 390:64]
  wire [1:0] _GEN_67379 = _T_6446 ? _GEN_67339 : _GEN_67359; // @[FanCtrl.scala 390:64]
  wire [1:0] _GEN_67380 = _T_6446 ? _GEN_67340 : _GEN_67360; // @[FanCtrl.scala 390:64]
  wire [1:0] _GEN_67381 = _T_6446 ? _GEN_67341 : _GEN_67361; // @[FanCtrl.scala 390:64]
  wire [1:0] _GEN_67382 = _T_6446 ? _GEN_67342 : _GEN_67362; // @[FanCtrl.scala 390:64]
  wire  _T_6645 = _T_6495 & _T_6357; // @[FanCtrl.scala 417:67]
  wire  _T_6653 = _T_6645 & _T_6365; // @[FanCtrl.scala 418:66]
  wire  _T_6661 = _T_6653 & _T_6373; // @[FanCtrl.scala 419:66]
  wire [2:0] _GEN_68579 = _T_6536 ? 3'h3 : 3'h0; // @[FanCtrl.scala 432:71]
  wire [2:0] _GEN_68610 = _T_6399 ? 3'h4 : _GEN_68579; // @[FanCtrl.scala 426:72]
  wire [2:0] _GEN_68641 = _T_6661 ? 3'h5 : _GEN_68610; // @[FanCtrl.scala 420:67]
  wire [2:0] _GEN_68765 = r_valid_1 ? _GEN_68641 : 3'h0; // @[FanCtrl.scala 408:33]
  wire [1:0] _GEN_69079 = r_valid_1 ? _GEN_67363 : _GEN_67343; // @[FanCtrl.scala 459:33]
  wire [1:0] _GEN_69080 = r_valid_1 ? _GEN_67364 : _GEN_67344; // @[FanCtrl.scala 459:33]
  wire [1:0] _GEN_69081 = r_valid_1 ? _GEN_67365 : _GEN_67345; // @[FanCtrl.scala 459:33]
  wire [1:0] _GEN_69082 = r_valid_1 ? _GEN_67366 : _GEN_67346; // @[FanCtrl.scala 459:33]
  wire [1:0] _GEN_69083 = r_valid_1 ? _GEN_67367 : _GEN_67347; // @[FanCtrl.scala 459:33]
  wire [1:0] _GEN_69084 = r_valid_1 ? _GEN_67368 : _GEN_67348; // @[FanCtrl.scala 459:33]
  wire [1:0] _GEN_69085 = r_valid_1 ? _GEN_67369 : _GEN_67349; // @[FanCtrl.scala 459:33]
  wire [1:0] _GEN_69086 = r_valid_1 ? _GEN_67370 : _GEN_67350; // @[FanCtrl.scala 459:33]
  wire [1:0] _GEN_69087 = r_valid_1 ? _GEN_67371 : _GEN_67351; // @[FanCtrl.scala 459:33]
  wire [1:0] _GEN_69088 = r_valid_1 ? _GEN_67372 : _GEN_67352; // @[FanCtrl.scala 459:33]
  wire [1:0] _GEN_69089 = r_valid_1 ? _GEN_67373 : _GEN_67353; // @[FanCtrl.scala 459:33]
  wire [1:0] _GEN_69090 = r_valid_1 ? _GEN_67374 : _GEN_67354; // @[FanCtrl.scala 459:33]
  wire [1:0] _GEN_69091 = r_valid_1 ? _GEN_67375 : _GEN_67355; // @[FanCtrl.scala 459:33]
  wire [1:0] _GEN_69092 = r_valid_1 ? _GEN_67376 : _GEN_67356; // @[FanCtrl.scala 459:33]
  wire [1:0] _GEN_69093 = r_valid_1 ? _GEN_67377 : _GEN_67357; // @[FanCtrl.scala 459:33]
  wire [1:0] _GEN_69094 = r_valid_1 ? _GEN_67378 : _GEN_67358; // @[FanCtrl.scala 459:33]
  wire [1:0] _GEN_69095 = r_valid_1 ? _GEN_67379 : _GEN_67359; // @[FanCtrl.scala 459:33]
  wire [1:0] _GEN_69096 = r_valid_1 ? _GEN_67380 : _GEN_67360; // @[FanCtrl.scala 459:33]
  wire [1:0] _GEN_69097 = r_valid_1 ? _GEN_67381 : _GEN_67361; // @[FanCtrl.scala 459:33]
  wire [1:0] _GEN_69098 = r_valid_1 ? _GEN_67382 : _GEN_67362; // @[FanCtrl.scala 459:33]
  wire [5:0] _T_6762 = 4'h8 * 2'h2; // @[FanCtrl.scala 276:23]
  wire [5:0] _T_6764 = _T_6762 + 6'h3; // @[FanCtrl.scala 276:29]
  wire [5:0] _T_6768 = _T_6762 + 6'h4; // @[FanCtrl.scala 276:56]
  wire [4:0] _GEN_69348 = 5'h3 == _T_6764[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_69349 = 5'h4 == _T_6764[4:0] ? w_vn_4 : _GEN_69348; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_69350 = 5'h5 == _T_6764[4:0] ? 5'h0 : _GEN_69349; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_69351 = 5'h6 == _T_6764[4:0] ? 5'h0 : _GEN_69350; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_69352 = 5'h7 == _T_6764[4:0] ? w_vn_7 : _GEN_69351; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_69353 = 5'h8 == _T_6764[4:0] ? w_vn_8 : _GEN_69352; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_69354 = 5'h9 == _T_6764[4:0] ? 5'h0 : _GEN_69353; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_69355 = 5'ha == _T_6764[4:0] ? 5'h0 : _GEN_69354; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_69356 = 5'hb == _T_6764[4:0] ? w_vn_11 : _GEN_69355; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_69357 = 5'hc == _T_6764[4:0] ? w_vn_12 : _GEN_69356; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_69358 = 5'hd == _T_6764[4:0] ? w_vn_13 : _GEN_69357; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_69359 = 5'he == _T_6764[4:0] ? 5'h0 : _GEN_69358; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_69360 = 5'hf == _T_6764[4:0] ? w_vn_15 : _GEN_69359; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_69361 = 5'h10 == _T_6764[4:0] ? w_vn_16 : _GEN_69360; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_69362 = 5'h11 == _T_6764[4:0] ? 5'h0 : _GEN_69361; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_69363 = 5'h12 == _T_6764[4:0] ? w_vn_18 : _GEN_69362; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_69364 = 5'h13 == _T_6764[4:0] ? 5'h0 : _GEN_69363; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_69365 = 5'h14 == _T_6764[4:0] ? 5'h0 : _GEN_69364; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_69366 = 5'h15 == _T_6764[4:0] ? 5'h0 : _GEN_69365; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_69367 = 5'h16 == _T_6764[4:0] ? 5'h0 : _GEN_69366; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_69368 = 5'h17 == _T_6764[4:0] ? w_vn_23 : _GEN_69367; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_69369 = 5'h18 == _T_6764[4:0] ? w_vn_24 : _GEN_69368; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_69370 = 5'h19 == _T_6764[4:0] ? 5'h0 : _GEN_69369; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_69371 = 5'h1a == _T_6764[4:0] ? 5'h0 : _GEN_69370; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_69372 = 5'h1b == _T_6764[4:0] ? 5'h0 : _GEN_69371; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_69373 = 5'h1c == _T_6764[4:0] ? 5'h0 : _GEN_69372; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_69374 = 5'h1d == _T_6764[4:0] ? 5'h0 : _GEN_69373; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_69375 = 5'h1e == _T_6764[4:0] ? 5'h0 : _GEN_69374; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_69376 = 5'h1f == _T_6764[4:0] ? 5'h0 : _GEN_69375; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_69380 = 5'h3 == _T_6768[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_69381 = 5'h4 == _T_6768[4:0] ? w_vn_4 : _GEN_69380; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_69382 = 5'h5 == _T_6768[4:0] ? 5'h0 : _GEN_69381; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_69383 = 5'h6 == _T_6768[4:0] ? 5'h0 : _GEN_69382; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_69384 = 5'h7 == _T_6768[4:0] ? w_vn_7 : _GEN_69383; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_69385 = 5'h8 == _T_6768[4:0] ? w_vn_8 : _GEN_69384; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_69386 = 5'h9 == _T_6768[4:0] ? 5'h0 : _GEN_69385; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_69387 = 5'ha == _T_6768[4:0] ? 5'h0 : _GEN_69386; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_69388 = 5'hb == _T_6768[4:0] ? w_vn_11 : _GEN_69387; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_69389 = 5'hc == _T_6768[4:0] ? w_vn_12 : _GEN_69388; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_69390 = 5'hd == _T_6768[4:0] ? w_vn_13 : _GEN_69389; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_69391 = 5'he == _T_6768[4:0] ? 5'h0 : _GEN_69390; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_69392 = 5'hf == _T_6768[4:0] ? w_vn_15 : _GEN_69391; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_69393 = 5'h10 == _T_6768[4:0] ? w_vn_16 : _GEN_69392; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_69394 = 5'h11 == _T_6768[4:0] ? 5'h0 : _GEN_69393; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_69395 = 5'h12 == _T_6768[4:0] ? w_vn_18 : _GEN_69394; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_69396 = 5'h13 == _T_6768[4:0] ? 5'h0 : _GEN_69395; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_69397 = 5'h14 == _T_6768[4:0] ? 5'h0 : _GEN_69396; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_69398 = 5'h15 == _T_6768[4:0] ? 5'h0 : _GEN_69397; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_69399 = 5'h16 == _T_6768[4:0] ? 5'h0 : _GEN_69398; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_69400 = 5'h17 == _T_6768[4:0] ? w_vn_23 : _GEN_69399; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_69401 = 5'h18 == _T_6768[4:0] ? w_vn_24 : _GEN_69400; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_69402 = 5'h19 == _T_6768[4:0] ? 5'h0 : _GEN_69401; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_69403 = 5'h1a == _T_6768[4:0] ? 5'h0 : _GEN_69402; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_69404 = 5'h1b == _T_6768[4:0] ? 5'h0 : _GEN_69403; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_69405 = 5'h1c == _T_6768[4:0] ? 5'h0 : _GEN_69404; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_69406 = 5'h1d == _T_6768[4:0] ? 5'h0 : _GEN_69405; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_69407 = 5'h1e == _T_6768[4:0] ? 5'h0 : _GEN_69406; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_69408 = 5'h1f == _T_6768[4:0] ? 5'h0 : _GEN_69407; // @[FanCtrl.scala 276:{37,37}]
  wire  _T_6770 = _GEN_69376 == _GEN_69408; // @[FanCtrl.scala 276:37]
  wire [5:0] _T_6777 = _T_6762 + 6'h1; // @[FanCtrl.scala 282:30]
  wire [5:0] _T_6781 = _T_6762 + 6'h2; // @[FanCtrl.scala 282:56]
  wire [4:0] _GEN_69505 = 5'h3 == _T_6777[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_69506 = 5'h4 == _T_6777[4:0] ? w_vn_4 : _GEN_69505; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_69507 = 5'h5 == _T_6777[4:0] ? 5'h0 : _GEN_69506; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_69508 = 5'h6 == _T_6777[4:0] ? 5'h0 : _GEN_69507; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_69509 = 5'h7 == _T_6777[4:0] ? w_vn_7 : _GEN_69508; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_69510 = 5'h8 == _T_6777[4:0] ? w_vn_8 : _GEN_69509; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_69511 = 5'h9 == _T_6777[4:0] ? 5'h0 : _GEN_69510; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_69512 = 5'ha == _T_6777[4:0] ? 5'h0 : _GEN_69511; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_69513 = 5'hb == _T_6777[4:0] ? w_vn_11 : _GEN_69512; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_69514 = 5'hc == _T_6777[4:0] ? w_vn_12 : _GEN_69513; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_69515 = 5'hd == _T_6777[4:0] ? w_vn_13 : _GEN_69514; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_69516 = 5'he == _T_6777[4:0] ? 5'h0 : _GEN_69515; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_69517 = 5'hf == _T_6777[4:0] ? w_vn_15 : _GEN_69516; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_69518 = 5'h10 == _T_6777[4:0] ? w_vn_16 : _GEN_69517; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_69519 = 5'h11 == _T_6777[4:0] ? 5'h0 : _GEN_69518; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_69520 = 5'h12 == _T_6777[4:0] ? w_vn_18 : _GEN_69519; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_69521 = 5'h13 == _T_6777[4:0] ? 5'h0 : _GEN_69520; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_69522 = 5'h14 == _T_6777[4:0] ? 5'h0 : _GEN_69521; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_69523 = 5'h15 == _T_6777[4:0] ? 5'h0 : _GEN_69522; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_69524 = 5'h16 == _T_6777[4:0] ? 5'h0 : _GEN_69523; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_69525 = 5'h17 == _T_6777[4:0] ? w_vn_23 : _GEN_69524; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_69526 = 5'h18 == _T_6777[4:0] ? w_vn_24 : _GEN_69525; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_69527 = 5'h19 == _T_6777[4:0] ? 5'h0 : _GEN_69526; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_69528 = 5'h1a == _T_6777[4:0] ? 5'h0 : _GEN_69527; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_69529 = 5'h1b == _T_6777[4:0] ? 5'h0 : _GEN_69528; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_69530 = 5'h1c == _T_6777[4:0] ? 5'h0 : _GEN_69529; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_69531 = 5'h1d == _T_6777[4:0] ? 5'h0 : _GEN_69530; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_69532 = 5'h1e == _T_6777[4:0] ? 5'h0 : _GEN_69531; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_69533 = 5'h1f == _T_6777[4:0] ? 5'h0 : _GEN_69532; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_69537 = 5'h3 == _T_6781[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_69538 = 5'h4 == _T_6781[4:0] ? w_vn_4 : _GEN_69537; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_69539 = 5'h5 == _T_6781[4:0] ? 5'h0 : _GEN_69538; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_69540 = 5'h6 == _T_6781[4:0] ? 5'h0 : _GEN_69539; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_69541 = 5'h7 == _T_6781[4:0] ? w_vn_7 : _GEN_69540; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_69542 = 5'h8 == _T_6781[4:0] ? w_vn_8 : _GEN_69541; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_69543 = 5'h9 == _T_6781[4:0] ? 5'h0 : _GEN_69542; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_69544 = 5'ha == _T_6781[4:0] ? 5'h0 : _GEN_69543; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_69545 = 5'hb == _T_6781[4:0] ? w_vn_11 : _GEN_69544; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_69546 = 5'hc == _T_6781[4:0] ? w_vn_12 : _GEN_69545; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_69547 = 5'hd == _T_6781[4:0] ? w_vn_13 : _GEN_69546; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_69548 = 5'he == _T_6781[4:0] ? 5'h0 : _GEN_69547; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_69549 = 5'hf == _T_6781[4:0] ? w_vn_15 : _GEN_69548; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_69550 = 5'h10 == _T_6781[4:0] ? w_vn_16 : _GEN_69549; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_69551 = 5'h11 == _T_6781[4:0] ? 5'h0 : _GEN_69550; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_69552 = 5'h12 == _T_6781[4:0] ? w_vn_18 : _GEN_69551; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_69553 = 5'h13 == _T_6781[4:0] ? 5'h0 : _GEN_69552; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_69554 = 5'h14 == _T_6781[4:0] ? 5'h0 : _GEN_69553; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_69555 = 5'h15 == _T_6781[4:0] ? 5'h0 : _GEN_69554; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_69556 = 5'h16 == _T_6781[4:0] ? 5'h0 : _GEN_69555; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_69557 = 5'h17 == _T_6781[4:0] ? w_vn_23 : _GEN_69556; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_69558 = 5'h18 == _T_6781[4:0] ? w_vn_24 : _GEN_69557; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_69559 = 5'h19 == _T_6781[4:0] ? 5'h0 : _GEN_69558; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_69560 = 5'h1a == _T_6781[4:0] ? 5'h0 : _GEN_69559; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_69561 = 5'h1b == _T_6781[4:0] ? 5'h0 : _GEN_69560; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_69562 = 5'h1c == _T_6781[4:0] ? 5'h0 : _GEN_69561; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_69563 = 5'h1d == _T_6781[4:0] ? 5'h0 : _GEN_69562; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_69564 = 5'h1e == _T_6781[4:0] ? 5'h0 : _GEN_69563; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_69565 = 5'h1f == _T_6781[4:0] ? 5'h0 : _GEN_69564; // @[FanCtrl.scala 282:{37,37}]
  wire  _T_6783 = _GEN_69533 == _GEN_69565; // @[FanCtrl.scala 282:37]
  wire [5:0] _T_6786 = _T_6762 + 6'h5; // @[FanCtrl.scala 283:29]
  wire [5:0] _T_6790 = _T_6762 + 6'h6; // @[FanCtrl.scala 283:56]
  wire [4:0] _GEN_69569 = 5'h3 == _T_6786[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_69570 = 5'h4 == _T_6786[4:0] ? w_vn_4 : _GEN_69569; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_69571 = 5'h5 == _T_6786[4:0] ? 5'h0 : _GEN_69570; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_69572 = 5'h6 == _T_6786[4:0] ? 5'h0 : _GEN_69571; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_69573 = 5'h7 == _T_6786[4:0] ? w_vn_7 : _GEN_69572; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_69574 = 5'h8 == _T_6786[4:0] ? w_vn_8 : _GEN_69573; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_69575 = 5'h9 == _T_6786[4:0] ? 5'h0 : _GEN_69574; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_69576 = 5'ha == _T_6786[4:0] ? 5'h0 : _GEN_69575; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_69577 = 5'hb == _T_6786[4:0] ? w_vn_11 : _GEN_69576; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_69578 = 5'hc == _T_6786[4:0] ? w_vn_12 : _GEN_69577; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_69579 = 5'hd == _T_6786[4:0] ? w_vn_13 : _GEN_69578; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_69580 = 5'he == _T_6786[4:0] ? 5'h0 : _GEN_69579; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_69581 = 5'hf == _T_6786[4:0] ? w_vn_15 : _GEN_69580; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_69582 = 5'h10 == _T_6786[4:0] ? w_vn_16 : _GEN_69581; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_69583 = 5'h11 == _T_6786[4:0] ? 5'h0 : _GEN_69582; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_69584 = 5'h12 == _T_6786[4:0] ? w_vn_18 : _GEN_69583; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_69585 = 5'h13 == _T_6786[4:0] ? 5'h0 : _GEN_69584; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_69586 = 5'h14 == _T_6786[4:0] ? 5'h0 : _GEN_69585; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_69587 = 5'h15 == _T_6786[4:0] ? 5'h0 : _GEN_69586; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_69588 = 5'h16 == _T_6786[4:0] ? 5'h0 : _GEN_69587; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_69589 = 5'h17 == _T_6786[4:0] ? w_vn_23 : _GEN_69588; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_69590 = 5'h18 == _T_6786[4:0] ? w_vn_24 : _GEN_69589; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_69591 = 5'h19 == _T_6786[4:0] ? 5'h0 : _GEN_69590; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_69592 = 5'h1a == _T_6786[4:0] ? 5'h0 : _GEN_69591; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_69593 = 5'h1b == _T_6786[4:0] ? 5'h0 : _GEN_69592; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_69594 = 5'h1c == _T_6786[4:0] ? 5'h0 : _GEN_69593; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_69595 = 5'h1d == _T_6786[4:0] ? 5'h0 : _GEN_69594; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_69596 = 5'h1e == _T_6786[4:0] ? 5'h0 : _GEN_69595; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_69597 = 5'h1f == _T_6786[4:0] ? 5'h0 : _GEN_69596; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_69601 = 5'h3 == _T_6790[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_69602 = 5'h4 == _T_6790[4:0] ? w_vn_4 : _GEN_69601; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_69603 = 5'h5 == _T_6790[4:0] ? 5'h0 : _GEN_69602; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_69604 = 5'h6 == _T_6790[4:0] ? 5'h0 : _GEN_69603; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_69605 = 5'h7 == _T_6790[4:0] ? w_vn_7 : _GEN_69604; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_69606 = 5'h8 == _T_6790[4:0] ? w_vn_8 : _GEN_69605; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_69607 = 5'h9 == _T_6790[4:0] ? 5'h0 : _GEN_69606; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_69608 = 5'ha == _T_6790[4:0] ? 5'h0 : _GEN_69607; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_69609 = 5'hb == _T_6790[4:0] ? w_vn_11 : _GEN_69608; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_69610 = 5'hc == _T_6790[4:0] ? w_vn_12 : _GEN_69609; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_69611 = 5'hd == _T_6790[4:0] ? w_vn_13 : _GEN_69610; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_69612 = 5'he == _T_6790[4:0] ? 5'h0 : _GEN_69611; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_69613 = 5'hf == _T_6790[4:0] ? w_vn_15 : _GEN_69612; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_69614 = 5'h10 == _T_6790[4:0] ? w_vn_16 : _GEN_69613; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_69615 = 5'h11 == _T_6790[4:0] ? 5'h0 : _GEN_69614; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_69616 = 5'h12 == _T_6790[4:0] ? w_vn_18 : _GEN_69615; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_69617 = 5'h13 == _T_6790[4:0] ? 5'h0 : _GEN_69616; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_69618 = 5'h14 == _T_6790[4:0] ? 5'h0 : _GEN_69617; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_69619 = 5'h15 == _T_6790[4:0] ? 5'h0 : _GEN_69618; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_69620 = 5'h16 == _T_6790[4:0] ? 5'h0 : _GEN_69619; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_69621 = 5'h17 == _T_6790[4:0] ? w_vn_23 : _GEN_69620; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_69622 = 5'h18 == _T_6790[4:0] ? w_vn_24 : _GEN_69621; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_69623 = 5'h19 == _T_6790[4:0] ? 5'h0 : _GEN_69622; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_69624 = 5'h1a == _T_6790[4:0] ? 5'h0 : _GEN_69623; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_69625 = 5'h1b == _T_6790[4:0] ? 5'h0 : _GEN_69624; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_69626 = 5'h1c == _T_6790[4:0] ? 5'h0 : _GEN_69625; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_69627 = 5'h1d == _T_6790[4:0] ? 5'h0 : _GEN_69626; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_69628 = 5'h1e == _T_6790[4:0] ? 5'h0 : _GEN_69627; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_69629 = 5'h1f == _T_6790[4:0] ? 5'h0 : _GEN_69628; // @[FanCtrl.scala 283:{37,37}]
  wire  _T_6792 = _GEN_69597 == _GEN_69629; // @[FanCtrl.scala 283:37]
  wire  _T_6793 = _GEN_69533 == _GEN_69565 & _T_6792; // @[FanCtrl.scala 282:64]
  wire [5:0] _T_6796 = _T_6762 + 6'h8; // @[FanCtrl.scala 284:29]
  wire [4:0] _GEN_69633 = 5'h3 == _T_6796[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_69634 = 5'h4 == _T_6796[4:0] ? w_vn_4 : _GEN_69633; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_69635 = 5'h5 == _T_6796[4:0] ? 5'h0 : _GEN_69634; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_69636 = 5'h6 == _T_6796[4:0] ? 5'h0 : _GEN_69635; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_69637 = 5'h7 == _T_6796[4:0] ? w_vn_7 : _GEN_69636; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_69638 = 5'h8 == _T_6796[4:0] ? w_vn_8 : _GEN_69637; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_69639 = 5'h9 == _T_6796[4:0] ? 5'h0 : _GEN_69638; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_69640 = 5'ha == _T_6796[4:0] ? 5'h0 : _GEN_69639; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_69641 = 5'hb == _T_6796[4:0] ? w_vn_11 : _GEN_69640; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_69642 = 5'hc == _T_6796[4:0] ? w_vn_12 : _GEN_69641; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_69643 = 5'hd == _T_6796[4:0] ? w_vn_13 : _GEN_69642; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_69644 = 5'he == _T_6796[4:0] ? 5'h0 : _GEN_69643; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_69645 = 5'hf == _T_6796[4:0] ? w_vn_15 : _GEN_69644; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_69646 = 5'h10 == _T_6796[4:0] ? w_vn_16 : _GEN_69645; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_69647 = 5'h11 == _T_6796[4:0] ? 5'h0 : _GEN_69646; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_69648 = 5'h12 == _T_6796[4:0] ? w_vn_18 : _GEN_69647; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_69649 = 5'h13 == _T_6796[4:0] ? 5'h0 : _GEN_69648; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_69650 = 5'h14 == _T_6796[4:0] ? 5'h0 : _GEN_69649; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_69651 = 5'h15 == _T_6796[4:0] ? 5'h0 : _GEN_69650; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_69652 = 5'h16 == _T_6796[4:0] ? 5'h0 : _GEN_69651; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_69653 = 5'h17 == _T_6796[4:0] ? w_vn_23 : _GEN_69652; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_69654 = 5'h18 == _T_6796[4:0] ? w_vn_24 : _GEN_69653; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_69655 = 5'h19 == _T_6796[4:0] ? 5'h0 : _GEN_69654; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_69656 = 5'h1a == _T_6796[4:0] ? 5'h0 : _GEN_69655; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_69657 = 5'h1b == _T_6796[4:0] ? 5'h0 : _GEN_69656; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_69658 = 5'h1c == _T_6796[4:0] ? 5'h0 : _GEN_69657; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_69659 = 5'h1d == _T_6796[4:0] ? 5'h0 : _GEN_69658; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_69660 = 5'h1e == _T_6796[4:0] ? 5'h0 : _GEN_69659; // @[FanCtrl.scala 284:{36,36}]
  wire [4:0] _GEN_69661 = 5'h1f == _T_6796[4:0] ? 5'h0 : _GEN_69660; // @[FanCtrl.scala 284:{36,36}]
  wire  _T_6802 = _GEN_69661 != _GEN_69629; // @[FanCtrl.scala 284:36]
  wire  _T_6812 = _GEN_69565 != _GEN_69408; // @[FanCtrl.scala 285:36]
  wire  _T_6822 = _GEN_69597 != _GEN_69376; // @[FanCtrl.scala 286:37]
  wire  _T_6844 = _T_6792 & _T_6802; // @[FanCtrl.scala 290:71]
  wire  _T_6854 = _T_6844 & _T_6822; // @[FanCtrl.scala 291:70]
  wire  _GEN_70447 = r_valid_1 & _T_6770; // @[FanCtrl.scala 274:32]
  wire  _T_6893 = _GEN_69376 == _GEN_69533; // @[FanCtrl.scala 313:39]
  wire  _T_6909 = _GEN_69408 == _GEN_69629; // @[FanCtrl.scala 325:39]
  wire [1:0] _GEN_70873 = 4'h0 == _T_357[3:0] ? 2'h0 : _GEN_69079; // @[FanCtrl.scala 338:{42,42}]
  wire [1:0] _GEN_70874 = 4'h1 == _T_357[3:0] ? 2'h0 : _GEN_69080; // @[FanCtrl.scala 338:{42,42}]
  wire [1:0] _GEN_70875 = 4'h2 == _T_357[3:0] ? 2'h0 : _GEN_69081; // @[FanCtrl.scala 338:{42,42}]
  wire [1:0] _GEN_70876 = 4'h3 == _T_357[3:0] ? 2'h0 : _GEN_69082; // @[FanCtrl.scala 338:{42,42}]
  wire [1:0] _GEN_70877 = 4'h4 == _T_357[3:0] ? 2'h0 : _GEN_69083; // @[FanCtrl.scala 338:{42,42}]
  wire [1:0] _GEN_70878 = 4'h5 == _T_357[3:0] ? 2'h0 : _GEN_69084; // @[FanCtrl.scala 338:{42,42}]
  wire [1:0] _GEN_70879 = 4'h6 == _T_357[3:0] ? 2'h0 : _GEN_69085; // @[FanCtrl.scala 338:{42,42}]
  wire [1:0] _GEN_70880 = 4'h7 == _T_357[3:0] ? 2'h0 : _GEN_69086; // @[FanCtrl.scala 338:{42,42}]
  wire [1:0] _GEN_70881 = 4'h8 == _T_357[3:0] ? 2'h0 : _GEN_69087; // @[FanCtrl.scala 338:{42,42}]
  wire [1:0] _GEN_70882 = 4'h9 == _T_357[3:0] ? 2'h0 : _GEN_69088; // @[FanCtrl.scala 338:{42,42}]
  wire [1:0] _GEN_70883 = 4'ha == _T_357[3:0] ? 2'h0 : _GEN_69089; // @[FanCtrl.scala 338:{42,42}]
  wire [1:0] _GEN_70884 = 4'hb == _T_357[3:0] ? 2'h0 : _GEN_69090; // @[FanCtrl.scala 338:{42,42}]
  wire [1:0] _GEN_70885 = 4'hc == _T_357[3:0] ? 2'h0 : _GEN_69091; // @[FanCtrl.scala 338:{42,42}]
  wire [1:0] _GEN_70886 = 4'hd == _T_357[3:0] ? 2'h0 : _GEN_69092; // @[FanCtrl.scala 338:{42,42}]
  wire [1:0] _GEN_70887 = 4'he == _T_357[3:0] ? 2'h0 : _GEN_69093; // @[FanCtrl.scala 338:{42,42}]
  wire [1:0] _GEN_70888 = 4'hf == _T_357[3:0] ? 2'h0 : _GEN_69094; // @[FanCtrl.scala 338:{42,42}]
  wire [1:0] _GEN_70889 = 5'h10 == _GEN_94094 ? 2'h0 : _GEN_69095; // @[FanCtrl.scala 338:{42,42}]
  wire [1:0] _GEN_70890 = 5'h11 == _GEN_94094 ? 2'h0 : _GEN_69096; // @[FanCtrl.scala 338:{42,42}]
  wire [1:0] _GEN_70891 = 5'h12 == _GEN_94094 ? 2'h0 : _GEN_69097; // @[FanCtrl.scala 338:{42,42}]
  wire [1:0] _GEN_70892 = 5'h13 == _GEN_94094 ? 2'h0 : _GEN_69098; // @[FanCtrl.scala 338:{42,42}]
  wire [5:0] _T_6963 = _T_6762 - 6'h1; // @[FanCtrl.scala 349:58]
  wire [4:0] _GEN_71213 = 5'h3 == _T_6963[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_71214 = 5'h4 == _T_6963[4:0] ? w_vn_4 : _GEN_71213; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_71215 = 5'h5 == _T_6963[4:0] ? 5'h0 : _GEN_71214; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_71216 = 5'h6 == _T_6963[4:0] ? 5'h0 : _GEN_71215; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_71217 = 5'h7 == _T_6963[4:0] ? w_vn_7 : _GEN_71216; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_71218 = 5'h8 == _T_6963[4:0] ? w_vn_8 : _GEN_71217; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_71219 = 5'h9 == _T_6963[4:0] ? 5'h0 : _GEN_71218; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_71220 = 5'ha == _T_6963[4:0] ? 5'h0 : _GEN_71219; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_71221 = 5'hb == _T_6963[4:0] ? w_vn_11 : _GEN_71220; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_71222 = 5'hc == _T_6963[4:0] ? w_vn_12 : _GEN_71221; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_71223 = 5'hd == _T_6963[4:0] ? w_vn_13 : _GEN_71222; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_71224 = 5'he == _T_6963[4:0] ? 5'h0 : _GEN_71223; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_71225 = 5'hf == _T_6963[4:0] ? w_vn_15 : _GEN_71224; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_71226 = 5'h10 == _T_6963[4:0] ? w_vn_16 : _GEN_71225; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_71227 = 5'h11 == _T_6963[4:0] ? 5'h0 : _GEN_71226; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_71228 = 5'h12 == _T_6963[4:0] ? w_vn_18 : _GEN_71227; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_71229 = 5'h13 == _T_6963[4:0] ? 5'h0 : _GEN_71228; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_71230 = 5'h14 == _T_6963[4:0] ? 5'h0 : _GEN_71229; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_71231 = 5'h15 == _T_6963[4:0] ? 5'h0 : _GEN_71230; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_71232 = 5'h16 == _T_6963[4:0] ? 5'h0 : _GEN_71231; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_71233 = 5'h17 == _T_6963[4:0] ? w_vn_23 : _GEN_71232; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_71234 = 5'h18 == _T_6963[4:0] ? w_vn_24 : _GEN_71233; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_71235 = 5'h19 == _T_6963[4:0] ? 5'h0 : _GEN_71234; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_71236 = 5'h1a == _T_6963[4:0] ? 5'h0 : _GEN_71235; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_71237 = 5'h1b == _T_6963[4:0] ? 5'h0 : _GEN_71236; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_71238 = 5'h1c == _T_6963[4:0] ? 5'h0 : _GEN_71237; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_71239 = 5'h1d == _T_6963[4:0] ? 5'h0 : _GEN_71238; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_71240 = 5'h1e == _T_6963[4:0] ? 5'h0 : _GEN_71239; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_71241 = 5'h1f == _T_6963[4:0] ? 5'h0 : _GEN_71240; // @[FanCtrl.scala 349:{39,39}]
  wire  _T_6965 = _GEN_69533 != _GEN_71241; // @[FanCtrl.scala 349:39]
  wire  _T_6966 = _T_6793 & _T_6965; // @[FanCtrl.scala 348:67]
  wire  _T_7007 = _T_6783 & _T_6965; // @[FanCtrl.scala 355:73]
  wire  _T_7016 = _GEN_69408 != _GEN_69565; // @[FanCtrl.scala 357:42]
  wire  _T_7017 = _T_7007 & _T_7016; // @[FanCtrl.scala 356:71]
  wire [1:0] _GEN_72095 = 4'h0 == _T_357[3:0] ? 2'h0 : _GEN_70873; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_72096 = 4'h1 == _T_357[3:0] ? 2'h0 : _GEN_70874; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_72097 = 4'h2 == _T_357[3:0] ? 2'h0 : _GEN_70875; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_72098 = 4'h3 == _T_357[3:0] ? 2'h0 : _GEN_70876; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_72099 = 4'h4 == _T_357[3:0] ? 2'h0 : _GEN_70877; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_72100 = 4'h5 == _T_357[3:0] ? 2'h0 : _GEN_70878; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_72101 = 4'h6 == _T_357[3:0] ? 2'h0 : _GEN_70879; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_72102 = 4'h7 == _T_357[3:0] ? 2'h0 : _GEN_70880; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_72103 = 4'h8 == _T_357[3:0] ? 2'h0 : _GEN_70881; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_72104 = 4'h9 == _T_357[3:0] ? 2'h0 : _GEN_70882; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_72105 = 4'ha == _T_357[3:0] ? 2'h0 : _GEN_70883; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_72106 = 4'hb == _T_357[3:0] ? 2'h0 : _GEN_70884; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_72107 = 4'hc == _T_357[3:0] ? 2'h0 : _GEN_70885; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_72108 = 4'hd == _T_357[3:0] ? 2'h0 : _GEN_70886; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_72109 = 4'he == _T_357[3:0] ? 2'h0 : _GEN_70887; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_72110 = 4'hf == _T_357[3:0] ? 2'h0 : _GEN_70888; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_72111 = 5'h10 == _GEN_94094 ? 2'h0 : _GEN_70889; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_72112 = 5'h11 == _GEN_94094 ? 2'h0 : _GEN_70890; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_72113 = 5'h12 == _GEN_94094 ? 2'h0 : _GEN_70891; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_72114 = 5'h13 == _GEN_94094 ? 2'h0 : _GEN_70892; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_72115 = 4'h0 == _T_357[3:0] ? 2'h1 : _GEN_70873; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_72116 = 4'h1 == _T_357[3:0] ? 2'h1 : _GEN_70874; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_72117 = 4'h2 == _T_357[3:0] ? 2'h1 : _GEN_70875; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_72118 = 4'h3 == _T_357[3:0] ? 2'h1 : _GEN_70876; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_72119 = 4'h4 == _T_357[3:0] ? 2'h1 : _GEN_70877; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_72120 = 4'h5 == _T_357[3:0] ? 2'h1 : _GEN_70878; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_72121 = 4'h6 == _T_357[3:0] ? 2'h1 : _GEN_70879; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_72122 = 4'h7 == _T_357[3:0] ? 2'h1 : _GEN_70880; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_72123 = 4'h8 == _T_357[3:0] ? 2'h1 : _GEN_70881; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_72124 = 4'h9 == _T_357[3:0] ? 2'h1 : _GEN_70882; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_72125 = 4'ha == _T_357[3:0] ? 2'h1 : _GEN_70883; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_72126 = 4'hb == _T_357[3:0] ? 2'h1 : _GEN_70884; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_72127 = 4'hc == _T_357[3:0] ? 2'h1 : _GEN_70885; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_72128 = 4'hd == _T_357[3:0] ? 2'h1 : _GEN_70886; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_72129 = 4'he == _T_357[3:0] ? 2'h1 : _GEN_70887; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_72130 = 4'hf == _T_357[3:0] ? 2'h1 : _GEN_70888; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_72131 = 5'h10 == _GEN_94094 ? 2'h1 : _GEN_70889; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_72132 = 5'h11 == _GEN_94094 ? 2'h1 : _GEN_70890; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_72133 = 5'h12 == _GEN_94094 ? 2'h1 : _GEN_70891; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_72134 = 5'h13 == _GEN_94094 ? 2'h1 : _GEN_70892; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_72135 = _T_6893 ? _GEN_72095 : _GEN_72115; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_72136 = _T_6893 ? _GEN_72096 : _GEN_72116; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_72137 = _T_6893 ? _GEN_72097 : _GEN_72117; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_72138 = _T_6893 ? _GEN_72098 : _GEN_72118; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_72139 = _T_6893 ? _GEN_72099 : _GEN_72119; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_72140 = _T_6893 ? _GEN_72100 : _GEN_72120; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_72141 = _T_6893 ? _GEN_72101 : _GEN_72121; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_72142 = _T_6893 ? _GEN_72102 : _GEN_72122; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_72143 = _T_6893 ? _GEN_72103 : _GEN_72123; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_72144 = _T_6893 ? _GEN_72104 : _GEN_72124; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_72145 = _T_6893 ? _GEN_72105 : _GEN_72125; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_72146 = _T_6893 ? _GEN_72106 : _GEN_72126; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_72147 = _T_6893 ? _GEN_72107 : _GEN_72127; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_72148 = _T_6893 ? _GEN_72108 : _GEN_72128; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_72149 = _T_6893 ? _GEN_72109 : _GEN_72129; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_72150 = _T_6893 ? _GEN_72110 : _GEN_72130; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_72151 = _T_6893 ? _GEN_72111 : _GEN_72131; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_72152 = _T_6893 ? _GEN_72112 : _GEN_72132; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_72153 = _T_6893 ? _GEN_72113 : _GEN_72133; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_72154 = _T_6893 ? _GEN_72114 : _GEN_72134; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_72175 = r_valid_1 ? _GEN_72135 : _GEN_72095; // @[FanCtrl.scala 376:33]
  wire [1:0] _GEN_72176 = r_valid_1 ? _GEN_72136 : _GEN_72096; // @[FanCtrl.scala 376:33]
  wire [1:0] _GEN_72177 = r_valid_1 ? _GEN_72137 : _GEN_72097; // @[FanCtrl.scala 376:33]
  wire [1:0] _GEN_72178 = r_valid_1 ? _GEN_72138 : _GEN_72098; // @[FanCtrl.scala 376:33]
  wire [1:0] _GEN_72179 = r_valid_1 ? _GEN_72139 : _GEN_72099; // @[FanCtrl.scala 376:33]
  wire [1:0] _GEN_72180 = r_valid_1 ? _GEN_72140 : _GEN_72100; // @[FanCtrl.scala 376:33]
  wire [1:0] _GEN_72181 = r_valid_1 ? _GEN_72141 : _GEN_72101; // @[FanCtrl.scala 376:33]
  wire [1:0] _GEN_72182 = r_valid_1 ? _GEN_72142 : _GEN_72102; // @[FanCtrl.scala 376:33]
  wire [1:0] _GEN_72183 = r_valid_1 ? _GEN_72143 : _GEN_72103; // @[FanCtrl.scala 376:33]
  wire [1:0] _GEN_72184 = r_valid_1 ? _GEN_72144 : _GEN_72104; // @[FanCtrl.scala 376:33]
  wire [1:0] _GEN_72185 = r_valid_1 ? _GEN_72145 : _GEN_72105; // @[FanCtrl.scala 376:33]
  wire [1:0] _GEN_72186 = r_valid_1 ? _GEN_72146 : _GEN_72106; // @[FanCtrl.scala 376:33]
  wire [1:0] _GEN_72187 = r_valid_1 ? _GEN_72147 : _GEN_72107; // @[FanCtrl.scala 376:33]
  wire [1:0] _GEN_72188 = r_valid_1 ? _GEN_72148 : _GEN_72108; // @[FanCtrl.scala 376:33]
  wire [1:0] _GEN_72189 = r_valid_1 ? _GEN_72149 : _GEN_72109; // @[FanCtrl.scala 376:33]
  wire [1:0] _GEN_72190 = r_valid_1 ? _GEN_72150 : _GEN_72110; // @[FanCtrl.scala 376:33]
  wire [1:0] _GEN_72191 = r_valid_1 ? _GEN_72151 : _GEN_72111; // @[FanCtrl.scala 376:33]
  wire [1:0] _GEN_72192 = r_valid_1 ? _GEN_72152 : _GEN_72112; // @[FanCtrl.scala 376:33]
  wire [1:0] _GEN_72193 = r_valid_1 ? _GEN_72153 : _GEN_72113; // @[FanCtrl.scala 376:33]
  wire [1:0] _GEN_72194 = r_valid_1 ? _GEN_72154 : _GEN_72114; // @[FanCtrl.scala 376:33]
  wire [1:0] _GEN_72259 = 4'h0 == _T_361 ? 2'h1 : _GEN_72175; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_72260 = 4'h1 == _T_361 ? 2'h1 : _GEN_72176; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_72261 = 4'h2 == _T_361 ? 2'h1 : _GEN_72177; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_72262 = 4'h3 == _T_361 ? 2'h1 : _GEN_72178; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_72263 = 4'h4 == _T_361 ? 2'h1 : _GEN_72179; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_72264 = 4'h5 == _T_361 ? 2'h1 : _GEN_72180; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_72265 = 4'h6 == _T_361 ? 2'h1 : _GEN_72181; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_72266 = 4'h7 == _T_361 ? 2'h1 : _GEN_72182; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_72267 = 4'h8 == _T_361 ? 2'h1 : _GEN_72183; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_72268 = 4'h9 == _T_361 ? 2'h1 : _GEN_72184; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_72269 = 4'ha == _T_361 ? 2'h1 : _GEN_72185; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_72270 = 4'hb == _T_361 ? 2'h1 : _GEN_72186; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_72271 = 4'hc == _T_361 ? 2'h1 : _GEN_72187; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_72272 = 4'hd == _T_361 ? 2'h1 : _GEN_72188; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_72273 = 4'he == _T_361 ? 2'h1 : _GEN_72189; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_72274 = 4'hf == _T_361 ? 2'h1 : _GEN_72190; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_72275 = 5'h10 == _GEN_94110 ? 2'h1 : _GEN_72191; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_72276 = 5'h11 == _GEN_94110 ? 2'h1 : _GEN_72192; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_72277 = 5'h12 == _GEN_94110 ? 2'h1 : _GEN_72193; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_72278 = 5'h13 == _GEN_94110 ? 2'h1 : _GEN_72194; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_72279 = 4'h0 == _T_361 ? 2'h0 : _GEN_72175; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_72280 = 4'h1 == _T_361 ? 2'h0 : _GEN_72176; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_72281 = 4'h2 == _T_361 ? 2'h0 : _GEN_72177; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_72282 = 4'h3 == _T_361 ? 2'h0 : _GEN_72178; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_72283 = 4'h4 == _T_361 ? 2'h0 : _GEN_72179; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_72284 = 4'h5 == _T_361 ? 2'h0 : _GEN_72180; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_72285 = 4'h6 == _T_361 ? 2'h0 : _GEN_72181; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_72286 = 4'h7 == _T_361 ? 2'h0 : _GEN_72182; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_72287 = 4'h8 == _T_361 ? 2'h0 : _GEN_72183; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_72288 = 4'h9 == _T_361 ? 2'h0 : _GEN_72184; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_72289 = 4'ha == _T_361 ? 2'h0 : _GEN_72185; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_72290 = 4'hb == _T_361 ? 2'h0 : _GEN_72186; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_72291 = 4'hc == _T_361 ? 2'h0 : _GEN_72187; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_72292 = 4'hd == _T_361 ? 2'h0 : _GEN_72188; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_72293 = 4'he == _T_361 ? 2'h0 : _GEN_72189; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_72294 = 4'hf == _T_361 ? 2'h0 : _GEN_72190; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_72295 = 5'h10 == _GEN_94110 ? 2'h0 : _GEN_72191; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_72296 = 5'h11 == _GEN_94110 ? 2'h0 : _GEN_72192; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_72297 = 5'h12 == _GEN_94110 ? 2'h0 : _GEN_72193; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_72298 = 5'h13 == _GEN_94110 ? 2'h0 : _GEN_72194; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_72299 = _T_6909 ? _GEN_72259 : _GEN_72279; // @[FanCtrl.scala 390:64]
  wire [1:0] _GEN_72300 = _T_6909 ? _GEN_72260 : _GEN_72280; // @[FanCtrl.scala 390:64]
  wire [1:0] _GEN_72301 = _T_6909 ? _GEN_72261 : _GEN_72281; // @[FanCtrl.scala 390:64]
  wire [1:0] _GEN_72302 = _T_6909 ? _GEN_72262 : _GEN_72282; // @[FanCtrl.scala 390:64]
  wire [1:0] _GEN_72303 = _T_6909 ? _GEN_72263 : _GEN_72283; // @[FanCtrl.scala 390:64]
  wire [1:0] _GEN_72304 = _T_6909 ? _GEN_72264 : _GEN_72284; // @[FanCtrl.scala 390:64]
  wire [1:0] _GEN_72305 = _T_6909 ? _GEN_72265 : _GEN_72285; // @[FanCtrl.scala 390:64]
  wire [1:0] _GEN_72306 = _T_6909 ? _GEN_72266 : _GEN_72286; // @[FanCtrl.scala 390:64]
  wire [1:0] _GEN_72307 = _T_6909 ? _GEN_72267 : _GEN_72287; // @[FanCtrl.scala 390:64]
  wire [1:0] _GEN_72308 = _T_6909 ? _GEN_72268 : _GEN_72288; // @[FanCtrl.scala 390:64]
  wire [1:0] _GEN_72309 = _T_6909 ? _GEN_72269 : _GEN_72289; // @[FanCtrl.scala 390:64]
  wire [1:0] _GEN_72310 = _T_6909 ? _GEN_72270 : _GEN_72290; // @[FanCtrl.scala 390:64]
  wire [1:0] _GEN_72311 = _T_6909 ? _GEN_72271 : _GEN_72291; // @[FanCtrl.scala 390:64]
  wire [1:0] _GEN_72312 = _T_6909 ? _GEN_72272 : _GEN_72292; // @[FanCtrl.scala 390:64]
  wire [1:0] _GEN_72313 = _T_6909 ? _GEN_72273 : _GEN_72293; // @[FanCtrl.scala 390:64]
  wire [1:0] _GEN_72314 = _T_6909 ? _GEN_72274 : _GEN_72294; // @[FanCtrl.scala 390:64]
  wire [1:0] _GEN_72315 = _T_6909 ? _GEN_72275 : _GEN_72295; // @[FanCtrl.scala 390:64]
  wire [1:0] _GEN_72316 = _T_6909 ? _GEN_72276 : _GEN_72296; // @[FanCtrl.scala 390:64]
  wire [1:0] _GEN_72317 = _T_6909 ? _GEN_72277 : _GEN_72297; // @[FanCtrl.scala 390:64]
  wire [1:0] _GEN_72318 = _T_6909 ? _GEN_72278 : _GEN_72298; // @[FanCtrl.scala 390:64]
  wire  _T_7144 = _T_6966 & _T_6802; // @[FanCtrl.scala 417:67]
  wire  _T_7154 = _T_7144 & _T_6812; // @[FanCtrl.scala 418:66]
  wire  _T_7164 = _T_7154 & _T_6822; // @[FanCtrl.scala 419:66]
  wire [2:0] _GEN_73516 = _T_7017 ? 3'h3 : 3'h0; // @[FanCtrl.scala 432:71]
  wire [2:0] _GEN_73547 = _T_6854 ? 3'h4 : _GEN_73516; // @[FanCtrl.scala 426:72]
  wire [2:0] _GEN_73578 = _T_7164 ? 3'h5 : _GEN_73547; // @[FanCtrl.scala 420:67]
  wire [2:0] _GEN_73702 = r_valid_1 ? _GEN_73578 : 3'h0; // @[FanCtrl.scala 408:33]
  wire [1:0] _GEN_74015 = r_valid_1 ? _GEN_72299 : _GEN_72279; // @[FanCtrl.scala 459:33]
  wire [1:0] _GEN_74016 = r_valid_1 ? _GEN_72300 : _GEN_72280; // @[FanCtrl.scala 459:33]
  wire [1:0] _GEN_74017 = r_valid_1 ? _GEN_72301 : _GEN_72281; // @[FanCtrl.scala 459:33]
  wire [1:0] _GEN_74018 = r_valid_1 ? _GEN_72302 : _GEN_72282; // @[FanCtrl.scala 459:33]
  wire [1:0] _GEN_74019 = r_valid_1 ? _GEN_72303 : _GEN_72283; // @[FanCtrl.scala 459:33]
  wire [1:0] _GEN_74020 = r_valid_1 ? _GEN_72304 : _GEN_72284; // @[FanCtrl.scala 459:33]
  wire [1:0] _GEN_74021 = r_valid_1 ? _GEN_72305 : _GEN_72285; // @[FanCtrl.scala 459:33]
  wire [1:0] _GEN_74022 = r_valid_1 ? _GEN_72306 : _GEN_72286; // @[FanCtrl.scala 459:33]
  wire [1:0] _GEN_74023 = r_valid_1 ? _GEN_72307 : _GEN_72287; // @[FanCtrl.scala 459:33]
  wire [1:0] _GEN_74024 = r_valid_1 ? _GEN_72308 : _GEN_72288; // @[FanCtrl.scala 459:33]
  wire [1:0] _GEN_74025 = r_valid_1 ? _GEN_72309 : _GEN_72289; // @[FanCtrl.scala 459:33]
  wire [1:0] _GEN_74026 = r_valid_1 ? _GEN_72310 : _GEN_72290; // @[FanCtrl.scala 459:33]
  wire [1:0] _GEN_74027 = r_valid_1 ? _GEN_72311 : _GEN_72291; // @[FanCtrl.scala 459:33]
  wire [1:0] _GEN_74028 = r_valid_1 ? _GEN_72312 : _GEN_72292; // @[FanCtrl.scala 459:33]
  wire [1:0] _GEN_74029 = r_valid_1 ? _GEN_72313 : _GEN_72293; // @[FanCtrl.scala 459:33]
  wire [1:0] _GEN_74030 = r_valid_1 ? _GEN_72314 : _GEN_72294; // @[FanCtrl.scala 459:33]
  wire [1:0] _GEN_74031 = r_valid_1 ? _GEN_72315 : _GEN_72295; // @[FanCtrl.scala 459:33]
  wire [1:0] _GEN_74032 = r_valid_1 ? _GEN_72316 : _GEN_72296; // @[FanCtrl.scala 459:33]
  wire [1:0] _GEN_74033 = r_valid_1 ? _GEN_72317 : _GEN_72297; // @[FanCtrl.scala 459:33]
  wire [1:0] _GEN_74034 = r_valid_1 ? _GEN_72318 : _GEN_72298; // @[FanCtrl.scala 459:33]
  wire [5:0] _T_7281 = 4'h8 * 2'h3; // @[FanCtrl.scala 276:23]
  wire [5:0] _T_7283 = _T_7281 + 6'h3; // @[FanCtrl.scala 276:29]
  wire [5:0] _T_7287 = _T_7281 + 6'h4; // @[FanCtrl.scala 276:56]
  wire [4:0] _GEN_74284 = 5'h3 == _T_7283[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_74285 = 5'h4 == _T_7283[4:0] ? w_vn_4 : _GEN_74284; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_74286 = 5'h5 == _T_7283[4:0] ? 5'h0 : _GEN_74285; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_74287 = 5'h6 == _T_7283[4:0] ? 5'h0 : _GEN_74286; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_74288 = 5'h7 == _T_7283[4:0] ? w_vn_7 : _GEN_74287; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_74289 = 5'h8 == _T_7283[4:0] ? w_vn_8 : _GEN_74288; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_74290 = 5'h9 == _T_7283[4:0] ? 5'h0 : _GEN_74289; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_74291 = 5'ha == _T_7283[4:0] ? 5'h0 : _GEN_74290; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_74292 = 5'hb == _T_7283[4:0] ? w_vn_11 : _GEN_74291; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_74293 = 5'hc == _T_7283[4:0] ? w_vn_12 : _GEN_74292; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_74294 = 5'hd == _T_7283[4:0] ? w_vn_13 : _GEN_74293; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_74295 = 5'he == _T_7283[4:0] ? 5'h0 : _GEN_74294; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_74296 = 5'hf == _T_7283[4:0] ? w_vn_15 : _GEN_74295; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_74297 = 5'h10 == _T_7283[4:0] ? w_vn_16 : _GEN_74296; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_74298 = 5'h11 == _T_7283[4:0] ? 5'h0 : _GEN_74297; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_74299 = 5'h12 == _T_7283[4:0] ? w_vn_18 : _GEN_74298; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_74300 = 5'h13 == _T_7283[4:0] ? 5'h0 : _GEN_74299; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_74301 = 5'h14 == _T_7283[4:0] ? 5'h0 : _GEN_74300; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_74302 = 5'h15 == _T_7283[4:0] ? 5'h0 : _GEN_74301; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_74303 = 5'h16 == _T_7283[4:0] ? 5'h0 : _GEN_74302; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_74304 = 5'h17 == _T_7283[4:0] ? w_vn_23 : _GEN_74303; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_74305 = 5'h18 == _T_7283[4:0] ? w_vn_24 : _GEN_74304; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_74306 = 5'h19 == _T_7283[4:0] ? 5'h0 : _GEN_74305; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_74307 = 5'h1a == _T_7283[4:0] ? 5'h0 : _GEN_74306; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_74308 = 5'h1b == _T_7283[4:0] ? 5'h0 : _GEN_74307; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_74309 = 5'h1c == _T_7283[4:0] ? 5'h0 : _GEN_74308; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_74310 = 5'h1d == _T_7283[4:0] ? 5'h0 : _GEN_74309; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_74311 = 5'h1e == _T_7283[4:0] ? 5'h0 : _GEN_74310; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_74312 = 5'h1f == _T_7283[4:0] ? 5'h0 : _GEN_74311; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_74316 = 5'h3 == _T_7287[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_74317 = 5'h4 == _T_7287[4:0] ? w_vn_4 : _GEN_74316; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_74318 = 5'h5 == _T_7287[4:0] ? 5'h0 : _GEN_74317; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_74319 = 5'h6 == _T_7287[4:0] ? 5'h0 : _GEN_74318; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_74320 = 5'h7 == _T_7287[4:0] ? w_vn_7 : _GEN_74319; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_74321 = 5'h8 == _T_7287[4:0] ? w_vn_8 : _GEN_74320; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_74322 = 5'h9 == _T_7287[4:0] ? 5'h0 : _GEN_74321; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_74323 = 5'ha == _T_7287[4:0] ? 5'h0 : _GEN_74322; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_74324 = 5'hb == _T_7287[4:0] ? w_vn_11 : _GEN_74323; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_74325 = 5'hc == _T_7287[4:0] ? w_vn_12 : _GEN_74324; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_74326 = 5'hd == _T_7287[4:0] ? w_vn_13 : _GEN_74325; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_74327 = 5'he == _T_7287[4:0] ? 5'h0 : _GEN_74326; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_74328 = 5'hf == _T_7287[4:0] ? w_vn_15 : _GEN_74327; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_74329 = 5'h10 == _T_7287[4:0] ? w_vn_16 : _GEN_74328; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_74330 = 5'h11 == _T_7287[4:0] ? 5'h0 : _GEN_74329; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_74331 = 5'h12 == _T_7287[4:0] ? w_vn_18 : _GEN_74330; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_74332 = 5'h13 == _T_7287[4:0] ? 5'h0 : _GEN_74331; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_74333 = 5'h14 == _T_7287[4:0] ? 5'h0 : _GEN_74332; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_74334 = 5'h15 == _T_7287[4:0] ? 5'h0 : _GEN_74333; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_74335 = 5'h16 == _T_7287[4:0] ? 5'h0 : _GEN_74334; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_74336 = 5'h17 == _T_7287[4:0] ? w_vn_23 : _GEN_74335; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_74337 = 5'h18 == _T_7287[4:0] ? w_vn_24 : _GEN_74336; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_74338 = 5'h19 == _T_7287[4:0] ? 5'h0 : _GEN_74337; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_74339 = 5'h1a == _T_7287[4:0] ? 5'h0 : _GEN_74338; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_74340 = 5'h1b == _T_7287[4:0] ? 5'h0 : _GEN_74339; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_74341 = 5'h1c == _T_7287[4:0] ? 5'h0 : _GEN_74340; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_74342 = 5'h1d == _T_7287[4:0] ? 5'h0 : _GEN_74341; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_74343 = 5'h1e == _T_7287[4:0] ? 5'h0 : _GEN_74342; // @[FanCtrl.scala 276:{37,37}]
  wire [4:0] _GEN_74344 = 5'h1f == _T_7287[4:0] ? 5'h0 : _GEN_74343; // @[FanCtrl.scala 276:{37,37}]
  wire  _T_7289 = _GEN_74312 == _GEN_74344; // @[FanCtrl.scala 276:37]
  wire [5:0] _T_7296 = _T_7281 + 6'h1; // @[FanCtrl.scala 282:30]
  wire [5:0] _T_7300 = _T_7281 + 6'h2; // @[FanCtrl.scala 282:56]
  wire [4:0] _GEN_74441 = 5'h3 == _T_7296[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_74442 = 5'h4 == _T_7296[4:0] ? w_vn_4 : _GEN_74441; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_74443 = 5'h5 == _T_7296[4:0] ? 5'h0 : _GEN_74442; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_74444 = 5'h6 == _T_7296[4:0] ? 5'h0 : _GEN_74443; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_74445 = 5'h7 == _T_7296[4:0] ? w_vn_7 : _GEN_74444; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_74446 = 5'h8 == _T_7296[4:0] ? w_vn_8 : _GEN_74445; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_74447 = 5'h9 == _T_7296[4:0] ? 5'h0 : _GEN_74446; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_74448 = 5'ha == _T_7296[4:0] ? 5'h0 : _GEN_74447; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_74449 = 5'hb == _T_7296[4:0] ? w_vn_11 : _GEN_74448; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_74450 = 5'hc == _T_7296[4:0] ? w_vn_12 : _GEN_74449; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_74451 = 5'hd == _T_7296[4:0] ? w_vn_13 : _GEN_74450; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_74452 = 5'he == _T_7296[4:0] ? 5'h0 : _GEN_74451; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_74453 = 5'hf == _T_7296[4:0] ? w_vn_15 : _GEN_74452; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_74454 = 5'h10 == _T_7296[4:0] ? w_vn_16 : _GEN_74453; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_74455 = 5'h11 == _T_7296[4:0] ? 5'h0 : _GEN_74454; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_74456 = 5'h12 == _T_7296[4:0] ? w_vn_18 : _GEN_74455; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_74457 = 5'h13 == _T_7296[4:0] ? 5'h0 : _GEN_74456; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_74458 = 5'h14 == _T_7296[4:0] ? 5'h0 : _GEN_74457; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_74459 = 5'h15 == _T_7296[4:0] ? 5'h0 : _GEN_74458; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_74460 = 5'h16 == _T_7296[4:0] ? 5'h0 : _GEN_74459; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_74461 = 5'h17 == _T_7296[4:0] ? w_vn_23 : _GEN_74460; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_74462 = 5'h18 == _T_7296[4:0] ? w_vn_24 : _GEN_74461; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_74463 = 5'h19 == _T_7296[4:0] ? 5'h0 : _GEN_74462; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_74464 = 5'h1a == _T_7296[4:0] ? 5'h0 : _GEN_74463; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_74465 = 5'h1b == _T_7296[4:0] ? 5'h0 : _GEN_74464; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_74466 = 5'h1c == _T_7296[4:0] ? 5'h0 : _GEN_74465; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_74467 = 5'h1d == _T_7296[4:0] ? 5'h0 : _GEN_74466; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_74468 = 5'h1e == _T_7296[4:0] ? 5'h0 : _GEN_74467; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_74469 = 5'h1f == _T_7296[4:0] ? 5'h0 : _GEN_74468; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_74473 = 5'h3 == _T_7300[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_74474 = 5'h4 == _T_7300[4:0] ? w_vn_4 : _GEN_74473; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_74475 = 5'h5 == _T_7300[4:0] ? 5'h0 : _GEN_74474; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_74476 = 5'h6 == _T_7300[4:0] ? 5'h0 : _GEN_74475; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_74477 = 5'h7 == _T_7300[4:0] ? w_vn_7 : _GEN_74476; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_74478 = 5'h8 == _T_7300[4:0] ? w_vn_8 : _GEN_74477; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_74479 = 5'h9 == _T_7300[4:0] ? 5'h0 : _GEN_74478; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_74480 = 5'ha == _T_7300[4:0] ? 5'h0 : _GEN_74479; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_74481 = 5'hb == _T_7300[4:0] ? w_vn_11 : _GEN_74480; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_74482 = 5'hc == _T_7300[4:0] ? w_vn_12 : _GEN_74481; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_74483 = 5'hd == _T_7300[4:0] ? w_vn_13 : _GEN_74482; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_74484 = 5'he == _T_7300[4:0] ? 5'h0 : _GEN_74483; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_74485 = 5'hf == _T_7300[4:0] ? w_vn_15 : _GEN_74484; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_74486 = 5'h10 == _T_7300[4:0] ? w_vn_16 : _GEN_74485; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_74487 = 5'h11 == _T_7300[4:0] ? 5'h0 : _GEN_74486; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_74488 = 5'h12 == _T_7300[4:0] ? w_vn_18 : _GEN_74487; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_74489 = 5'h13 == _T_7300[4:0] ? 5'h0 : _GEN_74488; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_74490 = 5'h14 == _T_7300[4:0] ? 5'h0 : _GEN_74489; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_74491 = 5'h15 == _T_7300[4:0] ? 5'h0 : _GEN_74490; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_74492 = 5'h16 == _T_7300[4:0] ? 5'h0 : _GEN_74491; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_74493 = 5'h17 == _T_7300[4:0] ? w_vn_23 : _GEN_74492; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_74494 = 5'h18 == _T_7300[4:0] ? w_vn_24 : _GEN_74493; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_74495 = 5'h19 == _T_7300[4:0] ? 5'h0 : _GEN_74494; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_74496 = 5'h1a == _T_7300[4:0] ? 5'h0 : _GEN_74495; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_74497 = 5'h1b == _T_7300[4:0] ? 5'h0 : _GEN_74496; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_74498 = 5'h1c == _T_7300[4:0] ? 5'h0 : _GEN_74497; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_74499 = 5'h1d == _T_7300[4:0] ? 5'h0 : _GEN_74498; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_74500 = 5'h1e == _T_7300[4:0] ? 5'h0 : _GEN_74499; // @[FanCtrl.scala 282:{37,37}]
  wire [4:0] _GEN_74501 = 5'h1f == _T_7300[4:0] ? 5'h0 : _GEN_74500; // @[FanCtrl.scala 282:{37,37}]
  wire  _T_7302 = _GEN_74469 == _GEN_74501; // @[FanCtrl.scala 282:37]
  wire [5:0] _T_7305 = _T_7281 + 6'h5; // @[FanCtrl.scala 283:29]
  wire [5:0] _T_7309 = _T_7281 + 6'h6; // @[FanCtrl.scala 283:56]
  wire [4:0] _GEN_74505 = 5'h3 == _T_7305[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_74506 = 5'h4 == _T_7305[4:0] ? w_vn_4 : _GEN_74505; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_74507 = 5'h5 == _T_7305[4:0] ? 5'h0 : _GEN_74506; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_74508 = 5'h6 == _T_7305[4:0] ? 5'h0 : _GEN_74507; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_74509 = 5'h7 == _T_7305[4:0] ? w_vn_7 : _GEN_74508; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_74510 = 5'h8 == _T_7305[4:0] ? w_vn_8 : _GEN_74509; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_74511 = 5'h9 == _T_7305[4:0] ? 5'h0 : _GEN_74510; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_74512 = 5'ha == _T_7305[4:0] ? 5'h0 : _GEN_74511; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_74513 = 5'hb == _T_7305[4:0] ? w_vn_11 : _GEN_74512; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_74514 = 5'hc == _T_7305[4:0] ? w_vn_12 : _GEN_74513; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_74515 = 5'hd == _T_7305[4:0] ? w_vn_13 : _GEN_74514; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_74516 = 5'he == _T_7305[4:0] ? 5'h0 : _GEN_74515; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_74517 = 5'hf == _T_7305[4:0] ? w_vn_15 : _GEN_74516; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_74518 = 5'h10 == _T_7305[4:0] ? w_vn_16 : _GEN_74517; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_74519 = 5'h11 == _T_7305[4:0] ? 5'h0 : _GEN_74518; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_74520 = 5'h12 == _T_7305[4:0] ? w_vn_18 : _GEN_74519; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_74521 = 5'h13 == _T_7305[4:0] ? 5'h0 : _GEN_74520; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_74522 = 5'h14 == _T_7305[4:0] ? 5'h0 : _GEN_74521; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_74523 = 5'h15 == _T_7305[4:0] ? 5'h0 : _GEN_74522; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_74524 = 5'h16 == _T_7305[4:0] ? 5'h0 : _GEN_74523; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_74525 = 5'h17 == _T_7305[4:0] ? w_vn_23 : _GEN_74524; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_74526 = 5'h18 == _T_7305[4:0] ? w_vn_24 : _GEN_74525; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_74527 = 5'h19 == _T_7305[4:0] ? 5'h0 : _GEN_74526; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_74528 = 5'h1a == _T_7305[4:0] ? 5'h0 : _GEN_74527; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_74529 = 5'h1b == _T_7305[4:0] ? 5'h0 : _GEN_74528; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_74530 = 5'h1c == _T_7305[4:0] ? 5'h0 : _GEN_74529; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_74531 = 5'h1d == _T_7305[4:0] ? 5'h0 : _GEN_74530; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_74532 = 5'h1e == _T_7305[4:0] ? 5'h0 : _GEN_74531; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_74533 = 5'h1f == _T_7305[4:0] ? 5'h0 : _GEN_74532; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_74537 = 5'h3 == _T_7309[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_74538 = 5'h4 == _T_7309[4:0] ? w_vn_4 : _GEN_74537; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_74539 = 5'h5 == _T_7309[4:0] ? 5'h0 : _GEN_74538; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_74540 = 5'h6 == _T_7309[4:0] ? 5'h0 : _GEN_74539; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_74541 = 5'h7 == _T_7309[4:0] ? w_vn_7 : _GEN_74540; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_74542 = 5'h8 == _T_7309[4:0] ? w_vn_8 : _GEN_74541; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_74543 = 5'h9 == _T_7309[4:0] ? 5'h0 : _GEN_74542; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_74544 = 5'ha == _T_7309[4:0] ? 5'h0 : _GEN_74543; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_74545 = 5'hb == _T_7309[4:0] ? w_vn_11 : _GEN_74544; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_74546 = 5'hc == _T_7309[4:0] ? w_vn_12 : _GEN_74545; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_74547 = 5'hd == _T_7309[4:0] ? w_vn_13 : _GEN_74546; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_74548 = 5'he == _T_7309[4:0] ? 5'h0 : _GEN_74547; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_74549 = 5'hf == _T_7309[4:0] ? w_vn_15 : _GEN_74548; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_74550 = 5'h10 == _T_7309[4:0] ? w_vn_16 : _GEN_74549; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_74551 = 5'h11 == _T_7309[4:0] ? 5'h0 : _GEN_74550; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_74552 = 5'h12 == _T_7309[4:0] ? w_vn_18 : _GEN_74551; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_74553 = 5'h13 == _T_7309[4:0] ? 5'h0 : _GEN_74552; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_74554 = 5'h14 == _T_7309[4:0] ? 5'h0 : _GEN_74553; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_74555 = 5'h15 == _T_7309[4:0] ? 5'h0 : _GEN_74554; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_74556 = 5'h16 == _T_7309[4:0] ? 5'h0 : _GEN_74555; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_74557 = 5'h17 == _T_7309[4:0] ? w_vn_23 : _GEN_74556; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_74558 = 5'h18 == _T_7309[4:0] ? w_vn_24 : _GEN_74557; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_74559 = 5'h19 == _T_7309[4:0] ? 5'h0 : _GEN_74558; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_74560 = 5'h1a == _T_7309[4:0] ? 5'h0 : _GEN_74559; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_74561 = 5'h1b == _T_7309[4:0] ? 5'h0 : _GEN_74560; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_74562 = 5'h1c == _T_7309[4:0] ? 5'h0 : _GEN_74561; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_74563 = 5'h1d == _T_7309[4:0] ? 5'h0 : _GEN_74562; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_74564 = 5'h1e == _T_7309[4:0] ? 5'h0 : _GEN_74563; // @[FanCtrl.scala 283:{37,37}]
  wire [4:0] _GEN_74565 = 5'h1f == _T_7309[4:0] ? 5'h0 : _GEN_74564; // @[FanCtrl.scala 283:{37,37}]
  wire  _T_7311 = _GEN_74533 == _GEN_74565; // @[FanCtrl.scala 283:37]
  wire  _T_7312 = _GEN_74469 == _GEN_74501 & _T_7311; // @[FanCtrl.scala 282:64]
  wire  _T_7331 = _GEN_74501 != _GEN_74344; // @[FanCtrl.scala 285:36]
  wire  _T_7341 = _GEN_74533 != _GEN_74312; // @[FanCtrl.scala 286:37]
  wire  _GEN_75384 = r_valid_1 & _T_7289; // @[FanCtrl.scala 274:32]
  wire  _T_7412 = _GEN_74312 == _GEN_74469; // @[FanCtrl.scala 313:39]
  wire  _T_7428 = _GEN_74344 == _GEN_74565; // @[FanCtrl.scala 325:39]
  wire [3:0] _T_7440 = 2'h3 * 2'h2; // @[FanCtrl.scala 338:28]
  wire [4:0] _T_7441 = {{1'd0}, _T_7440}; // @[FanCtrl.scala 338:35]
  wire [1:0] _GEN_75809 = 4'h0 == _T_7441[3:0] ? 2'h0 : _GEN_74015; // @[FanCtrl.scala 338:{42,42}]
  wire [1:0] _GEN_75810 = 4'h1 == _T_7441[3:0] ? 2'h0 : _GEN_74016; // @[FanCtrl.scala 338:{42,42}]
  wire [1:0] _GEN_75811 = 4'h2 == _T_7441[3:0] ? 2'h0 : _GEN_74017; // @[FanCtrl.scala 338:{42,42}]
  wire [1:0] _GEN_75812 = 4'h3 == _T_7441[3:0] ? 2'h0 : _GEN_74018; // @[FanCtrl.scala 338:{42,42}]
  wire [1:0] _GEN_75813 = 4'h4 == _T_7441[3:0] ? 2'h0 : _GEN_74019; // @[FanCtrl.scala 338:{42,42}]
  wire [1:0] _GEN_75814 = 4'h5 == _T_7441[3:0] ? 2'h0 : _GEN_74020; // @[FanCtrl.scala 338:{42,42}]
  wire [1:0] _GEN_75815 = 4'h6 == _T_7441[3:0] ? 2'h0 : _GEN_74021; // @[FanCtrl.scala 338:{42,42}]
  wire [1:0] _GEN_75816 = 4'h7 == _T_7441[3:0] ? 2'h0 : _GEN_74022; // @[FanCtrl.scala 338:{42,42}]
  wire [1:0] _GEN_75817 = 4'h8 == _T_7441[3:0] ? 2'h0 : _GEN_74023; // @[FanCtrl.scala 338:{42,42}]
  wire [1:0] _GEN_75818 = 4'h9 == _T_7441[3:0] ? 2'h0 : _GEN_74024; // @[FanCtrl.scala 338:{42,42}]
  wire [1:0] _GEN_75819 = 4'ha == _T_7441[3:0] ? 2'h0 : _GEN_74025; // @[FanCtrl.scala 338:{42,42}]
  wire [1:0] _GEN_75820 = 4'hb == _T_7441[3:0] ? 2'h0 : _GEN_74026; // @[FanCtrl.scala 338:{42,42}]
  wire [1:0] _GEN_75821 = 4'hc == _T_7441[3:0] ? 2'h0 : _GEN_74027; // @[FanCtrl.scala 338:{42,42}]
  wire [1:0] _GEN_75822 = 4'hd == _T_7441[3:0] ? 2'h0 : _GEN_74028; // @[FanCtrl.scala 338:{42,42}]
  wire [1:0] _GEN_75823 = 4'he == _T_7441[3:0] ? 2'h0 : _GEN_74029; // @[FanCtrl.scala 338:{42,42}]
  wire [1:0] _GEN_75824 = 4'hf == _T_7441[3:0] ? 2'h0 : _GEN_74030; // @[FanCtrl.scala 338:{42,42}]
  wire [4:0] _GEN_97814 = {{1'd0}, _T_7441[3:0]}; // @[FanCtrl.scala 338:{42,42}]
  wire [1:0] _GEN_75825 = 5'h10 == _GEN_97814 ? 2'h0 : _GEN_74031; // @[FanCtrl.scala 338:{42,42}]
  wire [1:0] _GEN_75826 = 5'h11 == _GEN_97814 ? 2'h0 : _GEN_74032; // @[FanCtrl.scala 338:{42,42}]
  wire [1:0] _GEN_75827 = 5'h12 == _GEN_97814 ? 2'h0 : _GEN_74033; // @[FanCtrl.scala 338:{42,42}]
  wire [1:0] _GEN_75828 = 5'h13 == _GEN_97814 ? 2'h0 : _GEN_74034; // @[FanCtrl.scala 338:{42,42}]
  wire [5:0] _T_7482 = _T_7281 - 6'h1; // @[FanCtrl.scala 349:58]
  wire [4:0] _GEN_76149 = 5'h3 == _T_7482[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_76150 = 5'h4 == _T_7482[4:0] ? w_vn_4 : _GEN_76149; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_76151 = 5'h5 == _T_7482[4:0] ? 5'h0 : _GEN_76150; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_76152 = 5'h6 == _T_7482[4:0] ? 5'h0 : _GEN_76151; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_76153 = 5'h7 == _T_7482[4:0] ? w_vn_7 : _GEN_76152; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_76154 = 5'h8 == _T_7482[4:0] ? w_vn_8 : _GEN_76153; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_76155 = 5'h9 == _T_7482[4:0] ? 5'h0 : _GEN_76154; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_76156 = 5'ha == _T_7482[4:0] ? 5'h0 : _GEN_76155; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_76157 = 5'hb == _T_7482[4:0] ? w_vn_11 : _GEN_76156; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_76158 = 5'hc == _T_7482[4:0] ? w_vn_12 : _GEN_76157; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_76159 = 5'hd == _T_7482[4:0] ? w_vn_13 : _GEN_76158; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_76160 = 5'he == _T_7482[4:0] ? 5'h0 : _GEN_76159; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_76161 = 5'hf == _T_7482[4:0] ? w_vn_15 : _GEN_76160; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_76162 = 5'h10 == _T_7482[4:0] ? w_vn_16 : _GEN_76161; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_76163 = 5'h11 == _T_7482[4:0] ? 5'h0 : _GEN_76162; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_76164 = 5'h12 == _T_7482[4:0] ? w_vn_18 : _GEN_76163; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_76165 = 5'h13 == _T_7482[4:0] ? 5'h0 : _GEN_76164; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_76166 = 5'h14 == _T_7482[4:0] ? 5'h0 : _GEN_76165; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_76167 = 5'h15 == _T_7482[4:0] ? 5'h0 : _GEN_76166; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_76168 = 5'h16 == _T_7482[4:0] ? 5'h0 : _GEN_76167; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_76169 = 5'h17 == _T_7482[4:0] ? w_vn_23 : _GEN_76168; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_76170 = 5'h18 == _T_7482[4:0] ? w_vn_24 : _GEN_76169; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_76171 = 5'h19 == _T_7482[4:0] ? 5'h0 : _GEN_76170; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_76172 = 5'h1a == _T_7482[4:0] ? 5'h0 : _GEN_76171; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_76173 = 5'h1b == _T_7482[4:0] ? 5'h0 : _GEN_76172; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_76174 = 5'h1c == _T_7482[4:0] ? 5'h0 : _GEN_76173; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_76175 = 5'h1d == _T_7482[4:0] ? 5'h0 : _GEN_76174; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_76176 = 5'h1e == _T_7482[4:0] ? 5'h0 : _GEN_76175; // @[FanCtrl.scala 349:{39,39}]
  wire [4:0] _GEN_76177 = 5'h1f == _T_7482[4:0] ? 5'h0 : _GEN_76176; // @[FanCtrl.scala 349:{39,39}]
  wire  _T_7484 = _GEN_74469 != _GEN_76177; // @[FanCtrl.scala 349:39]
  wire  _T_7485 = _T_7312 & _T_7484; // @[FanCtrl.scala 348:67]
  wire  _T_7495 = _T_7485 & _T_7331; // @[FanCtrl.scala 349:67]
  wire  _T_7505 = _T_7495 & _T_7341; // @[FanCtrl.scala 350:67]
  wire  _T_7526 = _T_7302 & _T_7484; // @[FanCtrl.scala 355:73]
  wire  _T_7535 = _GEN_74344 != _GEN_74501; // @[FanCtrl.scala 357:42]
  wire  _T_7536 = _T_7526 & _T_7535; // @[FanCtrl.scala 356:71]
  wire  _T_7557 = _T_7311 & _T_7341; // @[FanCtrl.scala 361:72]
  wire [6:0] _T_7558 = 5'h18 * 2'h3; // @[FanCtrl.scala 364:33]
  wire [2:0] _GEN_76688 = 5'h0 == _T_7558[4:0] ? 3'h4 : _GEN_477; // @[FanCtrl.scala 364:{40,40}]
  wire [2:0] _GEN_76689 = 5'h1 == _T_7558[4:0] ? 3'h4 : _GEN_3697; // @[FanCtrl.scala 364:{40,40}]
  wire [2:0] _GEN_76690 = 5'h2 == _T_7558[4:0] ? 3'h4 : _GEN_5579; // @[FanCtrl.scala 364:{40,40}]
  wire [2:0] _GEN_76691 = 5'h3 == _T_7558[4:0] ? 3'h4 : _GEN_7461; // @[FanCtrl.scala 364:{40,40}]
  wire [2:0] _GEN_76692 = 5'h4 == _T_7558[4:0] ? 3'h4 : _GEN_9343; // @[FanCtrl.scala 364:{40,40}]
  wire [2:0] _GEN_76693 = 5'h5 == _T_7558[4:0] ? 3'h4 : _GEN_11225; // @[FanCtrl.scala 364:{40,40}]
  wire [2:0] _GEN_76694 = 5'h6 == _T_7558[4:0] ? 3'h4 : _GEN_13107; // @[FanCtrl.scala 364:{40,40}]
  wire [2:0] _GEN_76695 = 5'h7 == _T_7558[4:0] ? 3'h4 : _GEN_14989; // @[FanCtrl.scala 364:{40,40}]
  wire [2:0] _GEN_76696 = 5'h8 == _T_7558[4:0] ? 3'h4 : _GEN_16871; // @[FanCtrl.scala 364:{40,40}]
  wire [2:0] _GEN_76697 = 5'h9 == _T_7558[4:0] ? 3'h4 : _GEN_18753; // @[FanCtrl.scala 364:{40,40}]
  wire [2:0] _GEN_76698 = 5'ha == _T_7558[4:0] ? 3'h4 : _GEN_20635; // @[FanCtrl.scala 364:{40,40}]
  wire [2:0] _GEN_76699 = 5'hb == _T_7558[4:0] ? 3'h4 : _GEN_22517; // @[FanCtrl.scala 364:{40,40}]
  wire [2:0] _GEN_76700 = 5'hc == _T_7558[4:0] ? 3'h4 : _GEN_24399; // @[FanCtrl.scala 364:{40,40}]
  wire [2:0] _GEN_76701 = 5'hd == _T_7558[4:0] ? 3'h4 : _GEN_26281; // @[FanCtrl.scala 364:{40,40}]
  wire [2:0] _GEN_76702 = 5'he == _T_7558[4:0] ? 3'h4 : _GEN_28163; // @[FanCtrl.scala 364:{40,40}]
  wire [2:0] _GEN_76703 = 5'hf == _T_7558[4:0] ? 3'h4 : _GEN_29215; // @[FanCtrl.scala 364:{40,40}]
  wire [2:0] _GEN_76704 = 5'h10 == _T_7558[4:0] ? 3'h4 : _GEN_31232; // @[FanCtrl.scala 364:{40,40}]
  wire [2:0] _GEN_76705 = 5'h11 == _T_7558[4:0] ? 3'h4 : _GEN_37293; // @[FanCtrl.scala 364:{40,40}]
  wire [2:0] _GEN_76706 = 5'h12 == _T_7558[4:0] ? 3'h4 : _GEN_40954; // @[FanCtrl.scala 364:{40,40}]
  wire [2:0] _GEN_76707 = 5'h13 == _T_7558[4:0] ? 3'h4 : _GEN_44615; // @[FanCtrl.scala 364:{40,40}]
  wire [2:0] _GEN_76708 = 5'h14 == _T_7558[4:0] ? 3'h4 : _GEN_48276; // @[FanCtrl.scala 364:{40,40}]
  wire [2:0] _GEN_76709 = 5'h15 == _T_7558[4:0] ? 3'h4 : _GEN_51937; // @[FanCtrl.scala 364:{40,40}]
  wire [2:0] _GEN_76710 = 5'h16 == _T_7558[4:0] ? 3'h4 : _GEN_55598; // @[FanCtrl.scala 364:{40,40}]
  wire [2:0] _GEN_76711 = 5'h17 == _T_7558[4:0] ? 3'h4 : _GEN_57995; // @[FanCtrl.scala 364:{40,40}]
  wire [2:0] _GEN_76712 = 5'h18 == _T_7558[4:0] ? 3'h4 : _GEN_60604; // @[FanCtrl.scala 364:{40,40}]
  wire [2:0] _GEN_76713 = 5'h19 == _T_7558[4:0] ? 3'h4 : _GEN_68765; // @[FanCtrl.scala 364:{40,40}]
  wire [2:0] _GEN_76714 = 5'h1a == _T_7558[4:0] ? 3'h4 : _GEN_73702; // @[FanCtrl.scala 364:{40,40}]
  wire [2:0] _GEN_76715 = 5'h1b == _T_7558[4:0] ? 3'h4 : 3'h0; // @[FanCtrl.scala 364:{40,40}]
  wire [2:0] _GEN_76750 = _T_7557 ? _GEN_76688 : _GEN_477; // @[FanCtrl.scala 362:71]
  wire [2:0] _GEN_76751 = _T_7557 ? _GEN_76689 : _GEN_3697; // @[FanCtrl.scala 362:71]
  wire [2:0] _GEN_76752 = _T_7557 ? _GEN_76690 : _GEN_5579; // @[FanCtrl.scala 362:71]
  wire [2:0] _GEN_76753 = _T_7557 ? _GEN_76691 : _GEN_7461; // @[FanCtrl.scala 362:71]
  wire [2:0] _GEN_76754 = _T_7557 ? _GEN_76692 : _GEN_9343; // @[FanCtrl.scala 362:71]
  wire [2:0] _GEN_76755 = _T_7557 ? _GEN_76693 : _GEN_11225; // @[FanCtrl.scala 362:71]
  wire [2:0] _GEN_76756 = _T_7557 ? _GEN_76694 : _GEN_13107; // @[FanCtrl.scala 362:71]
  wire [2:0] _GEN_76757 = _T_7557 ? _GEN_76695 : _GEN_14989; // @[FanCtrl.scala 362:71]
  wire [2:0] _GEN_76758 = _T_7557 ? _GEN_76696 : _GEN_16871; // @[FanCtrl.scala 362:71]
  wire [2:0] _GEN_76759 = _T_7557 ? _GEN_76697 : _GEN_18753; // @[FanCtrl.scala 362:71]
  wire [2:0] _GEN_76760 = _T_7557 ? _GEN_76698 : _GEN_20635; // @[FanCtrl.scala 362:71]
  wire [2:0] _GEN_76761 = _T_7557 ? _GEN_76699 : _GEN_22517; // @[FanCtrl.scala 362:71]
  wire [2:0] _GEN_76762 = _T_7557 ? _GEN_76700 : _GEN_24399; // @[FanCtrl.scala 362:71]
  wire [2:0] _GEN_76763 = _T_7557 ? _GEN_76701 : _GEN_26281; // @[FanCtrl.scala 362:71]
  wire [2:0] _GEN_76764 = _T_7557 ? _GEN_76702 : _GEN_28163; // @[FanCtrl.scala 362:71]
  wire [2:0] _GEN_76765 = _T_7557 ? _GEN_76703 : _GEN_29215; // @[FanCtrl.scala 362:71]
  wire [2:0] _GEN_76766 = _T_7557 ? _GEN_76704 : _GEN_31232; // @[FanCtrl.scala 362:71]
  wire [2:0] _GEN_76767 = _T_7557 ? _GEN_76705 : _GEN_37293; // @[FanCtrl.scala 362:71]
  wire [2:0] _GEN_76768 = _T_7557 ? _GEN_76706 : _GEN_40954; // @[FanCtrl.scala 362:71]
  wire [2:0] _GEN_76769 = _T_7557 ? _GEN_76707 : _GEN_44615; // @[FanCtrl.scala 362:71]
  wire [2:0] _GEN_76770 = _T_7557 ? _GEN_76708 : _GEN_48276; // @[FanCtrl.scala 362:71]
  wire [2:0] _GEN_76771 = _T_7557 ? _GEN_76709 : _GEN_51937; // @[FanCtrl.scala 362:71]
  wire [2:0] _GEN_76772 = _T_7557 ? _GEN_76710 : _GEN_55598; // @[FanCtrl.scala 362:71]
  wire [2:0] _GEN_76773 = _T_7557 ? _GEN_76711 : _GEN_57995; // @[FanCtrl.scala 362:71]
  wire [2:0] _GEN_76774 = _T_7557 ? _GEN_76712 : _GEN_60604; // @[FanCtrl.scala 362:71]
  wire [2:0] _GEN_76775 = _T_7557 ? _GEN_76713 : _GEN_68765; // @[FanCtrl.scala 362:71]
  wire [2:0] _GEN_76776 = _T_7557 ? _GEN_76714 : _GEN_73702; // @[FanCtrl.scala 362:71]
  wire [2:0] _GEN_76777 = _T_7557 ? _GEN_76715 : 3'h0; // @[FanCtrl.scala 362:71]
  wire [1:0] _GEN_77031 = 4'h0 == _T_7441[3:0] ? 2'h0 : _GEN_75809; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_77032 = 4'h1 == _T_7441[3:0] ? 2'h0 : _GEN_75810; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_77033 = 4'h2 == _T_7441[3:0] ? 2'h0 : _GEN_75811; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_77034 = 4'h3 == _T_7441[3:0] ? 2'h0 : _GEN_75812; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_77035 = 4'h4 == _T_7441[3:0] ? 2'h0 : _GEN_75813; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_77036 = 4'h5 == _T_7441[3:0] ? 2'h0 : _GEN_75814; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_77037 = 4'h6 == _T_7441[3:0] ? 2'h0 : _GEN_75815; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_77038 = 4'h7 == _T_7441[3:0] ? 2'h0 : _GEN_75816; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_77039 = 4'h8 == _T_7441[3:0] ? 2'h0 : _GEN_75817; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_77040 = 4'h9 == _T_7441[3:0] ? 2'h0 : _GEN_75818; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_77041 = 4'ha == _T_7441[3:0] ? 2'h0 : _GEN_75819; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_77042 = 4'hb == _T_7441[3:0] ? 2'h0 : _GEN_75820; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_77043 = 4'hc == _T_7441[3:0] ? 2'h0 : _GEN_75821; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_77044 = 4'hd == _T_7441[3:0] ? 2'h0 : _GEN_75822; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_77045 = 4'he == _T_7441[3:0] ? 2'h0 : _GEN_75823; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_77046 = 4'hf == _T_7441[3:0] ? 2'h0 : _GEN_75824; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_77047 = 5'h10 == _GEN_97814 ? 2'h0 : _GEN_75825; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_77048 = 5'h11 == _GEN_97814 ? 2'h0 : _GEN_75826; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_77049 = 5'h12 == _GEN_97814 ? 2'h0 : _GEN_75827; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_77050 = 5'h13 == _GEN_97814 ? 2'h0 : _GEN_75828; // @[FanCtrl.scala 379:{46,46}]
  wire [1:0] _GEN_77051 = 4'h0 == _T_7441[3:0] ? 2'h1 : _GEN_75809; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_77052 = 4'h1 == _T_7441[3:0] ? 2'h1 : _GEN_75810; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_77053 = 4'h2 == _T_7441[3:0] ? 2'h1 : _GEN_75811; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_77054 = 4'h3 == _T_7441[3:0] ? 2'h1 : _GEN_75812; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_77055 = 4'h4 == _T_7441[3:0] ? 2'h1 : _GEN_75813; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_77056 = 4'h5 == _T_7441[3:0] ? 2'h1 : _GEN_75814; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_77057 = 4'h6 == _T_7441[3:0] ? 2'h1 : _GEN_75815; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_77058 = 4'h7 == _T_7441[3:0] ? 2'h1 : _GEN_75816; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_77059 = 4'h8 == _T_7441[3:0] ? 2'h1 : _GEN_75817; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_77060 = 4'h9 == _T_7441[3:0] ? 2'h1 : _GEN_75818; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_77061 = 4'ha == _T_7441[3:0] ? 2'h1 : _GEN_75819; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_77062 = 4'hb == _T_7441[3:0] ? 2'h1 : _GEN_75820; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_77063 = 4'hc == _T_7441[3:0] ? 2'h1 : _GEN_75821; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_77064 = 4'hd == _T_7441[3:0] ? 2'h1 : _GEN_75822; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_77065 = 4'he == _T_7441[3:0] ? 2'h1 : _GEN_75823; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_77066 = 4'hf == _T_7441[3:0] ? 2'h1 : _GEN_75824; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_77067 = 5'h10 == _GEN_97814 ? 2'h1 : _GEN_75825; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_77068 = 5'h11 == _GEN_97814 ? 2'h1 : _GEN_75826; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_77069 = 5'h12 == _GEN_97814 ? 2'h1 : _GEN_75827; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_77070 = 5'h13 == _GEN_97814 ? 2'h1 : _GEN_75828; // @[FanCtrl.scala 382:{46,46}]
  wire [1:0] _GEN_77071 = _T_7412 ? _GEN_77031 : _GEN_77051; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_77072 = _T_7412 ? _GEN_77032 : _GEN_77052; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_77073 = _T_7412 ? _GEN_77033 : _GEN_77053; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_77074 = _T_7412 ? _GEN_77034 : _GEN_77054; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_77075 = _T_7412 ? _GEN_77035 : _GEN_77055; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_77076 = _T_7412 ? _GEN_77036 : _GEN_77056; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_77077 = _T_7412 ? _GEN_77037 : _GEN_77057; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_77078 = _T_7412 ? _GEN_77038 : _GEN_77058; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_77079 = _T_7412 ? _GEN_77039 : _GEN_77059; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_77080 = _T_7412 ? _GEN_77040 : _GEN_77060; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_77081 = _T_7412 ? _GEN_77041 : _GEN_77061; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_77082 = _T_7412 ? _GEN_77042 : _GEN_77062; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_77083 = _T_7412 ? _GEN_77043 : _GEN_77063; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_77084 = _T_7412 ? _GEN_77044 : _GEN_77064; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_77085 = _T_7412 ? _GEN_77045 : _GEN_77065; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_77086 = _T_7412 ? _GEN_77046 : _GEN_77066; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_77087 = _T_7412 ? _GEN_77047 : _GEN_77067; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_77088 = _T_7412 ? _GEN_77048 : _GEN_77068; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_77089 = _T_7412 ? _GEN_77049 : _GEN_77069; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_77090 = _T_7412 ? _GEN_77050 : _GEN_77070; // @[FanCtrl.scala 377:65]
  wire [1:0] _GEN_77111 = r_valid_1 ? _GEN_77071 : _GEN_77031; // @[FanCtrl.scala 376:33]
  wire [1:0] _GEN_77112 = r_valid_1 ? _GEN_77072 : _GEN_77032; // @[FanCtrl.scala 376:33]
  wire [1:0] _GEN_77113 = r_valid_1 ? _GEN_77073 : _GEN_77033; // @[FanCtrl.scala 376:33]
  wire [1:0] _GEN_77114 = r_valid_1 ? _GEN_77074 : _GEN_77034; // @[FanCtrl.scala 376:33]
  wire [1:0] _GEN_77115 = r_valid_1 ? _GEN_77075 : _GEN_77035; // @[FanCtrl.scala 376:33]
  wire [1:0] _GEN_77116 = r_valid_1 ? _GEN_77076 : _GEN_77036; // @[FanCtrl.scala 376:33]
  wire [1:0] _GEN_77117 = r_valid_1 ? _GEN_77077 : _GEN_77037; // @[FanCtrl.scala 376:33]
  wire [1:0] _GEN_77118 = r_valid_1 ? _GEN_77078 : _GEN_77038; // @[FanCtrl.scala 376:33]
  wire [1:0] _GEN_77119 = r_valid_1 ? _GEN_77079 : _GEN_77039; // @[FanCtrl.scala 376:33]
  wire [1:0] _GEN_77120 = r_valid_1 ? _GEN_77080 : _GEN_77040; // @[FanCtrl.scala 376:33]
  wire [1:0] _GEN_77121 = r_valid_1 ? _GEN_77081 : _GEN_77041; // @[FanCtrl.scala 376:33]
  wire [1:0] _GEN_77122 = r_valid_1 ? _GEN_77082 : _GEN_77042; // @[FanCtrl.scala 376:33]
  wire [1:0] _GEN_77123 = r_valid_1 ? _GEN_77083 : _GEN_77043; // @[FanCtrl.scala 376:33]
  wire [1:0] _GEN_77124 = r_valid_1 ? _GEN_77084 : _GEN_77044; // @[FanCtrl.scala 376:33]
  wire [1:0] _GEN_77125 = r_valid_1 ? _GEN_77085 : _GEN_77045; // @[FanCtrl.scala 376:33]
  wire [1:0] _GEN_77126 = r_valid_1 ? _GEN_77086 : _GEN_77046; // @[FanCtrl.scala 376:33]
  wire [1:0] _GEN_77127 = r_valid_1 ? _GEN_77087 : _GEN_77047; // @[FanCtrl.scala 376:33]
  wire [1:0] _GEN_77128 = r_valid_1 ? _GEN_77088 : _GEN_77048; // @[FanCtrl.scala 376:33]
  wire [1:0] _GEN_77129 = r_valid_1 ? _GEN_77089 : _GEN_77049; // @[FanCtrl.scala 376:33]
  wire [1:0] _GEN_77130 = r_valid_1 ? _GEN_77090 : _GEN_77050; // @[FanCtrl.scala 376:33]
  wire [3:0] _T_7597 = _T_7440 + 4'h1; // @[FanCtrl.scala 392:39]
  wire [1:0] _GEN_77195 = 4'h0 == _T_7597 ? 2'h1 : _GEN_77111; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_77196 = 4'h1 == _T_7597 ? 2'h1 : _GEN_77112; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_77197 = 4'h2 == _T_7597 ? 2'h1 : _GEN_77113; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_77198 = 4'h3 == _T_7597 ? 2'h1 : _GEN_77114; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_77199 = 4'h4 == _T_7597 ? 2'h1 : _GEN_77115; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_77200 = 4'h5 == _T_7597 ? 2'h1 : _GEN_77116; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_77201 = 4'h6 == _T_7597 ? 2'h1 : _GEN_77117; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_77202 = 4'h7 == _T_7597 ? 2'h1 : _GEN_77118; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_77203 = 4'h8 == _T_7597 ? 2'h1 : _GEN_77119; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_77204 = 4'h9 == _T_7597 ? 2'h1 : _GEN_77120; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_77205 = 4'ha == _T_7597 ? 2'h1 : _GEN_77121; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_77206 = 4'hb == _T_7597 ? 2'h1 : _GEN_77122; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_77207 = 4'hc == _T_7597 ? 2'h1 : _GEN_77123; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_77208 = 4'hd == _T_7597 ? 2'h1 : _GEN_77124; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_77209 = 4'he == _T_7597 ? 2'h1 : _GEN_77125; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_77210 = 4'hf == _T_7597 ? 2'h1 : _GEN_77126; // @[FanCtrl.scala 392:{46,46}]
  wire [4:0] _GEN_97830 = {{1'd0}, _T_7597}; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_77211 = 5'h10 == _GEN_97830 ? 2'h1 : _GEN_77127; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_77212 = 5'h11 == _GEN_97830 ? 2'h1 : _GEN_77128; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_77213 = 5'h12 == _GEN_97830 ? 2'h1 : _GEN_77129; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_77214 = 5'h13 == _GEN_97830 ? 2'h1 : _GEN_77130; // @[FanCtrl.scala 392:{46,46}]
  wire [1:0] _GEN_77215 = 4'h0 == _T_7597 ? 2'h0 : _GEN_77111; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_77216 = 4'h1 == _T_7597 ? 2'h0 : _GEN_77112; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_77217 = 4'h2 == _T_7597 ? 2'h0 : _GEN_77113; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_77218 = 4'h3 == _T_7597 ? 2'h0 : _GEN_77114; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_77219 = 4'h4 == _T_7597 ? 2'h0 : _GEN_77115; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_77220 = 4'h5 == _T_7597 ? 2'h0 : _GEN_77116; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_77221 = 4'h6 == _T_7597 ? 2'h0 : _GEN_77117; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_77222 = 4'h7 == _T_7597 ? 2'h0 : _GEN_77118; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_77223 = 4'h8 == _T_7597 ? 2'h0 : _GEN_77119; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_77224 = 4'h9 == _T_7597 ? 2'h0 : _GEN_77120; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_77225 = 4'ha == _T_7597 ? 2'h0 : _GEN_77121; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_77226 = 4'hb == _T_7597 ? 2'h0 : _GEN_77122; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_77227 = 4'hc == _T_7597 ? 2'h0 : _GEN_77123; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_77228 = 4'hd == _T_7597 ? 2'h0 : _GEN_77124; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_77229 = 4'he == _T_7597 ? 2'h0 : _GEN_77125; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_77230 = 4'hf == _T_7597 ? 2'h0 : _GEN_77126; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_77231 = 5'h10 == _GEN_97830 ? 2'h0 : _GEN_77127; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_77232 = 5'h11 == _GEN_97830 ? 2'h0 : _GEN_77128; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_77233 = 5'h12 == _GEN_97830 ? 2'h0 : _GEN_77129; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_77234 = 5'h13 == _GEN_97830 ? 2'h0 : _GEN_77130; // @[FanCtrl.scala 395:{46,46}]
  wire [1:0] _GEN_77235 = _T_7428 ? _GEN_77195 : _GEN_77215; // @[FanCtrl.scala 390:64]
  wire [1:0] _GEN_77236 = _T_7428 ? _GEN_77196 : _GEN_77216; // @[FanCtrl.scala 390:64]
  wire [1:0] _GEN_77237 = _T_7428 ? _GEN_77197 : _GEN_77217; // @[FanCtrl.scala 390:64]
  wire [1:0] _GEN_77238 = _T_7428 ? _GEN_77198 : _GEN_77218; // @[FanCtrl.scala 390:64]
  wire [1:0] _GEN_77239 = _T_7428 ? _GEN_77199 : _GEN_77219; // @[FanCtrl.scala 390:64]
  wire [1:0] _GEN_77240 = _T_7428 ? _GEN_77200 : _GEN_77220; // @[FanCtrl.scala 390:64]
  wire [1:0] _GEN_77241 = _T_7428 ? _GEN_77201 : _GEN_77221; // @[FanCtrl.scala 390:64]
  wire [1:0] _GEN_77242 = _T_7428 ? _GEN_77202 : _GEN_77222; // @[FanCtrl.scala 390:64]
  wire [1:0] _GEN_77243 = _T_7428 ? _GEN_77203 : _GEN_77223; // @[FanCtrl.scala 390:64]
  wire [1:0] _GEN_77244 = _T_7428 ? _GEN_77204 : _GEN_77224; // @[FanCtrl.scala 390:64]
  wire [1:0] _GEN_77245 = _T_7428 ? _GEN_77205 : _GEN_77225; // @[FanCtrl.scala 390:64]
  wire [1:0] _GEN_77246 = _T_7428 ? _GEN_77206 : _GEN_77226; // @[FanCtrl.scala 390:64]
  wire [1:0] _GEN_77247 = _T_7428 ? _GEN_77207 : _GEN_77227; // @[FanCtrl.scala 390:64]
  wire [1:0] _GEN_77248 = _T_7428 ? _GEN_77208 : _GEN_77228; // @[FanCtrl.scala 390:64]
  wire [1:0] _GEN_77249 = _T_7428 ? _GEN_77209 : _GEN_77229; // @[FanCtrl.scala 390:64]
  wire [1:0] _GEN_77250 = _T_7428 ? _GEN_77210 : _GEN_77230; // @[FanCtrl.scala 390:64]
  wire [1:0] _GEN_77251 = _T_7428 ? _GEN_77211 : _GEN_77231; // @[FanCtrl.scala 390:64]
  wire [1:0] _GEN_77252 = _T_7428 ? _GEN_77212 : _GEN_77232; // @[FanCtrl.scala 390:64]
  wire [1:0] _GEN_77253 = _T_7428 ? _GEN_77213 : _GEN_77233; // @[FanCtrl.scala 390:64]
  wire [1:0] _GEN_77254 = _T_7428 ? _GEN_77214 : _GEN_77234; // @[FanCtrl.scala 390:64]
  wire [1:0] _GEN_77255 = 4'h0 == _T_7441[3:0] ? 2'h0 : _GEN_77111; // @[FanCtrl.scala 398:{44,44}]
  wire [1:0] _GEN_77256 = 4'h1 == _T_7441[3:0] ? 2'h0 : _GEN_77112; // @[FanCtrl.scala 398:{44,44}]
  wire [1:0] _GEN_77257 = 4'h2 == _T_7441[3:0] ? 2'h0 : _GEN_77113; // @[FanCtrl.scala 398:{44,44}]
  wire [1:0] _GEN_77258 = 4'h3 == _T_7441[3:0] ? 2'h0 : _GEN_77114; // @[FanCtrl.scala 398:{44,44}]
  wire [1:0] _GEN_77259 = 4'h4 == _T_7441[3:0] ? 2'h0 : _GEN_77115; // @[FanCtrl.scala 398:{44,44}]
  wire [1:0] _GEN_77260 = 4'h5 == _T_7441[3:0] ? 2'h0 : _GEN_77116; // @[FanCtrl.scala 398:{44,44}]
  wire [1:0] _GEN_77261 = 4'h6 == _T_7441[3:0] ? 2'h0 : _GEN_77117; // @[FanCtrl.scala 398:{44,44}]
  wire [1:0] _GEN_77262 = 4'h7 == _T_7441[3:0] ? 2'h0 : _GEN_77118; // @[FanCtrl.scala 398:{44,44}]
  wire [1:0] _GEN_77263 = 4'h8 == _T_7441[3:0] ? 2'h0 : _GEN_77119; // @[FanCtrl.scala 398:{44,44}]
  wire [1:0] _GEN_77264 = 4'h9 == _T_7441[3:0] ? 2'h0 : _GEN_77120; // @[FanCtrl.scala 398:{44,44}]
  wire [1:0] _GEN_77265 = 4'ha == _T_7441[3:0] ? 2'h0 : _GEN_77121; // @[FanCtrl.scala 398:{44,44}]
  wire [1:0] _GEN_77266 = 4'hb == _T_7441[3:0] ? 2'h0 : _GEN_77122; // @[FanCtrl.scala 398:{44,44}]
  wire [1:0] _GEN_77267 = 4'hc == _T_7441[3:0] ? 2'h0 : _GEN_77123; // @[FanCtrl.scala 398:{44,44}]
  wire [1:0] _GEN_77268 = 4'hd == _T_7441[3:0] ? 2'h0 : _GEN_77124; // @[FanCtrl.scala 398:{44,44}]
  wire [1:0] _GEN_77269 = 4'he == _T_7441[3:0] ? 2'h0 : _GEN_77125; // @[FanCtrl.scala 398:{44,44}]
  wire [1:0] _GEN_77270 = 4'hf == _T_7441[3:0] ? 2'h0 : _GEN_77126; // @[FanCtrl.scala 398:{44,44}]
  wire [1:0] _GEN_77271 = 5'h10 == _GEN_97814 ? 2'h0 : _GEN_77127; // @[FanCtrl.scala 398:{44,44}]
  wire [1:0] _GEN_77272 = 5'h11 == _GEN_97814 ? 2'h0 : _GEN_77128; // @[FanCtrl.scala 398:{44,44}]
  wire [1:0] _GEN_77273 = 5'h12 == _GEN_97814 ? 2'h0 : _GEN_77129; // @[FanCtrl.scala 398:{44,44}]
  wire [1:0] _GEN_77274 = 5'h13 == _GEN_97814 ? 2'h0 : _GEN_77130; // @[FanCtrl.scala 398:{44,44}]
  wire [1:0] _GEN_77275 = r_valid_1 ? _GEN_77235 : _GEN_77255; // @[FanCtrl.scala 389:33]
  wire [1:0] _GEN_77276 = r_valid_1 ? _GEN_77236 : _GEN_77256; // @[FanCtrl.scala 389:33]
  wire [1:0] _GEN_77277 = r_valid_1 ? _GEN_77237 : _GEN_77257; // @[FanCtrl.scala 389:33]
  wire [1:0] _GEN_77278 = r_valid_1 ? _GEN_77238 : _GEN_77258; // @[FanCtrl.scala 389:33]
  wire [1:0] _GEN_77279 = r_valid_1 ? _GEN_77239 : _GEN_77259; // @[FanCtrl.scala 389:33]
  wire [1:0] _GEN_77280 = r_valid_1 ? _GEN_77240 : _GEN_77260; // @[FanCtrl.scala 389:33]
  wire [1:0] _GEN_77281 = r_valid_1 ? _GEN_77241 : _GEN_77261; // @[FanCtrl.scala 389:33]
  wire [1:0] _GEN_77282 = r_valid_1 ? _GEN_77242 : _GEN_77262; // @[FanCtrl.scala 389:33]
  wire [1:0] _GEN_77283 = r_valid_1 ? _GEN_77243 : _GEN_77263; // @[FanCtrl.scala 389:33]
  wire [1:0] _GEN_77284 = r_valid_1 ? _GEN_77244 : _GEN_77264; // @[FanCtrl.scala 389:33]
  wire [1:0] _GEN_77285 = r_valid_1 ? _GEN_77245 : _GEN_77265; // @[FanCtrl.scala 389:33]
  wire [1:0] _GEN_77286 = r_valid_1 ? _GEN_77246 : _GEN_77266; // @[FanCtrl.scala 389:33]
  wire [1:0] _GEN_77287 = r_valid_1 ? _GEN_77247 : _GEN_77267; // @[FanCtrl.scala 389:33]
  wire [1:0] _GEN_77288 = r_valid_1 ? _GEN_77248 : _GEN_77268; // @[FanCtrl.scala 389:33]
  wire [1:0] _GEN_77289 = r_valid_1 ? _GEN_77249 : _GEN_77269; // @[FanCtrl.scala 389:33]
  wire [1:0] _GEN_77290 = r_valid_1 ? _GEN_77250 : _GEN_77270; // @[FanCtrl.scala 389:33]
  wire [1:0] _GEN_77291 = r_valid_1 ? _GEN_77251 : _GEN_77271; // @[FanCtrl.scala 389:33]
  wire [1:0] _GEN_77292 = r_valid_1 ? _GEN_77252 : _GEN_77272; // @[FanCtrl.scala 389:33]
  wire [1:0] _GEN_77293 = r_valid_1 ? _GEN_77253 : _GEN_77273; // @[FanCtrl.scala 389:33]
  wire [1:0] _GEN_77294 = r_valid_1 ? _GEN_77254 : _GEN_77274; // @[FanCtrl.scala 389:33]
  wire [3:0] _T_7797 = 1'h0 * 3'h4; // @[FanCtrl.scala 479:28]
  wire [3:0] _T_7799 = _T_7797 + 4'h8; // @[FanCtrl.scala 479:35]
  wire [1:0] _GEN_79197 = 4'h0 == _T_7799 ? 2'h0 : _GEN_77275; // @[FanCtrl.scala 479:{42,42}]
  wire [1:0] _GEN_79198 = 4'h1 == _T_7799 ? 2'h0 : _GEN_77276; // @[FanCtrl.scala 479:{42,42}]
  wire [1:0] _GEN_79199 = 4'h2 == _T_7799 ? 2'h0 : _GEN_77277; // @[FanCtrl.scala 479:{42,42}]
  wire [1:0] _GEN_79200 = 4'h3 == _T_7799 ? 2'h0 : _GEN_77278; // @[FanCtrl.scala 479:{42,42}]
  wire [1:0] _GEN_79201 = 4'h4 == _T_7799 ? 2'h0 : _GEN_77279; // @[FanCtrl.scala 479:{42,42}]
  wire [1:0] _GEN_79202 = 4'h5 == _T_7799 ? 2'h0 : _GEN_77280; // @[FanCtrl.scala 479:{42,42}]
  wire [1:0] _GEN_79203 = 4'h6 == _T_7799 ? 2'h0 : _GEN_77281; // @[FanCtrl.scala 479:{42,42}]
  wire [1:0] _GEN_79204 = 4'h7 == _T_7799 ? 2'h0 : _GEN_77282; // @[FanCtrl.scala 479:{42,42}]
  wire [1:0] _GEN_79205 = 4'h8 == _T_7799 ? 2'h0 : _GEN_77283; // @[FanCtrl.scala 479:{42,42}]
  wire [1:0] _GEN_79206 = 4'h9 == _T_7799 ? 2'h0 : _GEN_77284; // @[FanCtrl.scala 479:{42,42}]
  wire [1:0] _GEN_79207 = 4'ha == _T_7799 ? 2'h0 : _GEN_77285; // @[FanCtrl.scala 479:{42,42}]
  wire [1:0] _GEN_79208 = 4'hb == _T_7799 ? 2'h0 : _GEN_77286; // @[FanCtrl.scala 479:{42,42}]
  wire [1:0] _GEN_79209 = 4'hc == _T_7799 ? 2'h0 : _GEN_77287; // @[FanCtrl.scala 479:{42,42}]
  wire [1:0] _GEN_79210 = 4'hd == _T_7799 ? 2'h0 : _GEN_77288; // @[FanCtrl.scala 479:{42,42}]
  wire [1:0] _GEN_79211 = 4'he == _T_7799 ? 2'h0 : _GEN_77289; // @[FanCtrl.scala 479:{42,42}]
  wire [1:0] _GEN_79212 = 4'hf == _T_7799 ? 2'h0 : _GEN_77290; // @[FanCtrl.scala 479:{42,42}]
  wire [4:0] _GEN_97870 = {{1'd0}, _T_7799}; // @[FanCtrl.scala 479:{42,42}]
  wire [1:0] _GEN_79213 = 5'h10 == _GEN_97870 ? 2'h0 : _GEN_77291; // @[FanCtrl.scala 479:{42,42}]
  wire [1:0] _GEN_79214 = 5'h11 == _GEN_97870 ? 2'h0 : _GEN_77292; // @[FanCtrl.scala 479:{42,42}]
  wire [1:0] _GEN_79215 = 5'h12 == _GEN_97870 ? 2'h0 : _GEN_77293; // @[FanCtrl.scala 479:{42,42}]
  wire [1:0] _GEN_79216 = 5'h13 == _GEN_97870 ? 2'h0 : _GEN_77294; // @[FanCtrl.scala 479:{42,42}]
  wire [5:0] _T_7801 = 5'h10 * 1'h0; // @[FanCtrl.scala 483:25]
  wire [5:0] _T_7803 = _T_7801 + 6'h7; // @[FanCtrl.scala 483:31]
  wire [5:0] _T_7807 = _T_7801 + 6'h8; // @[FanCtrl.scala 483:59]
  wire [4:0] _GEN_79220 = 5'h3 == _T_7803[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_79221 = 5'h4 == _T_7803[4:0] ? w_vn_4 : _GEN_79220; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_79222 = 5'h5 == _T_7803[4:0] ? 5'h0 : _GEN_79221; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_79223 = 5'h6 == _T_7803[4:0] ? 5'h0 : _GEN_79222; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_79224 = 5'h7 == _T_7803[4:0] ? w_vn_7 : _GEN_79223; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_79225 = 5'h8 == _T_7803[4:0] ? w_vn_8 : _GEN_79224; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_79226 = 5'h9 == _T_7803[4:0] ? 5'h0 : _GEN_79225; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_79227 = 5'ha == _T_7803[4:0] ? 5'h0 : _GEN_79226; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_79228 = 5'hb == _T_7803[4:0] ? w_vn_11 : _GEN_79227; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_79229 = 5'hc == _T_7803[4:0] ? w_vn_12 : _GEN_79228; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_79230 = 5'hd == _T_7803[4:0] ? w_vn_13 : _GEN_79229; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_79231 = 5'he == _T_7803[4:0] ? 5'h0 : _GEN_79230; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_79232 = 5'hf == _T_7803[4:0] ? w_vn_15 : _GEN_79231; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_79233 = 5'h10 == _T_7803[4:0] ? w_vn_16 : _GEN_79232; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_79234 = 5'h11 == _T_7803[4:0] ? 5'h0 : _GEN_79233; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_79235 = 5'h12 == _T_7803[4:0] ? w_vn_18 : _GEN_79234; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_79236 = 5'h13 == _T_7803[4:0] ? 5'h0 : _GEN_79235; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_79237 = 5'h14 == _T_7803[4:0] ? 5'h0 : _GEN_79236; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_79238 = 5'h15 == _T_7803[4:0] ? 5'h0 : _GEN_79237; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_79239 = 5'h16 == _T_7803[4:0] ? 5'h0 : _GEN_79238; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_79240 = 5'h17 == _T_7803[4:0] ? w_vn_23 : _GEN_79239; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_79241 = 5'h18 == _T_7803[4:0] ? w_vn_24 : _GEN_79240; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_79242 = 5'h19 == _T_7803[4:0] ? 5'h0 : _GEN_79241; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_79243 = 5'h1a == _T_7803[4:0] ? 5'h0 : _GEN_79242; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_79244 = 5'h1b == _T_7803[4:0] ? 5'h0 : _GEN_79243; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_79245 = 5'h1c == _T_7803[4:0] ? 5'h0 : _GEN_79244; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_79246 = 5'h1d == _T_7803[4:0] ? 5'h0 : _GEN_79245; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_79247 = 5'h1e == _T_7803[4:0] ? 5'h0 : _GEN_79246; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_79248 = 5'h1f == _T_7803[4:0] ? 5'h0 : _GEN_79247; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_79252 = 5'h3 == _T_7807[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_79253 = 5'h4 == _T_7807[4:0] ? w_vn_4 : _GEN_79252; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_79254 = 5'h5 == _T_7807[4:0] ? 5'h0 : _GEN_79253; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_79255 = 5'h6 == _T_7807[4:0] ? 5'h0 : _GEN_79254; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_79256 = 5'h7 == _T_7807[4:0] ? w_vn_7 : _GEN_79255; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_79257 = 5'h8 == _T_7807[4:0] ? w_vn_8 : _GEN_79256; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_79258 = 5'h9 == _T_7807[4:0] ? 5'h0 : _GEN_79257; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_79259 = 5'ha == _T_7807[4:0] ? 5'h0 : _GEN_79258; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_79260 = 5'hb == _T_7807[4:0] ? w_vn_11 : _GEN_79259; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_79261 = 5'hc == _T_7807[4:0] ? w_vn_12 : _GEN_79260; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_79262 = 5'hd == _T_7807[4:0] ? w_vn_13 : _GEN_79261; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_79263 = 5'he == _T_7807[4:0] ? 5'h0 : _GEN_79262; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_79264 = 5'hf == _T_7807[4:0] ? w_vn_15 : _GEN_79263; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_79265 = 5'h10 == _T_7807[4:0] ? w_vn_16 : _GEN_79264; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_79266 = 5'h11 == _T_7807[4:0] ? 5'h0 : _GEN_79265; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_79267 = 5'h12 == _T_7807[4:0] ? w_vn_18 : _GEN_79266; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_79268 = 5'h13 == _T_7807[4:0] ? 5'h0 : _GEN_79267; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_79269 = 5'h14 == _T_7807[4:0] ? 5'h0 : _GEN_79268; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_79270 = 5'h15 == _T_7807[4:0] ? 5'h0 : _GEN_79269; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_79271 = 5'h16 == _T_7807[4:0] ? 5'h0 : _GEN_79270; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_79272 = 5'h17 == _T_7807[4:0] ? w_vn_23 : _GEN_79271; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_79273 = 5'h18 == _T_7807[4:0] ? w_vn_24 : _GEN_79272; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_79274 = 5'h19 == _T_7807[4:0] ? 5'h0 : _GEN_79273; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_79275 = 5'h1a == _T_7807[4:0] ? 5'h0 : _GEN_79274; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_79276 = 5'h1b == _T_7807[4:0] ? 5'h0 : _GEN_79275; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_79277 = 5'h1c == _T_7807[4:0] ? 5'h0 : _GEN_79276; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_79278 = 5'h1d == _T_7807[4:0] ? 5'h0 : _GEN_79277; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_79279 = 5'h1e == _T_7807[4:0] ? 5'h0 : _GEN_79278; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_79280 = 5'h1f == _T_7807[4:0] ? 5'h0 : _GEN_79279; // @[FanCtrl.scala 483:{39,39}]
  wire  _T_7809 = _GEN_79248 == _GEN_79280; // @[FanCtrl.scala 483:39]
  wire [5:0] _T_7816 = _T_7801 + 6'h3; // @[FanCtrl.scala 489:31]
  wire [5:0] _T_7820 = _T_7801 + 6'h4; // @[FanCtrl.scala 489:59]
  wire [4:0] _GEN_79377 = 5'h3 == _T_7816[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_79378 = 5'h4 == _T_7816[4:0] ? w_vn_4 : _GEN_79377; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_79379 = 5'h5 == _T_7816[4:0] ? 5'h0 : _GEN_79378; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_79380 = 5'h6 == _T_7816[4:0] ? 5'h0 : _GEN_79379; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_79381 = 5'h7 == _T_7816[4:0] ? w_vn_7 : _GEN_79380; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_79382 = 5'h8 == _T_7816[4:0] ? w_vn_8 : _GEN_79381; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_79383 = 5'h9 == _T_7816[4:0] ? 5'h0 : _GEN_79382; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_79384 = 5'ha == _T_7816[4:0] ? 5'h0 : _GEN_79383; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_79385 = 5'hb == _T_7816[4:0] ? w_vn_11 : _GEN_79384; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_79386 = 5'hc == _T_7816[4:0] ? w_vn_12 : _GEN_79385; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_79387 = 5'hd == _T_7816[4:0] ? w_vn_13 : _GEN_79386; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_79388 = 5'he == _T_7816[4:0] ? 5'h0 : _GEN_79387; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_79389 = 5'hf == _T_7816[4:0] ? w_vn_15 : _GEN_79388; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_79390 = 5'h10 == _T_7816[4:0] ? w_vn_16 : _GEN_79389; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_79391 = 5'h11 == _T_7816[4:0] ? 5'h0 : _GEN_79390; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_79392 = 5'h12 == _T_7816[4:0] ? w_vn_18 : _GEN_79391; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_79393 = 5'h13 == _T_7816[4:0] ? 5'h0 : _GEN_79392; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_79394 = 5'h14 == _T_7816[4:0] ? 5'h0 : _GEN_79393; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_79395 = 5'h15 == _T_7816[4:0] ? 5'h0 : _GEN_79394; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_79396 = 5'h16 == _T_7816[4:0] ? 5'h0 : _GEN_79395; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_79397 = 5'h17 == _T_7816[4:0] ? w_vn_23 : _GEN_79396; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_79398 = 5'h18 == _T_7816[4:0] ? w_vn_24 : _GEN_79397; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_79399 = 5'h19 == _T_7816[4:0] ? 5'h0 : _GEN_79398; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_79400 = 5'h1a == _T_7816[4:0] ? 5'h0 : _GEN_79399; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_79401 = 5'h1b == _T_7816[4:0] ? 5'h0 : _GEN_79400; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_79402 = 5'h1c == _T_7816[4:0] ? 5'h0 : _GEN_79401; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_79403 = 5'h1d == _T_7816[4:0] ? 5'h0 : _GEN_79402; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_79404 = 5'h1e == _T_7816[4:0] ? 5'h0 : _GEN_79403; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_79405 = 5'h1f == _T_7816[4:0] ? 5'h0 : _GEN_79404; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_79409 = 5'h3 == _T_7820[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_79410 = 5'h4 == _T_7820[4:0] ? w_vn_4 : _GEN_79409; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_79411 = 5'h5 == _T_7820[4:0] ? 5'h0 : _GEN_79410; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_79412 = 5'h6 == _T_7820[4:0] ? 5'h0 : _GEN_79411; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_79413 = 5'h7 == _T_7820[4:0] ? w_vn_7 : _GEN_79412; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_79414 = 5'h8 == _T_7820[4:0] ? w_vn_8 : _GEN_79413; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_79415 = 5'h9 == _T_7820[4:0] ? 5'h0 : _GEN_79414; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_79416 = 5'ha == _T_7820[4:0] ? 5'h0 : _GEN_79415; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_79417 = 5'hb == _T_7820[4:0] ? w_vn_11 : _GEN_79416; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_79418 = 5'hc == _T_7820[4:0] ? w_vn_12 : _GEN_79417; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_79419 = 5'hd == _T_7820[4:0] ? w_vn_13 : _GEN_79418; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_79420 = 5'he == _T_7820[4:0] ? 5'h0 : _GEN_79419; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_79421 = 5'hf == _T_7820[4:0] ? w_vn_15 : _GEN_79420; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_79422 = 5'h10 == _T_7820[4:0] ? w_vn_16 : _GEN_79421; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_79423 = 5'h11 == _T_7820[4:0] ? 5'h0 : _GEN_79422; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_79424 = 5'h12 == _T_7820[4:0] ? w_vn_18 : _GEN_79423; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_79425 = 5'h13 == _T_7820[4:0] ? 5'h0 : _GEN_79424; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_79426 = 5'h14 == _T_7820[4:0] ? 5'h0 : _GEN_79425; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_79427 = 5'h15 == _T_7820[4:0] ? 5'h0 : _GEN_79426; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_79428 = 5'h16 == _T_7820[4:0] ? 5'h0 : _GEN_79427; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_79429 = 5'h17 == _T_7820[4:0] ? w_vn_23 : _GEN_79428; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_79430 = 5'h18 == _T_7820[4:0] ? w_vn_24 : _GEN_79429; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_79431 = 5'h19 == _T_7820[4:0] ? 5'h0 : _GEN_79430; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_79432 = 5'h1a == _T_7820[4:0] ? 5'h0 : _GEN_79431; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_79433 = 5'h1b == _T_7820[4:0] ? 5'h0 : _GEN_79432; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_79434 = 5'h1c == _T_7820[4:0] ? 5'h0 : _GEN_79433; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_79435 = 5'h1d == _T_7820[4:0] ? 5'h0 : _GEN_79434; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_79436 = 5'h1e == _T_7820[4:0] ? 5'h0 : _GEN_79435; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_79437 = 5'h1f == _T_7820[4:0] ? 5'h0 : _GEN_79436; // @[FanCtrl.scala 489:{38,38}]
  wire  _T_7822 = _GEN_79405 == _GEN_79437; // @[FanCtrl.scala 489:38]
  wire [5:0] _T_7825 = _T_7801 + 6'hb; // @[FanCtrl.scala 490:32]
  wire [5:0] _T_7829 = _T_7801 + 6'hc; // @[FanCtrl.scala 490:61]
  wire [4:0] _GEN_79441 = 5'h3 == _T_7825[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_79442 = 5'h4 == _T_7825[4:0] ? w_vn_4 : _GEN_79441; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_79443 = 5'h5 == _T_7825[4:0] ? 5'h0 : _GEN_79442; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_79444 = 5'h6 == _T_7825[4:0] ? 5'h0 : _GEN_79443; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_79445 = 5'h7 == _T_7825[4:0] ? w_vn_7 : _GEN_79444; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_79446 = 5'h8 == _T_7825[4:0] ? w_vn_8 : _GEN_79445; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_79447 = 5'h9 == _T_7825[4:0] ? 5'h0 : _GEN_79446; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_79448 = 5'ha == _T_7825[4:0] ? 5'h0 : _GEN_79447; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_79449 = 5'hb == _T_7825[4:0] ? w_vn_11 : _GEN_79448; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_79450 = 5'hc == _T_7825[4:0] ? w_vn_12 : _GEN_79449; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_79451 = 5'hd == _T_7825[4:0] ? w_vn_13 : _GEN_79450; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_79452 = 5'he == _T_7825[4:0] ? 5'h0 : _GEN_79451; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_79453 = 5'hf == _T_7825[4:0] ? w_vn_15 : _GEN_79452; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_79454 = 5'h10 == _T_7825[4:0] ? w_vn_16 : _GEN_79453; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_79455 = 5'h11 == _T_7825[4:0] ? 5'h0 : _GEN_79454; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_79456 = 5'h12 == _T_7825[4:0] ? w_vn_18 : _GEN_79455; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_79457 = 5'h13 == _T_7825[4:0] ? 5'h0 : _GEN_79456; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_79458 = 5'h14 == _T_7825[4:0] ? 5'h0 : _GEN_79457; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_79459 = 5'h15 == _T_7825[4:0] ? 5'h0 : _GEN_79458; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_79460 = 5'h16 == _T_7825[4:0] ? 5'h0 : _GEN_79459; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_79461 = 5'h17 == _T_7825[4:0] ? w_vn_23 : _GEN_79460; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_79462 = 5'h18 == _T_7825[4:0] ? w_vn_24 : _GEN_79461; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_79463 = 5'h19 == _T_7825[4:0] ? 5'h0 : _GEN_79462; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_79464 = 5'h1a == _T_7825[4:0] ? 5'h0 : _GEN_79463; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_79465 = 5'h1b == _T_7825[4:0] ? 5'h0 : _GEN_79464; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_79466 = 5'h1c == _T_7825[4:0] ? 5'h0 : _GEN_79465; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_79467 = 5'h1d == _T_7825[4:0] ? 5'h0 : _GEN_79466; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_79468 = 5'h1e == _T_7825[4:0] ? 5'h0 : _GEN_79467; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_79469 = 5'h1f == _T_7825[4:0] ? 5'h0 : _GEN_79468; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_79473 = 5'h3 == _T_7829[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_79474 = 5'h4 == _T_7829[4:0] ? w_vn_4 : _GEN_79473; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_79475 = 5'h5 == _T_7829[4:0] ? 5'h0 : _GEN_79474; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_79476 = 5'h6 == _T_7829[4:0] ? 5'h0 : _GEN_79475; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_79477 = 5'h7 == _T_7829[4:0] ? w_vn_7 : _GEN_79476; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_79478 = 5'h8 == _T_7829[4:0] ? w_vn_8 : _GEN_79477; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_79479 = 5'h9 == _T_7829[4:0] ? 5'h0 : _GEN_79478; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_79480 = 5'ha == _T_7829[4:0] ? 5'h0 : _GEN_79479; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_79481 = 5'hb == _T_7829[4:0] ? w_vn_11 : _GEN_79480; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_79482 = 5'hc == _T_7829[4:0] ? w_vn_12 : _GEN_79481; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_79483 = 5'hd == _T_7829[4:0] ? w_vn_13 : _GEN_79482; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_79484 = 5'he == _T_7829[4:0] ? 5'h0 : _GEN_79483; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_79485 = 5'hf == _T_7829[4:0] ? w_vn_15 : _GEN_79484; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_79486 = 5'h10 == _T_7829[4:0] ? w_vn_16 : _GEN_79485; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_79487 = 5'h11 == _T_7829[4:0] ? 5'h0 : _GEN_79486; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_79488 = 5'h12 == _T_7829[4:0] ? w_vn_18 : _GEN_79487; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_79489 = 5'h13 == _T_7829[4:0] ? 5'h0 : _GEN_79488; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_79490 = 5'h14 == _T_7829[4:0] ? 5'h0 : _GEN_79489; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_79491 = 5'h15 == _T_7829[4:0] ? 5'h0 : _GEN_79490; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_79492 = 5'h16 == _T_7829[4:0] ? 5'h0 : _GEN_79491; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_79493 = 5'h17 == _T_7829[4:0] ? w_vn_23 : _GEN_79492; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_79494 = 5'h18 == _T_7829[4:0] ? w_vn_24 : _GEN_79493; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_79495 = 5'h19 == _T_7829[4:0] ? 5'h0 : _GEN_79494; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_79496 = 5'h1a == _T_7829[4:0] ? 5'h0 : _GEN_79495; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_79497 = 5'h1b == _T_7829[4:0] ? 5'h0 : _GEN_79496; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_79498 = 5'h1c == _T_7829[4:0] ? 5'h0 : _GEN_79497; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_79499 = 5'h1d == _T_7829[4:0] ? 5'h0 : _GEN_79498; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_79500 = 5'h1e == _T_7829[4:0] ? 5'h0 : _GEN_79499; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_79501 = 5'h1f == _T_7829[4:0] ? 5'h0 : _GEN_79500; // @[FanCtrl.scala 490:{41,41}]
  wire  _T_7831 = _GEN_79469 == _GEN_79501; // @[FanCtrl.scala 490:41]
  wire  _T_7832 = _GEN_79405 == _GEN_79437 & _T_7831; // @[FanCtrl.scala 489:68]
  wire [5:0] _T_7835 = _T_7801 + 6'h10; // @[FanCtrl.scala 491:32]
  wire [4:0] _GEN_79505 = 5'h3 == _T_7835[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 491:{40,40}]
  wire [4:0] _GEN_79506 = 5'h4 == _T_7835[4:0] ? w_vn_4 : _GEN_79505; // @[FanCtrl.scala 491:{40,40}]
  wire [4:0] _GEN_79507 = 5'h5 == _T_7835[4:0] ? 5'h0 : _GEN_79506; // @[FanCtrl.scala 491:{40,40}]
  wire [4:0] _GEN_79508 = 5'h6 == _T_7835[4:0] ? 5'h0 : _GEN_79507; // @[FanCtrl.scala 491:{40,40}]
  wire [4:0] _GEN_79509 = 5'h7 == _T_7835[4:0] ? w_vn_7 : _GEN_79508; // @[FanCtrl.scala 491:{40,40}]
  wire [4:0] _GEN_79510 = 5'h8 == _T_7835[4:0] ? w_vn_8 : _GEN_79509; // @[FanCtrl.scala 491:{40,40}]
  wire [4:0] _GEN_79511 = 5'h9 == _T_7835[4:0] ? 5'h0 : _GEN_79510; // @[FanCtrl.scala 491:{40,40}]
  wire [4:0] _GEN_79512 = 5'ha == _T_7835[4:0] ? 5'h0 : _GEN_79511; // @[FanCtrl.scala 491:{40,40}]
  wire [4:0] _GEN_79513 = 5'hb == _T_7835[4:0] ? w_vn_11 : _GEN_79512; // @[FanCtrl.scala 491:{40,40}]
  wire [4:0] _GEN_79514 = 5'hc == _T_7835[4:0] ? w_vn_12 : _GEN_79513; // @[FanCtrl.scala 491:{40,40}]
  wire [4:0] _GEN_79515 = 5'hd == _T_7835[4:0] ? w_vn_13 : _GEN_79514; // @[FanCtrl.scala 491:{40,40}]
  wire [4:0] _GEN_79516 = 5'he == _T_7835[4:0] ? 5'h0 : _GEN_79515; // @[FanCtrl.scala 491:{40,40}]
  wire [4:0] _GEN_79517 = 5'hf == _T_7835[4:0] ? w_vn_15 : _GEN_79516; // @[FanCtrl.scala 491:{40,40}]
  wire [4:0] _GEN_79518 = 5'h10 == _T_7835[4:0] ? w_vn_16 : _GEN_79517; // @[FanCtrl.scala 491:{40,40}]
  wire [4:0] _GEN_79519 = 5'h11 == _T_7835[4:0] ? 5'h0 : _GEN_79518; // @[FanCtrl.scala 491:{40,40}]
  wire [4:0] _GEN_79520 = 5'h12 == _T_7835[4:0] ? w_vn_18 : _GEN_79519; // @[FanCtrl.scala 491:{40,40}]
  wire [4:0] _GEN_79521 = 5'h13 == _T_7835[4:0] ? 5'h0 : _GEN_79520; // @[FanCtrl.scala 491:{40,40}]
  wire [4:0] _GEN_79522 = 5'h14 == _T_7835[4:0] ? 5'h0 : _GEN_79521; // @[FanCtrl.scala 491:{40,40}]
  wire [4:0] _GEN_79523 = 5'h15 == _T_7835[4:0] ? 5'h0 : _GEN_79522; // @[FanCtrl.scala 491:{40,40}]
  wire [4:0] _GEN_79524 = 5'h16 == _T_7835[4:0] ? 5'h0 : _GEN_79523; // @[FanCtrl.scala 491:{40,40}]
  wire [4:0] _GEN_79525 = 5'h17 == _T_7835[4:0] ? w_vn_23 : _GEN_79524; // @[FanCtrl.scala 491:{40,40}]
  wire [4:0] _GEN_79526 = 5'h18 == _T_7835[4:0] ? w_vn_24 : _GEN_79525; // @[FanCtrl.scala 491:{40,40}]
  wire [4:0] _GEN_79527 = 5'h19 == _T_7835[4:0] ? 5'h0 : _GEN_79526; // @[FanCtrl.scala 491:{40,40}]
  wire [4:0] _GEN_79528 = 5'h1a == _T_7835[4:0] ? 5'h0 : _GEN_79527; // @[FanCtrl.scala 491:{40,40}]
  wire [4:0] _GEN_79529 = 5'h1b == _T_7835[4:0] ? 5'h0 : _GEN_79528; // @[FanCtrl.scala 491:{40,40}]
  wire [4:0] _GEN_79530 = 5'h1c == _T_7835[4:0] ? 5'h0 : _GEN_79529; // @[FanCtrl.scala 491:{40,40}]
  wire [4:0] _GEN_79531 = 5'h1d == _T_7835[4:0] ? 5'h0 : _GEN_79530; // @[FanCtrl.scala 491:{40,40}]
  wire [4:0] _GEN_79532 = 5'h1e == _T_7835[4:0] ? 5'h0 : _GEN_79531; // @[FanCtrl.scala 491:{40,40}]
  wire [4:0] _GEN_79533 = 5'h1f == _T_7835[4:0] ? 5'h0 : _GEN_79532; // @[FanCtrl.scala 491:{40,40}]
  wire  _T_7841 = _GEN_79533 != _GEN_79501; // @[FanCtrl.scala 491:40]
  wire  _T_7842 = _T_7832 & _T_7841; // @[FanCtrl.scala 490:71]
  wire  _T_7851 = _GEN_79437 != _GEN_79280; // @[FanCtrl.scala 492:40]
  wire  _T_7852 = _T_7842 & _T_7851; // @[FanCtrl.scala 491:69]
  wire  _T_7861 = _GEN_79469 != _GEN_79248; // @[FanCtrl.scala 493:41]
  wire  _T_7862 = _T_7852 & _T_7861; // @[FanCtrl.scala 492:69]
  wire  _T_7883 = _T_7831 & _T_7841; // @[FanCtrl.scala 497:74]
  wire  _T_7893 = _T_7883 & _T_7861; // @[FanCtrl.scala 498:74]
  wire  _T_7914 = _T_7822 & _T_7851; // @[FanCtrl.scala 503:73]
  wire [2:0] _GEN_80166 = _T_7914 ? 3'h3 : 3'h0; // @[FanCtrl.scala 504:74]
  wire  _GEN_80321 = r_valid_1 & _T_7809; // @[FanCtrl.scala 482:33]
  wire [1:0] _GEN_80419 = 4'h0 == _T_7799 ? 2'h0 : _GEN_79197; // @[FanCtrl.scala 520:{46,46}]
  wire [1:0] _GEN_80420 = 4'h1 == _T_7799 ? 2'h0 : _GEN_79198; // @[FanCtrl.scala 520:{46,46}]
  wire [1:0] _GEN_80421 = 4'h2 == _T_7799 ? 2'h0 : _GEN_79199; // @[FanCtrl.scala 520:{46,46}]
  wire [1:0] _GEN_80422 = 4'h3 == _T_7799 ? 2'h0 : _GEN_79200; // @[FanCtrl.scala 520:{46,46}]
  wire [1:0] _GEN_80423 = 4'h4 == _T_7799 ? 2'h0 : _GEN_79201; // @[FanCtrl.scala 520:{46,46}]
  wire [1:0] _GEN_80424 = 4'h5 == _T_7799 ? 2'h0 : _GEN_79202; // @[FanCtrl.scala 520:{46,46}]
  wire [1:0] _GEN_80425 = 4'h6 == _T_7799 ? 2'h0 : _GEN_79203; // @[FanCtrl.scala 520:{46,46}]
  wire [1:0] _GEN_80426 = 4'h7 == _T_7799 ? 2'h0 : _GEN_79204; // @[FanCtrl.scala 520:{46,46}]
  wire [1:0] _GEN_80427 = 4'h8 == _T_7799 ? 2'h0 : _GEN_79205; // @[FanCtrl.scala 520:{46,46}]
  wire [1:0] _GEN_80428 = 4'h9 == _T_7799 ? 2'h0 : _GEN_79206; // @[FanCtrl.scala 520:{46,46}]
  wire [1:0] _GEN_80429 = 4'ha == _T_7799 ? 2'h0 : _GEN_79207; // @[FanCtrl.scala 520:{46,46}]
  wire [1:0] _GEN_80430 = 4'hb == _T_7799 ? 2'h0 : _GEN_79208; // @[FanCtrl.scala 520:{46,46}]
  wire [1:0] _GEN_80431 = 4'hc == _T_7799 ? 2'h0 : _GEN_79209; // @[FanCtrl.scala 520:{46,46}]
  wire [1:0] _GEN_80432 = 4'hd == _T_7799 ? 2'h0 : _GEN_79210; // @[FanCtrl.scala 520:{46,46}]
  wire [1:0] _GEN_80433 = 4'he == _T_7799 ? 2'h0 : _GEN_79211; // @[FanCtrl.scala 520:{46,46}]
  wire [1:0] _GEN_80434 = 4'hf == _T_7799 ? 2'h0 : _GEN_79212; // @[FanCtrl.scala 520:{46,46}]
  wire [1:0] _GEN_80435 = 5'h10 == _GEN_97870 ? 2'h0 : _GEN_79213; // @[FanCtrl.scala 520:{46,46}]
  wire [1:0] _GEN_80436 = 5'h11 == _GEN_97870 ? 2'h0 : _GEN_79214; // @[FanCtrl.scala 520:{46,46}]
  wire [1:0] _GEN_80437 = 5'h12 == _GEN_97870 ? 2'h0 : _GEN_79215; // @[FanCtrl.scala 520:{46,46}]
  wire [1:0] _GEN_80438 = 5'h13 == _GEN_97870 ? 2'h0 : _GEN_79216; // @[FanCtrl.scala 520:{46,46}]
  wire [5:0] _T_7942 = _T_7801 + 6'h5; // @[FanCtrl.scala 522:65]
  wire [4:0] _GEN_80474 = 5'h3 == _T_7942[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 522:{45,45}]
  wire [4:0] _GEN_80475 = 5'h4 == _T_7942[4:0] ? w_vn_4 : _GEN_80474; // @[FanCtrl.scala 522:{45,45}]
  wire [4:0] _GEN_80476 = 5'h5 == _T_7942[4:0] ? 5'h0 : _GEN_80475; // @[FanCtrl.scala 522:{45,45}]
  wire [4:0] _GEN_80477 = 5'h6 == _T_7942[4:0] ? 5'h0 : _GEN_80476; // @[FanCtrl.scala 522:{45,45}]
  wire [4:0] _GEN_80478 = 5'h7 == _T_7942[4:0] ? w_vn_7 : _GEN_80477; // @[FanCtrl.scala 522:{45,45}]
  wire [4:0] _GEN_80479 = 5'h8 == _T_7942[4:0] ? w_vn_8 : _GEN_80478; // @[FanCtrl.scala 522:{45,45}]
  wire [4:0] _GEN_80480 = 5'h9 == _T_7942[4:0] ? 5'h0 : _GEN_80479; // @[FanCtrl.scala 522:{45,45}]
  wire [4:0] _GEN_80481 = 5'ha == _T_7942[4:0] ? 5'h0 : _GEN_80480; // @[FanCtrl.scala 522:{45,45}]
  wire [4:0] _GEN_80482 = 5'hb == _T_7942[4:0] ? w_vn_11 : _GEN_80481; // @[FanCtrl.scala 522:{45,45}]
  wire [4:0] _GEN_80483 = 5'hc == _T_7942[4:0] ? w_vn_12 : _GEN_80482; // @[FanCtrl.scala 522:{45,45}]
  wire [4:0] _GEN_80484 = 5'hd == _T_7942[4:0] ? w_vn_13 : _GEN_80483; // @[FanCtrl.scala 522:{45,45}]
  wire [4:0] _GEN_80485 = 5'he == _T_7942[4:0] ? 5'h0 : _GEN_80484; // @[FanCtrl.scala 522:{45,45}]
  wire [4:0] _GEN_80486 = 5'hf == _T_7942[4:0] ? w_vn_15 : _GEN_80485; // @[FanCtrl.scala 522:{45,45}]
  wire [4:0] _GEN_80487 = 5'h10 == _T_7942[4:0] ? w_vn_16 : _GEN_80486; // @[FanCtrl.scala 522:{45,45}]
  wire [4:0] _GEN_80488 = 5'h11 == _T_7942[4:0] ? 5'h0 : _GEN_80487; // @[FanCtrl.scala 522:{45,45}]
  wire [4:0] _GEN_80489 = 5'h12 == _T_7942[4:0] ? w_vn_18 : _GEN_80488; // @[FanCtrl.scala 522:{45,45}]
  wire [4:0] _GEN_80490 = 5'h13 == _T_7942[4:0] ? 5'h0 : _GEN_80489; // @[FanCtrl.scala 522:{45,45}]
  wire [4:0] _GEN_80491 = 5'h14 == _T_7942[4:0] ? 5'h0 : _GEN_80490; // @[FanCtrl.scala 522:{45,45}]
  wire [4:0] _GEN_80492 = 5'h15 == _T_7942[4:0] ? 5'h0 : _GEN_80491; // @[FanCtrl.scala 522:{45,45}]
  wire [4:0] _GEN_80493 = 5'h16 == _T_7942[4:0] ? 5'h0 : _GEN_80492; // @[FanCtrl.scala 522:{45,45}]
  wire [4:0] _GEN_80494 = 5'h17 == _T_7942[4:0] ? w_vn_23 : _GEN_80493; // @[FanCtrl.scala 522:{45,45}]
  wire [4:0] _GEN_80495 = 5'h18 == _T_7942[4:0] ? w_vn_24 : _GEN_80494; // @[FanCtrl.scala 522:{45,45}]
  wire [4:0] _GEN_80496 = 5'h19 == _T_7942[4:0] ? 5'h0 : _GEN_80495; // @[FanCtrl.scala 522:{45,45}]
  wire [4:0] _GEN_80497 = 5'h1a == _T_7942[4:0] ? 5'h0 : _GEN_80496; // @[FanCtrl.scala 522:{45,45}]
  wire [4:0] _GEN_80498 = 5'h1b == _T_7942[4:0] ? 5'h0 : _GEN_80497; // @[FanCtrl.scala 522:{45,45}]
  wire [4:0] _GEN_80499 = 5'h1c == _T_7942[4:0] ? 5'h0 : _GEN_80498; // @[FanCtrl.scala 522:{45,45}]
  wire [4:0] _GEN_80500 = 5'h1d == _T_7942[4:0] ? 5'h0 : _GEN_80499; // @[FanCtrl.scala 522:{45,45}]
  wire [4:0] _GEN_80501 = 5'h1e == _T_7942[4:0] ? 5'h0 : _GEN_80500; // @[FanCtrl.scala 522:{45,45}]
  wire [4:0] _GEN_80502 = 5'h1f == _T_7942[4:0] ? 5'h0 : _GEN_80501; // @[FanCtrl.scala 522:{45,45}]
  wire [1:0] _GEN_80503 = 4'h0 == _T_7799 ? 2'h1 : _GEN_79197; // @[FanCtrl.scala 524:{45,45}]
  wire [1:0] _GEN_80504 = 4'h1 == _T_7799 ? 2'h1 : _GEN_79198; // @[FanCtrl.scala 524:{45,45}]
  wire [1:0] _GEN_80505 = 4'h2 == _T_7799 ? 2'h1 : _GEN_79199; // @[FanCtrl.scala 524:{45,45}]
  wire [1:0] _GEN_80506 = 4'h3 == _T_7799 ? 2'h1 : _GEN_79200; // @[FanCtrl.scala 524:{45,45}]
  wire [1:0] _GEN_80507 = 4'h4 == _T_7799 ? 2'h1 : _GEN_79201; // @[FanCtrl.scala 524:{45,45}]
  wire [1:0] _GEN_80508 = 4'h5 == _T_7799 ? 2'h1 : _GEN_79202; // @[FanCtrl.scala 524:{45,45}]
  wire [1:0] _GEN_80509 = 4'h6 == _T_7799 ? 2'h1 : _GEN_79203; // @[FanCtrl.scala 524:{45,45}]
  wire [1:0] _GEN_80510 = 4'h7 == _T_7799 ? 2'h1 : _GEN_79204; // @[FanCtrl.scala 524:{45,45}]
  wire [1:0] _GEN_80511 = 4'h8 == _T_7799 ? 2'h1 : _GEN_79205; // @[FanCtrl.scala 524:{45,45}]
  wire [1:0] _GEN_80512 = 4'h9 == _T_7799 ? 2'h1 : _GEN_79206; // @[FanCtrl.scala 524:{45,45}]
  wire [1:0] _GEN_80513 = 4'ha == _T_7799 ? 2'h1 : _GEN_79207; // @[FanCtrl.scala 524:{45,45}]
  wire [1:0] _GEN_80514 = 4'hb == _T_7799 ? 2'h1 : _GEN_79208; // @[FanCtrl.scala 524:{45,45}]
  wire [1:0] _GEN_80515 = 4'hc == _T_7799 ? 2'h1 : _GEN_79209; // @[FanCtrl.scala 524:{45,45}]
  wire [1:0] _GEN_80516 = 4'hd == _T_7799 ? 2'h1 : _GEN_79210; // @[FanCtrl.scala 524:{45,45}]
  wire [1:0] _GEN_80517 = 4'he == _T_7799 ? 2'h1 : _GEN_79211; // @[FanCtrl.scala 524:{45,45}]
  wire [1:0] _GEN_80518 = 4'hf == _T_7799 ? 2'h1 : _GEN_79212; // @[FanCtrl.scala 524:{45,45}]
  wire [1:0] _GEN_80519 = 5'h10 == _GEN_97870 ? 2'h1 : _GEN_79213; // @[FanCtrl.scala 524:{45,45}]
  wire [1:0] _GEN_80520 = 5'h11 == _GEN_97870 ? 2'h1 : _GEN_79214; // @[FanCtrl.scala 524:{45,45}]
  wire [1:0] _GEN_80521 = 5'h12 == _GEN_97870 ? 2'h1 : _GEN_79215; // @[FanCtrl.scala 524:{45,45}]
  wire [1:0] _GEN_80522 = 5'h13 == _GEN_97870 ? 2'h1 : _GEN_79216; // @[FanCtrl.scala 524:{45,45}]
  wire [1:0] _GEN_80523 = 4'h0 == _T_7799 ? 2'h2 : _GEN_79197; // @[FanCtrl.scala 528:{46,46}]
  wire [1:0] _GEN_80524 = 4'h1 == _T_7799 ? 2'h2 : _GEN_79198; // @[FanCtrl.scala 528:{46,46}]
  wire [1:0] _GEN_80525 = 4'h2 == _T_7799 ? 2'h2 : _GEN_79199; // @[FanCtrl.scala 528:{46,46}]
  wire [1:0] _GEN_80526 = 4'h3 == _T_7799 ? 2'h2 : _GEN_79200; // @[FanCtrl.scala 528:{46,46}]
  wire [1:0] _GEN_80527 = 4'h4 == _T_7799 ? 2'h2 : _GEN_79201; // @[FanCtrl.scala 528:{46,46}]
  wire [1:0] _GEN_80528 = 4'h5 == _T_7799 ? 2'h2 : _GEN_79202; // @[FanCtrl.scala 528:{46,46}]
  wire [1:0] _GEN_80529 = 4'h6 == _T_7799 ? 2'h2 : _GEN_79203; // @[FanCtrl.scala 528:{46,46}]
  wire [1:0] _GEN_80530 = 4'h7 == _T_7799 ? 2'h2 : _GEN_79204; // @[FanCtrl.scala 528:{46,46}]
  wire [1:0] _GEN_80531 = 4'h8 == _T_7799 ? 2'h2 : _GEN_79205; // @[FanCtrl.scala 528:{46,46}]
  wire [1:0] _GEN_80532 = 4'h9 == _T_7799 ? 2'h2 : _GEN_79206; // @[FanCtrl.scala 528:{46,46}]
  wire [1:0] _GEN_80533 = 4'ha == _T_7799 ? 2'h2 : _GEN_79207; // @[FanCtrl.scala 528:{46,46}]
  wire [1:0] _GEN_80534 = 4'hb == _T_7799 ? 2'h2 : _GEN_79208; // @[FanCtrl.scala 528:{46,46}]
  wire [1:0] _GEN_80535 = 4'hc == _T_7799 ? 2'h2 : _GEN_79209; // @[FanCtrl.scala 528:{46,46}]
  wire [1:0] _GEN_80536 = 4'hd == _T_7799 ? 2'h2 : _GEN_79210; // @[FanCtrl.scala 528:{46,46}]
  wire [1:0] _GEN_80537 = 4'he == _T_7799 ? 2'h2 : _GEN_79211; // @[FanCtrl.scala 528:{46,46}]
  wire [1:0] _GEN_80538 = 4'hf == _T_7799 ? 2'h2 : _GEN_79212; // @[FanCtrl.scala 528:{46,46}]
  wire [1:0] _GEN_80539 = 5'h10 == _GEN_97870 ? 2'h2 : _GEN_79213; // @[FanCtrl.scala 528:{46,46}]
  wire [1:0] _GEN_80540 = 5'h11 == _GEN_97870 ? 2'h2 : _GEN_79214; // @[FanCtrl.scala 528:{46,46}]
  wire [1:0] _GEN_80541 = 5'h12 == _GEN_97870 ? 2'h2 : _GEN_79215; // @[FanCtrl.scala 528:{46,46}]
  wire [1:0] _GEN_80542 = 5'h13 == _GEN_97870 ? 2'h2 : _GEN_79216; // @[FanCtrl.scala 528:{46,46}]
  wire [1:0] _GEN_80543 = _GEN_79248 == _GEN_80502 ? _GEN_80503 : _GEN_80523; // @[FanCtrl.scala 522:74]
  wire [1:0] _GEN_80544 = _GEN_79248 == _GEN_80502 ? _GEN_80504 : _GEN_80524; // @[FanCtrl.scala 522:74]
  wire [1:0] _GEN_80545 = _GEN_79248 == _GEN_80502 ? _GEN_80505 : _GEN_80525; // @[FanCtrl.scala 522:74]
  wire [1:0] _GEN_80546 = _GEN_79248 == _GEN_80502 ? _GEN_80506 : _GEN_80526; // @[FanCtrl.scala 522:74]
  wire [1:0] _GEN_80547 = _GEN_79248 == _GEN_80502 ? _GEN_80507 : _GEN_80527; // @[FanCtrl.scala 522:74]
  wire [1:0] _GEN_80548 = _GEN_79248 == _GEN_80502 ? _GEN_80508 : _GEN_80528; // @[FanCtrl.scala 522:74]
  wire [1:0] _GEN_80549 = _GEN_79248 == _GEN_80502 ? _GEN_80509 : _GEN_80529; // @[FanCtrl.scala 522:74]
  wire [1:0] _GEN_80550 = _GEN_79248 == _GEN_80502 ? _GEN_80510 : _GEN_80530; // @[FanCtrl.scala 522:74]
  wire [1:0] _GEN_80551 = _GEN_79248 == _GEN_80502 ? _GEN_80511 : _GEN_80531; // @[FanCtrl.scala 522:74]
  wire [1:0] _GEN_80552 = _GEN_79248 == _GEN_80502 ? _GEN_80512 : _GEN_80532; // @[FanCtrl.scala 522:74]
  wire [1:0] _GEN_80553 = _GEN_79248 == _GEN_80502 ? _GEN_80513 : _GEN_80533; // @[FanCtrl.scala 522:74]
  wire [1:0] _GEN_80554 = _GEN_79248 == _GEN_80502 ? _GEN_80514 : _GEN_80534; // @[FanCtrl.scala 522:74]
  wire [1:0] _GEN_80555 = _GEN_79248 == _GEN_80502 ? _GEN_80515 : _GEN_80535; // @[FanCtrl.scala 522:74]
  wire [1:0] _GEN_80556 = _GEN_79248 == _GEN_80502 ? _GEN_80516 : _GEN_80536; // @[FanCtrl.scala 522:74]
  wire [1:0] _GEN_80557 = _GEN_79248 == _GEN_80502 ? _GEN_80517 : _GEN_80537; // @[FanCtrl.scala 522:74]
  wire [1:0] _GEN_80558 = _GEN_79248 == _GEN_80502 ? _GEN_80518 : _GEN_80538; // @[FanCtrl.scala 522:74]
  wire [1:0] _GEN_80559 = _GEN_79248 == _GEN_80502 ? _GEN_80519 : _GEN_80539; // @[FanCtrl.scala 522:74]
  wire [1:0] _GEN_80560 = _GEN_79248 == _GEN_80502 ? _GEN_80520 : _GEN_80540; // @[FanCtrl.scala 522:74]
  wire [1:0] _GEN_80561 = _GEN_79248 == _GEN_80502 ? _GEN_80521 : _GEN_80541; // @[FanCtrl.scala 522:74]
  wire [1:0] _GEN_80562 = _GEN_79248 == _GEN_80502 ? _GEN_80522 : _GEN_80542; // @[FanCtrl.scala 522:74]
  wire [1:0] _GEN_80563 = _GEN_79248 == _GEN_79405 ? _GEN_80419 : _GEN_80543; // @[FanCtrl.scala 518:68]
  wire [1:0] _GEN_80564 = _GEN_79248 == _GEN_79405 ? _GEN_80420 : _GEN_80544; // @[FanCtrl.scala 518:68]
  wire [1:0] _GEN_80565 = _GEN_79248 == _GEN_79405 ? _GEN_80421 : _GEN_80545; // @[FanCtrl.scala 518:68]
  wire [1:0] _GEN_80566 = _GEN_79248 == _GEN_79405 ? _GEN_80422 : _GEN_80546; // @[FanCtrl.scala 518:68]
  wire [1:0] _GEN_80567 = _GEN_79248 == _GEN_79405 ? _GEN_80423 : _GEN_80547; // @[FanCtrl.scala 518:68]
  wire [1:0] _GEN_80568 = _GEN_79248 == _GEN_79405 ? _GEN_80424 : _GEN_80548; // @[FanCtrl.scala 518:68]
  wire [1:0] _GEN_80569 = _GEN_79248 == _GEN_79405 ? _GEN_80425 : _GEN_80549; // @[FanCtrl.scala 518:68]
  wire [1:0] _GEN_80570 = _GEN_79248 == _GEN_79405 ? _GEN_80426 : _GEN_80550; // @[FanCtrl.scala 518:68]
  wire [1:0] _GEN_80571 = _GEN_79248 == _GEN_79405 ? _GEN_80427 : _GEN_80551; // @[FanCtrl.scala 518:68]
  wire [1:0] _GEN_80572 = _GEN_79248 == _GEN_79405 ? _GEN_80428 : _GEN_80552; // @[FanCtrl.scala 518:68]
  wire [1:0] _GEN_80573 = _GEN_79248 == _GEN_79405 ? _GEN_80429 : _GEN_80553; // @[FanCtrl.scala 518:68]
  wire [1:0] _GEN_80574 = _GEN_79248 == _GEN_79405 ? _GEN_80430 : _GEN_80554; // @[FanCtrl.scala 518:68]
  wire [1:0] _GEN_80575 = _GEN_79248 == _GEN_79405 ? _GEN_80431 : _GEN_80555; // @[FanCtrl.scala 518:68]
  wire [1:0] _GEN_80576 = _GEN_79248 == _GEN_79405 ? _GEN_80432 : _GEN_80556; // @[FanCtrl.scala 518:68]
  wire [1:0] _GEN_80577 = _GEN_79248 == _GEN_79405 ? _GEN_80433 : _GEN_80557; // @[FanCtrl.scala 518:68]
  wire [1:0] _GEN_80578 = _GEN_79248 == _GEN_79405 ? _GEN_80434 : _GEN_80558; // @[FanCtrl.scala 518:68]
  wire [1:0] _GEN_80579 = _GEN_79248 == _GEN_79405 ? _GEN_80435 : _GEN_80559; // @[FanCtrl.scala 518:68]
  wire [1:0] _GEN_80580 = _GEN_79248 == _GEN_79405 ? _GEN_80436 : _GEN_80560; // @[FanCtrl.scala 518:68]
  wire [1:0] _GEN_80581 = _GEN_79248 == _GEN_79405 ? _GEN_80437 : _GEN_80561; // @[FanCtrl.scala 518:68]
  wire [1:0] _GEN_80582 = _GEN_79248 == _GEN_79405 ? _GEN_80438 : _GEN_80562; // @[FanCtrl.scala 518:68]
  wire [1:0] _GEN_80603 = r_valid_1 ? _GEN_80563 : _GEN_80419; // @[FanCtrl.scala 517:33]
  wire [1:0] _GEN_80604 = r_valid_1 ? _GEN_80564 : _GEN_80420; // @[FanCtrl.scala 517:33]
  wire [1:0] _GEN_80605 = r_valid_1 ? _GEN_80565 : _GEN_80421; // @[FanCtrl.scala 517:33]
  wire [1:0] _GEN_80606 = r_valid_1 ? _GEN_80566 : _GEN_80422; // @[FanCtrl.scala 517:33]
  wire [1:0] _GEN_80607 = r_valid_1 ? _GEN_80567 : _GEN_80423; // @[FanCtrl.scala 517:33]
  wire [1:0] _GEN_80608 = r_valid_1 ? _GEN_80568 : _GEN_80424; // @[FanCtrl.scala 517:33]
  wire [1:0] _GEN_80609 = r_valid_1 ? _GEN_80569 : _GEN_80425; // @[FanCtrl.scala 517:33]
  wire [1:0] _GEN_80610 = r_valid_1 ? _GEN_80570 : _GEN_80426; // @[FanCtrl.scala 517:33]
  wire [1:0] _GEN_80611 = r_valid_1 ? _GEN_80571 : _GEN_80427; // @[FanCtrl.scala 517:33]
  wire [1:0] _GEN_80612 = r_valid_1 ? _GEN_80572 : _GEN_80428; // @[FanCtrl.scala 517:33]
  wire [1:0] _GEN_80613 = r_valid_1 ? _GEN_80573 : _GEN_80429; // @[FanCtrl.scala 517:33]
  wire [1:0] _GEN_80614 = r_valid_1 ? _GEN_80574 : _GEN_80430; // @[FanCtrl.scala 517:33]
  wire [1:0] _GEN_80615 = r_valid_1 ? _GEN_80575 : _GEN_80431; // @[FanCtrl.scala 517:33]
  wire [1:0] _GEN_80616 = r_valid_1 ? _GEN_80576 : _GEN_80432; // @[FanCtrl.scala 517:33]
  wire [1:0] _GEN_80617 = r_valid_1 ? _GEN_80577 : _GEN_80433; // @[FanCtrl.scala 517:33]
  wire [1:0] _GEN_80618 = r_valid_1 ? _GEN_80578 : _GEN_80434; // @[FanCtrl.scala 517:33]
  wire [1:0] _GEN_80619 = r_valid_1 ? _GEN_80579 : _GEN_80435; // @[FanCtrl.scala 517:33]
  wire [1:0] _GEN_80620 = r_valid_1 ? _GEN_80580 : _GEN_80436; // @[FanCtrl.scala 517:33]
  wire [1:0] _GEN_80621 = r_valid_1 ? _GEN_80581 : _GEN_80437; // @[FanCtrl.scala 517:33]
  wire [1:0] _GEN_80622 = r_valid_1 ? _GEN_80582 : _GEN_80438; // @[FanCtrl.scala 517:33]
  wire [3:0] _T_7966 = _T_7797 + 4'ha; // @[FanCtrl.scala 538:39]
  wire [1:0] _GEN_80687 = 4'h0 == _T_7966 ? 2'h2 : _GEN_80603; // @[FanCtrl.scala 538:{47,47}]
  wire [1:0] _GEN_80688 = 4'h1 == _T_7966 ? 2'h2 : _GEN_80604; // @[FanCtrl.scala 538:{47,47}]
  wire [1:0] _GEN_80689 = 4'h2 == _T_7966 ? 2'h2 : _GEN_80605; // @[FanCtrl.scala 538:{47,47}]
  wire [1:0] _GEN_80690 = 4'h3 == _T_7966 ? 2'h2 : _GEN_80606; // @[FanCtrl.scala 538:{47,47}]
  wire [1:0] _GEN_80691 = 4'h4 == _T_7966 ? 2'h2 : _GEN_80607; // @[FanCtrl.scala 538:{47,47}]
  wire [1:0] _GEN_80692 = 4'h5 == _T_7966 ? 2'h2 : _GEN_80608; // @[FanCtrl.scala 538:{47,47}]
  wire [1:0] _GEN_80693 = 4'h6 == _T_7966 ? 2'h2 : _GEN_80609; // @[FanCtrl.scala 538:{47,47}]
  wire [1:0] _GEN_80694 = 4'h7 == _T_7966 ? 2'h2 : _GEN_80610; // @[FanCtrl.scala 538:{47,47}]
  wire [1:0] _GEN_80695 = 4'h8 == _T_7966 ? 2'h2 : _GEN_80611; // @[FanCtrl.scala 538:{47,47}]
  wire [1:0] _GEN_80696 = 4'h9 == _T_7966 ? 2'h2 : _GEN_80612; // @[FanCtrl.scala 538:{47,47}]
  wire [1:0] _GEN_80697 = 4'ha == _T_7966 ? 2'h2 : _GEN_80613; // @[FanCtrl.scala 538:{47,47}]
  wire [1:0] _GEN_80698 = 4'hb == _T_7966 ? 2'h2 : _GEN_80614; // @[FanCtrl.scala 538:{47,47}]
  wire [1:0] _GEN_80699 = 4'hc == _T_7966 ? 2'h2 : _GEN_80615; // @[FanCtrl.scala 538:{47,47}]
  wire [1:0] _GEN_80700 = 4'hd == _T_7966 ? 2'h2 : _GEN_80616; // @[FanCtrl.scala 538:{47,47}]
  wire [1:0] _GEN_80701 = 4'he == _T_7966 ? 2'h2 : _GEN_80617; // @[FanCtrl.scala 538:{47,47}]
  wire [1:0] _GEN_80702 = 4'hf == _T_7966 ? 2'h2 : _GEN_80618; // @[FanCtrl.scala 538:{47,47}]
  wire [4:0] _GEN_97890 = {{1'd0}, _T_7966}; // @[FanCtrl.scala 538:{47,47}]
  wire [1:0] _GEN_80703 = 5'h10 == _GEN_97890 ? 2'h2 : _GEN_80619; // @[FanCtrl.scala 538:{47,47}]
  wire [1:0] _GEN_80704 = 5'h11 == _GEN_97890 ? 2'h2 : _GEN_80620; // @[FanCtrl.scala 538:{47,47}]
  wire [1:0] _GEN_80705 = 5'h12 == _GEN_97890 ? 2'h2 : _GEN_80621; // @[FanCtrl.scala 538:{47,47}]
  wire [1:0] _GEN_80706 = 5'h13 == _GEN_97890 ? 2'h2 : _GEN_80622; // @[FanCtrl.scala 538:{47,47}]
  wire [5:0] _T_7973 = _T_7801 + 6'ha; // @[FanCtrl.scala 540:65]
  wire [4:0] _GEN_80742 = 5'h3 == _T_7973[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 540:{45,45}]
  wire [4:0] _GEN_80743 = 5'h4 == _T_7973[4:0] ? w_vn_4 : _GEN_80742; // @[FanCtrl.scala 540:{45,45}]
  wire [4:0] _GEN_80744 = 5'h5 == _T_7973[4:0] ? 5'h0 : _GEN_80743; // @[FanCtrl.scala 540:{45,45}]
  wire [4:0] _GEN_80745 = 5'h6 == _T_7973[4:0] ? 5'h0 : _GEN_80744; // @[FanCtrl.scala 540:{45,45}]
  wire [4:0] _GEN_80746 = 5'h7 == _T_7973[4:0] ? w_vn_7 : _GEN_80745; // @[FanCtrl.scala 540:{45,45}]
  wire [4:0] _GEN_80747 = 5'h8 == _T_7973[4:0] ? w_vn_8 : _GEN_80746; // @[FanCtrl.scala 540:{45,45}]
  wire [4:0] _GEN_80748 = 5'h9 == _T_7973[4:0] ? 5'h0 : _GEN_80747; // @[FanCtrl.scala 540:{45,45}]
  wire [4:0] _GEN_80749 = 5'ha == _T_7973[4:0] ? 5'h0 : _GEN_80748; // @[FanCtrl.scala 540:{45,45}]
  wire [4:0] _GEN_80750 = 5'hb == _T_7973[4:0] ? w_vn_11 : _GEN_80749; // @[FanCtrl.scala 540:{45,45}]
  wire [4:0] _GEN_80751 = 5'hc == _T_7973[4:0] ? w_vn_12 : _GEN_80750; // @[FanCtrl.scala 540:{45,45}]
  wire [4:0] _GEN_80752 = 5'hd == _T_7973[4:0] ? w_vn_13 : _GEN_80751; // @[FanCtrl.scala 540:{45,45}]
  wire [4:0] _GEN_80753 = 5'he == _T_7973[4:0] ? 5'h0 : _GEN_80752; // @[FanCtrl.scala 540:{45,45}]
  wire [4:0] _GEN_80754 = 5'hf == _T_7973[4:0] ? w_vn_15 : _GEN_80753; // @[FanCtrl.scala 540:{45,45}]
  wire [4:0] _GEN_80755 = 5'h10 == _T_7973[4:0] ? w_vn_16 : _GEN_80754; // @[FanCtrl.scala 540:{45,45}]
  wire [4:0] _GEN_80756 = 5'h11 == _T_7973[4:0] ? 5'h0 : _GEN_80755; // @[FanCtrl.scala 540:{45,45}]
  wire [4:0] _GEN_80757 = 5'h12 == _T_7973[4:0] ? w_vn_18 : _GEN_80756; // @[FanCtrl.scala 540:{45,45}]
  wire [4:0] _GEN_80758 = 5'h13 == _T_7973[4:0] ? 5'h0 : _GEN_80757; // @[FanCtrl.scala 540:{45,45}]
  wire [4:0] _GEN_80759 = 5'h14 == _T_7973[4:0] ? 5'h0 : _GEN_80758; // @[FanCtrl.scala 540:{45,45}]
  wire [4:0] _GEN_80760 = 5'h15 == _T_7973[4:0] ? 5'h0 : _GEN_80759; // @[FanCtrl.scala 540:{45,45}]
  wire [4:0] _GEN_80761 = 5'h16 == _T_7973[4:0] ? 5'h0 : _GEN_80760; // @[FanCtrl.scala 540:{45,45}]
  wire [4:0] _GEN_80762 = 5'h17 == _T_7973[4:0] ? w_vn_23 : _GEN_80761; // @[FanCtrl.scala 540:{45,45}]
  wire [4:0] _GEN_80763 = 5'h18 == _T_7973[4:0] ? w_vn_24 : _GEN_80762; // @[FanCtrl.scala 540:{45,45}]
  wire [4:0] _GEN_80764 = 5'h19 == _T_7973[4:0] ? 5'h0 : _GEN_80763; // @[FanCtrl.scala 540:{45,45}]
  wire [4:0] _GEN_80765 = 5'h1a == _T_7973[4:0] ? 5'h0 : _GEN_80764; // @[FanCtrl.scala 540:{45,45}]
  wire [4:0] _GEN_80766 = 5'h1b == _T_7973[4:0] ? 5'h0 : _GEN_80765; // @[FanCtrl.scala 540:{45,45}]
  wire [4:0] _GEN_80767 = 5'h1c == _T_7973[4:0] ? 5'h0 : _GEN_80766; // @[FanCtrl.scala 540:{45,45}]
  wire [4:0] _GEN_80768 = 5'h1d == _T_7973[4:0] ? 5'h0 : _GEN_80767; // @[FanCtrl.scala 540:{45,45}]
  wire [4:0] _GEN_80769 = 5'h1e == _T_7973[4:0] ? 5'h0 : _GEN_80768; // @[FanCtrl.scala 540:{45,45}]
  wire [4:0] _GEN_80770 = 5'h1f == _T_7973[4:0] ? 5'h0 : _GEN_80769; // @[FanCtrl.scala 540:{45,45}]
  wire [1:0] _GEN_80771 = 4'h0 == _T_7966 ? 2'h1 : _GEN_80603; // @[FanCtrl.scala 542:{47,47}]
  wire [1:0] _GEN_80772 = 4'h1 == _T_7966 ? 2'h1 : _GEN_80604; // @[FanCtrl.scala 542:{47,47}]
  wire [1:0] _GEN_80773 = 4'h2 == _T_7966 ? 2'h1 : _GEN_80605; // @[FanCtrl.scala 542:{47,47}]
  wire [1:0] _GEN_80774 = 4'h3 == _T_7966 ? 2'h1 : _GEN_80606; // @[FanCtrl.scala 542:{47,47}]
  wire [1:0] _GEN_80775 = 4'h4 == _T_7966 ? 2'h1 : _GEN_80607; // @[FanCtrl.scala 542:{47,47}]
  wire [1:0] _GEN_80776 = 4'h5 == _T_7966 ? 2'h1 : _GEN_80608; // @[FanCtrl.scala 542:{47,47}]
  wire [1:0] _GEN_80777 = 4'h6 == _T_7966 ? 2'h1 : _GEN_80609; // @[FanCtrl.scala 542:{47,47}]
  wire [1:0] _GEN_80778 = 4'h7 == _T_7966 ? 2'h1 : _GEN_80610; // @[FanCtrl.scala 542:{47,47}]
  wire [1:0] _GEN_80779 = 4'h8 == _T_7966 ? 2'h1 : _GEN_80611; // @[FanCtrl.scala 542:{47,47}]
  wire [1:0] _GEN_80780 = 4'h9 == _T_7966 ? 2'h1 : _GEN_80612; // @[FanCtrl.scala 542:{47,47}]
  wire [1:0] _GEN_80781 = 4'ha == _T_7966 ? 2'h1 : _GEN_80613; // @[FanCtrl.scala 542:{47,47}]
  wire [1:0] _GEN_80782 = 4'hb == _T_7966 ? 2'h1 : _GEN_80614; // @[FanCtrl.scala 542:{47,47}]
  wire [1:0] _GEN_80783 = 4'hc == _T_7966 ? 2'h1 : _GEN_80615; // @[FanCtrl.scala 542:{47,47}]
  wire [1:0] _GEN_80784 = 4'hd == _T_7966 ? 2'h1 : _GEN_80616; // @[FanCtrl.scala 542:{47,47}]
  wire [1:0] _GEN_80785 = 4'he == _T_7966 ? 2'h1 : _GEN_80617; // @[FanCtrl.scala 542:{47,47}]
  wire [1:0] _GEN_80786 = 4'hf == _T_7966 ? 2'h1 : _GEN_80618; // @[FanCtrl.scala 542:{47,47}]
  wire [1:0] _GEN_80787 = 5'h10 == _GEN_97890 ? 2'h1 : _GEN_80619; // @[FanCtrl.scala 542:{47,47}]
  wire [1:0] _GEN_80788 = 5'h11 == _GEN_97890 ? 2'h1 : _GEN_80620; // @[FanCtrl.scala 542:{47,47}]
  wire [1:0] _GEN_80789 = 5'h12 == _GEN_97890 ? 2'h1 : _GEN_80621; // @[FanCtrl.scala 542:{47,47}]
  wire [1:0] _GEN_80790 = 5'h13 == _GEN_97890 ? 2'h1 : _GEN_80622; // @[FanCtrl.scala 542:{47,47}]
  wire [1:0] _GEN_80791 = 4'h0 == _T_7966 ? 2'h0 : _GEN_80603; // @[FanCtrl.scala 545:{47,47}]
  wire [1:0] _GEN_80792 = 4'h1 == _T_7966 ? 2'h0 : _GEN_80604; // @[FanCtrl.scala 545:{47,47}]
  wire [1:0] _GEN_80793 = 4'h2 == _T_7966 ? 2'h0 : _GEN_80605; // @[FanCtrl.scala 545:{47,47}]
  wire [1:0] _GEN_80794 = 4'h3 == _T_7966 ? 2'h0 : _GEN_80606; // @[FanCtrl.scala 545:{47,47}]
  wire [1:0] _GEN_80795 = 4'h4 == _T_7966 ? 2'h0 : _GEN_80607; // @[FanCtrl.scala 545:{47,47}]
  wire [1:0] _GEN_80796 = 4'h5 == _T_7966 ? 2'h0 : _GEN_80608; // @[FanCtrl.scala 545:{47,47}]
  wire [1:0] _GEN_80797 = 4'h6 == _T_7966 ? 2'h0 : _GEN_80609; // @[FanCtrl.scala 545:{47,47}]
  wire [1:0] _GEN_80798 = 4'h7 == _T_7966 ? 2'h0 : _GEN_80610; // @[FanCtrl.scala 545:{47,47}]
  wire [1:0] _GEN_80799 = 4'h8 == _T_7966 ? 2'h0 : _GEN_80611; // @[FanCtrl.scala 545:{47,47}]
  wire [1:0] _GEN_80800 = 4'h9 == _T_7966 ? 2'h0 : _GEN_80612; // @[FanCtrl.scala 545:{47,47}]
  wire [1:0] _GEN_80801 = 4'ha == _T_7966 ? 2'h0 : _GEN_80613; // @[FanCtrl.scala 545:{47,47}]
  wire [1:0] _GEN_80802 = 4'hb == _T_7966 ? 2'h0 : _GEN_80614; // @[FanCtrl.scala 545:{47,47}]
  wire [1:0] _GEN_80803 = 4'hc == _T_7966 ? 2'h0 : _GEN_80615; // @[FanCtrl.scala 545:{47,47}]
  wire [1:0] _GEN_80804 = 4'hd == _T_7966 ? 2'h0 : _GEN_80616; // @[FanCtrl.scala 545:{47,47}]
  wire [1:0] _GEN_80805 = 4'he == _T_7966 ? 2'h0 : _GEN_80617; // @[FanCtrl.scala 545:{47,47}]
  wire [1:0] _GEN_80806 = 4'hf == _T_7966 ? 2'h0 : _GEN_80618; // @[FanCtrl.scala 545:{47,47}]
  wire [1:0] _GEN_80807 = 5'h10 == _GEN_97890 ? 2'h0 : _GEN_80619; // @[FanCtrl.scala 545:{47,47}]
  wire [1:0] _GEN_80808 = 5'h11 == _GEN_97890 ? 2'h0 : _GEN_80620; // @[FanCtrl.scala 545:{47,47}]
  wire [1:0] _GEN_80809 = 5'h12 == _GEN_97890 ? 2'h0 : _GEN_80621; // @[FanCtrl.scala 545:{47,47}]
  wire [1:0] _GEN_80810 = 5'h13 == _GEN_97890 ? 2'h0 : _GEN_80622; // @[FanCtrl.scala 545:{47,47}]
  wire [1:0] _GEN_80811 = _GEN_79280 == _GEN_80770 ? _GEN_80771 : _GEN_80791; // @[FanCtrl.scala 540:74]
  wire [1:0] _GEN_80812 = _GEN_79280 == _GEN_80770 ? _GEN_80772 : _GEN_80792; // @[FanCtrl.scala 540:74]
  wire [1:0] _GEN_80813 = _GEN_79280 == _GEN_80770 ? _GEN_80773 : _GEN_80793; // @[FanCtrl.scala 540:74]
  wire [1:0] _GEN_80814 = _GEN_79280 == _GEN_80770 ? _GEN_80774 : _GEN_80794; // @[FanCtrl.scala 540:74]
  wire [1:0] _GEN_80815 = _GEN_79280 == _GEN_80770 ? _GEN_80775 : _GEN_80795; // @[FanCtrl.scala 540:74]
  wire [1:0] _GEN_80816 = _GEN_79280 == _GEN_80770 ? _GEN_80776 : _GEN_80796; // @[FanCtrl.scala 540:74]
  wire [1:0] _GEN_80817 = _GEN_79280 == _GEN_80770 ? _GEN_80777 : _GEN_80797; // @[FanCtrl.scala 540:74]
  wire [1:0] _GEN_80818 = _GEN_79280 == _GEN_80770 ? _GEN_80778 : _GEN_80798; // @[FanCtrl.scala 540:74]
  wire [1:0] _GEN_80819 = _GEN_79280 == _GEN_80770 ? _GEN_80779 : _GEN_80799; // @[FanCtrl.scala 540:74]
  wire [1:0] _GEN_80820 = _GEN_79280 == _GEN_80770 ? _GEN_80780 : _GEN_80800; // @[FanCtrl.scala 540:74]
  wire [1:0] _GEN_80821 = _GEN_79280 == _GEN_80770 ? _GEN_80781 : _GEN_80801; // @[FanCtrl.scala 540:74]
  wire [1:0] _GEN_80822 = _GEN_79280 == _GEN_80770 ? _GEN_80782 : _GEN_80802; // @[FanCtrl.scala 540:74]
  wire [1:0] _GEN_80823 = _GEN_79280 == _GEN_80770 ? _GEN_80783 : _GEN_80803; // @[FanCtrl.scala 540:74]
  wire [1:0] _GEN_80824 = _GEN_79280 == _GEN_80770 ? _GEN_80784 : _GEN_80804; // @[FanCtrl.scala 540:74]
  wire [1:0] _GEN_80825 = _GEN_79280 == _GEN_80770 ? _GEN_80785 : _GEN_80805; // @[FanCtrl.scala 540:74]
  wire [1:0] _GEN_80826 = _GEN_79280 == _GEN_80770 ? _GEN_80786 : _GEN_80806; // @[FanCtrl.scala 540:74]
  wire [1:0] _GEN_80827 = _GEN_79280 == _GEN_80770 ? _GEN_80787 : _GEN_80807; // @[FanCtrl.scala 540:74]
  wire [1:0] _GEN_80828 = _GEN_79280 == _GEN_80770 ? _GEN_80788 : _GEN_80808; // @[FanCtrl.scala 540:74]
  wire [1:0] _GEN_80829 = _GEN_79280 == _GEN_80770 ? _GEN_80789 : _GEN_80809; // @[FanCtrl.scala 540:74]
  wire [1:0] _GEN_80830 = _GEN_79280 == _GEN_80770 ? _GEN_80790 : _GEN_80810; // @[FanCtrl.scala 540:74]
  wire [1:0] _GEN_80831 = _GEN_79280 == _GEN_79501 ? _GEN_80687 : _GEN_80811; // @[FanCtrl.scala 536:69]
  wire [1:0] _GEN_80832 = _GEN_79280 == _GEN_79501 ? _GEN_80688 : _GEN_80812; // @[FanCtrl.scala 536:69]
  wire [1:0] _GEN_80833 = _GEN_79280 == _GEN_79501 ? _GEN_80689 : _GEN_80813; // @[FanCtrl.scala 536:69]
  wire [1:0] _GEN_80834 = _GEN_79280 == _GEN_79501 ? _GEN_80690 : _GEN_80814; // @[FanCtrl.scala 536:69]
  wire [1:0] _GEN_80835 = _GEN_79280 == _GEN_79501 ? _GEN_80691 : _GEN_80815; // @[FanCtrl.scala 536:69]
  wire [1:0] _GEN_80836 = _GEN_79280 == _GEN_79501 ? _GEN_80692 : _GEN_80816; // @[FanCtrl.scala 536:69]
  wire [1:0] _GEN_80837 = _GEN_79280 == _GEN_79501 ? _GEN_80693 : _GEN_80817; // @[FanCtrl.scala 536:69]
  wire [1:0] _GEN_80838 = _GEN_79280 == _GEN_79501 ? _GEN_80694 : _GEN_80818; // @[FanCtrl.scala 536:69]
  wire [1:0] _GEN_80839 = _GEN_79280 == _GEN_79501 ? _GEN_80695 : _GEN_80819; // @[FanCtrl.scala 536:69]
  wire [1:0] _GEN_80840 = _GEN_79280 == _GEN_79501 ? _GEN_80696 : _GEN_80820; // @[FanCtrl.scala 536:69]
  wire [1:0] _GEN_80841 = _GEN_79280 == _GEN_79501 ? _GEN_80697 : _GEN_80821; // @[FanCtrl.scala 536:69]
  wire [1:0] _GEN_80842 = _GEN_79280 == _GEN_79501 ? _GEN_80698 : _GEN_80822; // @[FanCtrl.scala 536:69]
  wire [1:0] _GEN_80843 = _GEN_79280 == _GEN_79501 ? _GEN_80699 : _GEN_80823; // @[FanCtrl.scala 536:69]
  wire [1:0] _GEN_80844 = _GEN_79280 == _GEN_79501 ? _GEN_80700 : _GEN_80824; // @[FanCtrl.scala 536:69]
  wire [1:0] _GEN_80845 = _GEN_79280 == _GEN_79501 ? _GEN_80701 : _GEN_80825; // @[FanCtrl.scala 536:69]
  wire [1:0] _GEN_80846 = _GEN_79280 == _GEN_79501 ? _GEN_80702 : _GEN_80826; // @[FanCtrl.scala 536:69]
  wire [1:0] _GEN_80847 = _GEN_79280 == _GEN_79501 ? _GEN_80703 : _GEN_80827; // @[FanCtrl.scala 536:69]
  wire [1:0] _GEN_80848 = _GEN_79280 == _GEN_79501 ? _GEN_80704 : _GEN_80828; // @[FanCtrl.scala 536:69]
  wire [1:0] _GEN_80849 = _GEN_79280 == _GEN_79501 ? _GEN_80705 : _GEN_80829; // @[FanCtrl.scala 536:69]
  wire [1:0] _GEN_80850 = _GEN_79280 == _GEN_79501 ? _GEN_80706 : _GEN_80830; // @[FanCtrl.scala 536:69]
  wire [1:0] _GEN_80851 = 4'h0 == _T_7799 ? 2'h0 : _GEN_80603; // @[FanCtrl.scala 548:{44,44}]
  wire [1:0] _GEN_80852 = 4'h1 == _T_7799 ? 2'h0 : _GEN_80604; // @[FanCtrl.scala 548:{44,44}]
  wire [1:0] _GEN_80853 = 4'h2 == _T_7799 ? 2'h0 : _GEN_80605; // @[FanCtrl.scala 548:{44,44}]
  wire [1:0] _GEN_80854 = 4'h3 == _T_7799 ? 2'h0 : _GEN_80606; // @[FanCtrl.scala 548:{44,44}]
  wire [1:0] _GEN_80855 = 4'h4 == _T_7799 ? 2'h0 : _GEN_80607; // @[FanCtrl.scala 548:{44,44}]
  wire [1:0] _GEN_80856 = 4'h5 == _T_7799 ? 2'h0 : _GEN_80608; // @[FanCtrl.scala 548:{44,44}]
  wire [1:0] _GEN_80857 = 4'h6 == _T_7799 ? 2'h0 : _GEN_80609; // @[FanCtrl.scala 548:{44,44}]
  wire [1:0] _GEN_80858 = 4'h7 == _T_7799 ? 2'h0 : _GEN_80610; // @[FanCtrl.scala 548:{44,44}]
  wire [1:0] _GEN_80859 = 4'h8 == _T_7799 ? 2'h0 : _GEN_80611; // @[FanCtrl.scala 548:{44,44}]
  wire [1:0] _GEN_80860 = 4'h9 == _T_7799 ? 2'h0 : _GEN_80612; // @[FanCtrl.scala 548:{44,44}]
  wire [1:0] _GEN_80861 = 4'ha == _T_7799 ? 2'h0 : _GEN_80613; // @[FanCtrl.scala 548:{44,44}]
  wire [1:0] _GEN_80862 = 4'hb == _T_7799 ? 2'h0 : _GEN_80614; // @[FanCtrl.scala 548:{44,44}]
  wire [1:0] _GEN_80863 = 4'hc == _T_7799 ? 2'h0 : _GEN_80615; // @[FanCtrl.scala 548:{44,44}]
  wire [1:0] _GEN_80864 = 4'hd == _T_7799 ? 2'h0 : _GEN_80616; // @[FanCtrl.scala 548:{44,44}]
  wire [1:0] _GEN_80865 = 4'he == _T_7799 ? 2'h0 : _GEN_80617; // @[FanCtrl.scala 548:{44,44}]
  wire [1:0] _GEN_80866 = 4'hf == _T_7799 ? 2'h0 : _GEN_80618; // @[FanCtrl.scala 548:{44,44}]
  wire [1:0] _GEN_80867 = 5'h10 == _GEN_97870 ? 2'h0 : _GEN_80619; // @[FanCtrl.scala 548:{44,44}]
  wire [1:0] _GEN_80868 = 5'h11 == _GEN_97870 ? 2'h0 : _GEN_80620; // @[FanCtrl.scala 548:{44,44}]
  wire [1:0] _GEN_80869 = 5'h12 == _GEN_97870 ? 2'h0 : _GEN_80621; // @[FanCtrl.scala 548:{44,44}]
  wire [1:0] _GEN_80870 = 5'h13 == _GEN_97870 ? 2'h0 : _GEN_80622; // @[FanCtrl.scala 548:{44,44}]
  wire [1:0] _GEN_80871 = r_valid_1 ? _GEN_80831 : _GEN_80851; // @[FanCtrl.scala 535:33]
  wire [1:0] _GEN_80872 = r_valid_1 ? _GEN_80832 : _GEN_80852; // @[FanCtrl.scala 535:33]
  wire [1:0] _GEN_80873 = r_valid_1 ? _GEN_80833 : _GEN_80853; // @[FanCtrl.scala 535:33]
  wire [1:0] _GEN_80874 = r_valid_1 ? _GEN_80834 : _GEN_80854; // @[FanCtrl.scala 535:33]
  wire [1:0] _GEN_80875 = r_valid_1 ? _GEN_80835 : _GEN_80855; // @[FanCtrl.scala 535:33]
  wire [1:0] _GEN_80876 = r_valid_1 ? _GEN_80836 : _GEN_80856; // @[FanCtrl.scala 535:33]
  wire [1:0] _GEN_80877 = r_valid_1 ? _GEN_80837 : _GEN_80857; // @[FanCtrl.scala 535:33]
  wire [1:0] _GEN_80878 = r_valid_1 ? _GEN_80838 : _GEN_80858; // @[FanCtrl.scala 535:33]
  wire [1:0] _GEN_80879 = r_valid_1 ? _GEN_80839 : _GEN_80859; // @[FanCtrl.scala 535:33]
  wire [1:0] _GEN_80880 = r_valid_1 ? _GEN_80840 : _GEN_80860; // @[FanCtrl.scala 535:33]
  wire [1:0] _GEN_80881 = r_valid_1 ? _GEN_80841 : _GEN_80861; // @[FanCtrl.scala 535:33]
  wire [1:0] _GEN_80882 = r_valid_1 ? _GEN_80842 : _GEN_80862; // @[FanCtrl.scala 535:33]
  wire [1:0] _GEN_80883 = r_valid_1 ? _GEN_80843 : _GEN_80863; // @[FanCtrl.scala 535:33]
  wire [1:0] _GEN_80884 = r_valid_1 ? _GEN_80844 : _GEN_80864; // @[FanCtrl.scala 535:33]
  wire [1:0] _GEN_80885 = r_valid_1 ? _GEN_80845 : _GEN_80865; // @[FanCtrl.scala 535:33]
  wire [1:0] _GEN_80886 = r_valid_1 ? _GEN_80846 : _GEN_80866; // @[FanCtrl.scala 535:33]
  wire [1:0] _GEN_80887 = r_valid_1 ? _GEN_80847 : _GEN_80867; // @[FanCtrl.scala 535:33]
  wire [1:0] _GEN_80888 = r_valid_1 ? _GEN_80848 : _GEN_80868; // @[FanCtrl.scala 535:33]
  wire [1:0] _GEN_80889 = r_valid_1 ? _GEN_80849 : _GEN_80869; // @[FanCtrl.scala 535:33]
  wire [1:0] _GEN_80890 = r_valid_1 ? _GEN_80850 : _GEN_80870; // @[FanCtrl.scala 535:33]
  wire [3:0] _T_8395 = 1'h1 * 3'h4; // @[FanCtrl.scala 479:28]
  wire [3:0] _T_8397 = _T_8395 + 4'h8; // @[FanCtrl.scala 479:35]
  wire [1:0] _GEN_84757 = 4'h0 == _T_8397 ? 2'h0 : _GEN_80871; // @[FanCtrl.scala 479:{42,42}]
  wire [1:0] _GEN_84758 = 4'h1 == _T_8397 ? 2'h0 : _GEN_80872; // @[FanCtrl.scala 479:{42,42}]
  wire [1:0] _GEN_84759 = 4'h2 == _T_8397 ? 2'h0 : _GEN_80873; // @[FanCtrl.scala 479:{42,42}]
  wire [1:0] _GEN_84760 = 4'h3 == _T_8397 ? 2'h0 : _GEN_80874; // @[FanCtrl.scala 479:{42,42}]
  wire [1:0] _GEN_84761 = 4'h4 == _T_8397 ? 2'h0 : _GEN_80875; // @[FanCtrl.scala 479:{42,42}]
  wire [1:0] _GEN_84762 = 4'h5 == _T_8397 ? 2'h0 : _GEN_80876; // @[FanCtrl.scala 479:{42,42}]
  wire [1:0] _GEN_84763 = 4'h6 == _T_8397 ? 2'h0 : _GEN_80877; // @[FanCtrl.scala 479:{42,42}]
  wire [1:0] _GEN_84764 = 4'h7 == _T_8397 ? 2'h0 : _GEN_80878; // @[FanCtrl.scala 479:{42,42}]
  wire [1:0] _GEN_84765 = 4'h8 == _T_8397 ? 2'h0 : _GEN_80879; // @[FanCtrl.scala 479:{42,42}]
  wire [1:0] _GEN_84766 = 4'h9 == _T_8397 ? 2'h0 : _GEN_80880; // @[FanCtrl.scala 479:{42,42}]
  wire [1:0] _GEN_84767 = 4'ha == _T_8397 ? 2'h0 : _GEN_80881; // @[FanCtrl.scala 479:{42,42}]
  wire [1:0] _GEN_84768 = 4'hb == _T_8397 ? 2'h0 : _GEN_80882; // @[FanCtrl.scala 479:{42,42}]
  wire [1:0] _GEN_84769 = 4'hc == _T_8397 ? 2'h0 : _GEN_80883; // @[FanCtrl.scala 479:{42,42}]
  wire [1:0] _GEN_84770 = 4'hd == _T_8397 ? 2'h0 : _GEN_80884; // @[FanCtrl.scala 479:{42,42}]
  wire [1:0] _GEN_84771 = 4'he == _T_8397 ? 2'h0 : _GEN_80885; // @[FanCtrl.scala 479:{42,42}]
  wire [1:0] _GEN_84772 = 4'hf == _T_8397 ? 2'h0 : _GEN_80886; // @[FanCtrl.scala 479:{42,42}]
  wire [4:0] _GEN_97978 = {{1'd0}, _T_8397}; // @[FanCtrl.scala 479:{42,42}]
  wire [1:0] _GEN_84773 = 5'h10 == _GEN_97978 ? 2'h0 : _GEN_80887; // @[FanCtrl.scala 479:{42,42}]
  wire [1:0] _GEN_84774 = 5'h11 == _GEN_97978 ? 2'h0 : _GEN_80888; // @[FanCtrl.scala 479:{42,42}]
  wire [1:0] _GEN_84775 = 5'h12 == _GEN_97978 ? 2'h0 : _GEN_80889; // @[FanCtrl.scala 479:{42,42}]
  wire [1:0] _GEN_84776 = 5'h13 == _GEN_97978 ? 2'h0 : _GEN_80890; // @[FanCtrl.scala 479:{42,42}]
  wire [5:0] _T_8399 = 5'h10 * 1'h1; // @[FanCtrl.scala 483:25]
  wire [5:0] _T_8401 = _T_8399 + 6'h7; // @[FanCtrl.scala 483:31]
  wire [5:0] _T_8405 = _T_8399 + 6'h8; // @[FanCtrl.scala 483:59]
  wire [4:0] _GEN_84780 = 5'h3 == _T_8401[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_84781 = 5'h4 == _T_8401[4:0] ? w_vn_4 : _GEN_84780; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_84782 = 5'h5 == _T_8401[4:0] ? 5'h0 : _GEN_84781; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_84783 = 5'h6 == _T_8401[4:0] ? 5'h0 : _GEN_84782; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_84784 = 5'h7 == _T_8401[4:0] ? w_vn_7 : _GEN_84783; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_84785 = 5'h8 == _T_8401[4:0] ? w_vn_8 : _GEN_84784; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_84786 = 5'h9 == _T_8401[4:0] ? 5'h0 : _GEN_84785; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_84787 = 5'ha == _T_8401[4:0] ? 5'h0 : _GEN_84786; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_84788 = 5'hb == _T_8401[4:0] ? w_vn_11 : _GEN_84787; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_84789 = 5'hc == _T_8401[4:0] ? w_vn_12 : _GEN_84788; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_84790 = 5'hd == _T_8401[4:0] ? w_vn_13 : _GEN_84789; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_84791 = 5'he == _T_8401[4:0] ? 5'h0 : _GEN_84790; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_84792 = 5'hf == _T_8401[4:0] ? w_vn_15 : _GEN_84791; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_84793 = 5'h10 == _T_8401[4:0] ? w_vn_16 : _GEN_84792; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_84794 = 5'h11 == _T_8401[4:0] ? 5'h0 : _GEN_84793; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_84795 = 5'h12 == _T_8401[4:0] ? w_vn_18 : _GEN_84794; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_84796 = 5'h13 == _T_8401[4:0] ? 5'h0 : _GEN_84795; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_84797 = 5'h14 == _T_8401[4:0] ? 5'h0 : _GEN_84796; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_84798 = 5'h15 == _T_8401[4:0] ? 5'h0 : _GEN_84797; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_84799 = 5'h16 == _T_8401[4:0] ? 5'h0 : _GEN_84798; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_84800 = 5'h17 == _T_8401[4:0] ? w_vn_23 : _GEN_84799; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_84801 = 5'h18 == _T_8401[4:0] ? w_vn_24 : _GEN_84800; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_84802 = 5'h19 == _T_8401[4:0] ? 5'h0 : _GEN_84801; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_84803 = 5'h1a == _T_8401[4:0] ? 5'h0 : _GEN_84802; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_84804 = 5'h1b == _T_8401[4:0] ? 5'h0 : _GEN_84803; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_84805 = 5'h1c == _T_8401[4:0] ? 5'h0 : _GEN_84804; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_84806 = 5'h1d == _T_8401[4:0] ? 5'h0 : _GEN_84805; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_84807 = 5'h1e == _T_8401[4:0] ? 5'h0 : _GEN_84806; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_84808 = 5'h1f == _T_8401[4:0] ? 5'h0 : _GEN_84807; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_84812 = 5'h3 == _T_8405[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_84813 = 5'h4 == _T_8405[4:0] ? w_vn_4 : _GEN_84812; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_84814 = 5'h5 == _T_8405[4:0] ? 5'h0 : _GEN_84813; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_84815 = 5'h6 == _T_8405[4:0] ? 5'h0 : _GEN_84814; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_84816 = 5'h7 == _T_8405[4:0] ? w_vn_7 : _GEN_84815; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_84817 = 5'h8 == _T_8405[4:0] ? w_vn_8 : _GEN_84816; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_84818 = 5'h9 == _T_8405[4:0] ? 5'h0 : _GEN_84817; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_84819 = 5'ha == _T_8405[4:0] ? 5'h0 : _GEN_84818; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_84820 = 5'hb == _T_8405[4:0] ? w_vn_11 : _GEN_84819; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_84821 = 5'hc == _T_8405[4:0] ? w_vn_12 : _GEN_84820; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_84822 = 5'hd == _T_8405[4:0] ? w_vn_13 : _GEN_84821; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_84823 = 5'he == _T_8405[4:0] ? 5'h0 : _GEN_84822; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_84824 = 5'hf == _T_8405[4:0] ? w_vn_15 : _GEN_84823; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_84825 = 5'h10 == _T_8405[4:0] ? w_vn_16 : _GEN_84824; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_84826 = 5'h11 == _T_8405[4:0] ? 5'h0 : _GEN_84825; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_84827 = 5'h12 == _T_8405[4:0] ? w_vn_18 : _GEN_84826; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_84828 = 5'h13 == _T_8405[4:0] ? 5'h0 : _GEN_84827; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_84829 = 5'h14 == _T_8405[4:0] ? 5'h0 : _GEN_84828; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_84830 = 5'h15 == _T_8405[4:0] ? 5'h0 : _GEN_84829; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_84831 = 5'h16 == _T_8405[4:0] ? 5'h0 : _GEN_84830; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_84832 = 5'h17 == _T_8405[4:0] ? w_vn_23 : _GEN_84831; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_84833 = 5'h18 == _T_8405[4:0] ? w_vn_24 : _GEN_84832; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_84834 = 5'h19 == _T_8405[4:0] ? 5'h0 : _GEN_84833; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_84835 = 5'h1a == _T_8405[4:0] ? 5'h0 : _GEN_84834; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_84836 = 5'h1b == _T_8405[4:0] ? 5'h0 : _GEN_84835; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_84837 = 5'h1c == _T_8405[4:0] ? 5'h0 : _GEN_84836; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_84838 = 5'h1d == _T_8405[4:0] ? 5'h0 : _GEN_84837; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_84839 = 5'h1e == _T_8405[4:0] ? 5'h0 : _GEN_84838; // @[FanCtrl.scala 483:{39,39}]
  wire [4:0] _GEN_84840 = 5'h1f == _T_8405[4:0] ? 5'h0 : _GEN_84839; // @[FanCtrl.scala 483:{39,39}]
  wire  _T_8407 = _GEN_84808 == _GEN_84840; // @[FanCtrl.scala 483:39]
  wire [5:0] _T_8414 = _T_8399 + 6'h3; // @[FanCtrl.scala 489:31]
  wire [5:0] _T_8418 = _T_8399 + 6'h4; // @[FanCtrl.scala 489:59]
  wire [4:0] _GEN_84937 = 5'h3 == _T_8414[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_84938 = 5'h4 == _T_8414[4:0] ? w_vn_4 : _GEN_84937; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_84939 = 5'h5 == _T_8414[4:0] ? 5'h0 : _GEN_84938; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_84940 = 5'h6 == _T_8414[4:0] ? 5'h0 : _GEN_84939; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_84941 = 5'h7 == _T_8414[4:0] ? w_vn_7 : _GEN_84940; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_84942 = 5'h8 == _T_8414[4:0] ? w_vn_8 : _GEN_84941; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_84943 = 5'h9 == _T_8414[4:0] ? 5'h0 : _GEN_84942; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_84944 = 5'ha == _T_8414[4:0] ? 5'h0 : _GEN_84943; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_84945 = 5'hb == _T_8414[4:0] ? w_vn_11 : _GEN_84944; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_84946 = 5'hc == _T_8414[4:0] ? w_vn_12 : _GEN_84945; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_84947 = 5'hd == _T_8414[4:0] ? w_vn_13 : _GEN_84946; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_84948 = 5'he == _T_8414[4:0] ? 5'h0 : _GEN_84947; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_84949 = 5'hf == _T_8414[4:0] ? w_vn_15 : _GEN_84948; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_84950 = 5'h10 == _T_8414[4:0] ? w_vn_16 : _GEN_84949; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_84951 = 5'h11 == _T_8414[4:0] ? 5'h0 : _GEN_84950; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_84952 = 5'h12 == _T_8414[4:0] ? w_vn_18 : _GEN_84951; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_84953 = 5'h13 == _T_8414[4:0] ? 5'h0 : _GEN_84952; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_84954 = 5'h14 == _T_8414[4:0] ? 5'h0 : _GEN_84953; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_84955 = 5'h15 == _T_8414[4:0] ? 5'h0 : _GEN_84954; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_84956 = 5'h16 == _T_8414[4:0] ? 5'h0 : _GEN_84955; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_84957 = 5'h17 == _T_8414[4:0] ? w_vn_23 : _GEN_84956; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_84958 = 5'h18 == _T_8414[4:0] ? w_vn_24 : _GEN_84957; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_84959 = 5'h19 == _T_8414[4:0] ? 5'h0 : _GEN_84958; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_84960 = 5'h1a == _T_8414[4:0] ? 5'h0 : _GEN_84959; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_84961 = 5'h1b == _T_8414[4:0] ? 5'h0 : _GEN_84960; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_84962 = 5'h1c == _T_8414[4:0] ? 5'h0 : _GEN_84961; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_84963 = 5'h1d == _T_8414[4:0] ? 5'h0 : _GEN_84962; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_84964 = 5'h1e == _T_8414[4:0] ? 5'h0 : _GEN_84963; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_84965 = 5'h1f == _T_8414[4:0] ? 5'h0 : _GEN_84964; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_84969 = 5'h3 == _T_8418[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_84970 = 5'h4 == _T_8418[4:0] ? w_vn_4 : _GEN_84969; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_84971 = 5'h5 == _T_8418[4:0] ? 5'h0 : _GEN_84970; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_84972 = 5'h6 == _T_8418[4:0] ? 5'h0 : _GEN_84971; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_84973 = 5'h7 == _T_8418[4:0] ? w_vn_7 : _GEN_84972; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_84974 = 5'h8 == _T_8418[4:0] ? w_vn_8 : _GEN_84973; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_84975 = 5'h9 == _T_8418[4:0] ? 5'h0 : _GEN_84974; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_84976 = 5'ha == _T_8418[4:0] ? 5'h0 : _GEN_84975; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_84977 = 5'hb == _T_8418[4:0] ? w_vn_11 : _GEN_84976; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_84978 = 5'hc == _T_8418[4:0] ? w_vn_12 : _GEN_84977; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_84979 = 5'hd == _T_8418[4:0] ? w_vn_13 : _GEN_84978; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_84980 = 5'he == _T_8418[4:0] ? 5'h0 : _GEN_84979; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_84981 = 5'hf == _T_8418[4:0] ? w_vn_15 : _GEN_84980; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_84982 = 5'h10 == _T_8418[4:0] ? w_vn_16 : _GEN_84981; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_84983 = 5'h11 == _T_8418[4:0] ? 5'h0 : _GEN_84982; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_84984 = 5'h12 == _T_8418[4:0] ? w_vn_18 : _GEN_84983; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_84985 = 5'h13 == _T_8418[4:0] ? 5'h0 : _GEN_84984; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_84986 = 5'h14 == _T_8418[4:0] ? 5'h0 : _GEN_84985; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_84987 = 5'h15 == _T_8418[4:0] ? 5'h0 : _GEN_84986; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_84988 = 5'h16 == _T_8418[4:0] ? 5'h0 : _GEN_84987; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_84989 = 5'h17 == _T_8418[4:0] ? w_vn_23 : _GEN_84988; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_84990 = 5'h18 == _T_8418[4:0] ? w_vn_24 : _GEN_84989; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_84991 = 5'h19 == _T_8418[4:0] ? 5'h0 : _GEN_84990; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_84992 = 5'h1a == _T_8418[4:0] ? 5'h0 : _GEN_84991; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_84993 = 5'h1b == _T_8418[4:0] ? 5'h0 : _GEN_84992; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_84994 = 5'h1c == _T_8418[4:0] ? 5'h0 : _GEN_84993; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_84995 = 5'h1d == _T_8418[4:0] ? 5'h0 : _GEN_84994; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_84996 = 5'h1e == _T_8418[4:0] ? 5'h0 : _GEN_84995; // @[FanCtrl.scala 489:{38,38}]
  wire [4:0] _GEN_84997 = 5'h1f == _T_8418[4:0] ? 5'h0 : _GEN_84996; // @[FanCtrl.scala 489:{38,38}]
  wire  _T_8420 = _GEN_84965 == _GEN_84997; // @[FanCtrl.scala 489:38]
  wire [5:0] _T_8423 = _T_8399 + 6'hb; // @[FanCtrl.scala 490:32]
  wire [5:0] _T_8427 = _T_8399 + 6'hc; // @[FanCtrl.scala 490:61]
  wire [4:0] _GEN_85001 = 5'h3 == _T_8423[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_85002 = 5'h4 == _T_8423[4:0] ? w_vn_4 : _GEN_85001; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_85003 = 5'h5 == _T_8423[4:0] ? 5'h0 : _GEN_85002; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_85004 = 5'h6 == _T_8423[4:0] ? 5'h0 : _GEN_85003; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_85005 = 5'h7 == _T_8423[4:0] ? w_vn_7 : _GEN_85004; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_85006 = 5'h8 == _T_8423[4:0] ? w_vn_8 : _GEN_85005; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_85007 = 5'h9 == _T_8423[4:0] ? 5'h0 : _GEN_85006; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_85008 = 5'ha == _T_8423[4:0] ? 5'h0 : _GEN_85007; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_85009 = 5'hb == _T_8423[4:0] ? w_vn_11 : _GEN_85008; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_85010 = 5'hc == _T_8423[4:0] ? w_vn_12 : _GEN_85009; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_85011 = 5'hd == _T_8423[4:0] ? w_vn_13 : _GEN_85010; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_85012 = 5'he == _T_8423[4:0] ? 5'h0 : _GEN_85011; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_85013 = 5'hf == _T_8423[4:0] ? w_vn_15 : _GEN_85012; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_85014 = 5'h10 == _T_8423[4:0] ? w_vn_16 : _GEN_85013; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_85015 = 5'h11 == _T_8423[4:0] ? 5'h0 : _GEN_85014; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_85016 = 5'h12 == _T_8423[4:0] ? w_vn_18 : _GEN_85015; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_85017 = 5'h13 == _T_8423[4:0] ? 5'h0 : _GEN_85016; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_85018 = 5'h14 == _T_8423[4:0] ? 5'h0 : _GEN_85017; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_85019 = 5'h15 == _T_8423[4:0] ? 5'h0 : _GEN_85018; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_85020 = 5'h16 == _T_8423[4:0] ? 5'h0 : _GEN_85019; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_85021 = 5'h17 == _T_8423[4:0] ? w_vn_23 : _GEN_85020; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_85022 = 5'h18 == _T_8423[4:0] ? w_vn_24 : _GEN_85021; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_85023 = 5'h19 == _T_8423[4:0] ? 5'h0 : _GEN_85022; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_85024 = 5'h1a == _T_8423[4:0] ? 5'h0 : _GEN_85023; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_85025 = 5'h1b == _T_8423[4:0] ? 5'h0 : _GEN_85024; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_85026 = 5'h1c == _T_8423[4:0] ? 5'h0 : _GEN_85025; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_85027 = 5'h1d == _T_8423[4:0] ? 5'h0 : _GEN_85026; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_85028 = 5'h1e == _T_8423[4:0] ? 5'h0 : _GEN_85027; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_85029 = 5'h1f == _T_8423[4:0] ? 5'h0 : _GEN_85028; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_85033 = 5'h3 == _T_8427[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_85034 = 5'h4 == _T_8427[4:0] ? w_vn_4 : _GEN_85033; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_85035 = 5'h5 == _T_8427[4:0] ? 5'h0 : _GEN_85034; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_85036 = 5'h6 == _T_8427[4:0] ? 5'h0 : _GEN_85035; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_85037 = 5'h7 == _T_8427[4:0] ? w_vn_7 : _GEN_85036; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_85038 = 5'h8 == _T_8427[4:0] ? w_vn_8 : _GEN_85037; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_85039 = 5'h9 == _T_8427[4:0] ? 5'h0 : _GEN_85038; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_85040 = 5'ha == _T_8427[4:0] ? 5'h0 : _GEN_85039; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_85041 = 5'hb == _T_8427[4:0] ? w_vn_11 : _GEN_85040; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_85042 = 5'hc == _T_8427[4:0] ? w_vn_12 : _GEN_85041; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_85043 = 5'hd == _T_8427[4:0] ? w_vn_13 : _GEN_85042; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_85044 = 5'he == _T_8427[4:0] ? 5'h0 : _GEN_85043; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_85045 = 5'hf == _T_8427[4:0] ? w_vn_15 : _GEN_85044; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_85046 = 5'h10 == _T_8427[4:0] ? w_vn_16 : _GEN_85045; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_85047 = 5'h11 == _T_8427[4:0] ? 5'h0 : _GEN_85046; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_85048 = 5'h12 == _T_8427[4:0] ? w_vn_18 : _GEN_85047; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_85049 = 5'h13 == _T_8427[4:0] ? 5'h0 : _GEN_85048; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_85050 = 5'h14 == _T_8427[4:0] ? 5'h0 : _GEN_85049; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_85051 = 5'h15 == _T_8427[4:0] ? 5'h0 : _GEN_85050; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_85052 = 5'h16 == _T_8427[4:0] ? 5'h0 : _GEN_85051; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_85053 = 5'h17 == _T_8427[4:0] ? w_vn_23 : _GEN_85052; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_85054 = 5'h18 == _T_8427[4:0] ? w_vn_24 : _GEN_85053; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_85055 = 5'h19 == _T_8427[4:0] ? 5'h0 : _GEN_85054; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_85056 = 5'h1a == _T_8427[4:0] ? 5'h0 : _GEN_85055; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_85057 = 5'h1b == _T_8427[4:0] ? 5'h0 : _GEN_85056; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_85058 = 5'h1c == _T_8427[4:0] ? 5'h0 : _GEN_85057; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_85059 = 5'h1d == _T_8427[4:0] ? 5'h0 : _GEN_85058; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_85060 = 5'h1e == _T_8427[4:0] ? 5'h0 : _GEN_85059; // @[FanCtrl.scala 490:{41,41}]
  wire [4:0] _GEN_85061 = 5'h1f == _T_8427[4:0] ? 5'h0 : _GEN_85060; // @[FanCtrl.scala 490:{41,41}]
  wire  _T_8429 = _GEN_85029 == _GEN_85061; // @[FanCtrl.scala 490:41]
  wire  _T_8430 = _GEN_84965 == _GEN_84997 & _T_8429; // @[FanCtrl.scala 489:68]
  wire  _T_8449 = _GEN_84997 != _GEN_84840; // @[FanCtrl.scala 492:40]
  wire  _T_8459 = _GEN_85029 != _GEN_84808; // @[FanCtrl.scala 493:41]
  wire  _GEN_85882 = r_valid_1 & _T_8407; // @[FanCtrl.scala 482:33]
  wire [1:0] _GEN_85979 = 4'h0 == _T_8397 ? 2'h0 : _GEN_84757; // @[FanCtrl.scala 520:{46,46}]
  wire [1:0] _GEN_85980 = 4'h1 == _T_8397 ? 2'h0 : _GEN_84758; // @[FanCtrl.scala 520:{46,46}]
  wire [1:0] _GEN_85981 = 4'h2 == _T_8397 ? 2'h0 : _GEN_84759; // @[FanCtrl.scala 520:{46,46}]
  wire [1:0] _GEN_85982 = 4'h3 == _T_8397 ? 2'h0 : _GEN_84760; // @[FanCtrl.scala 520:{46,46}]
  wire [1:0] _GEN_85983 = 4'h4 == _T_8397 ? 2'h0 : _GEN_84761; // @[FanCtrl.scala 520:{46,46}]
  wire [1:0] _GEN_85984 = 4'h5 == _T_8397 ? 2'h0 : _GEN_84762; // @[FanCtrl.scala 520:{46,46}]
  wire [1:0] _GEN_85985 = 4'h6 == _T_8397 ? 2'h0 : _GEN_84763; // @[FanCtrl.scala 520:{46,46}]
  wire [1:0] _GEN_85986 = 4'h7 == _T_8397 ? 2'h0 : _GEN_84764; // @[FanCtrl.scala 520:{46,46}]
  wire [1:0] _GEN_85987 = 4'h8 == _T_8397 ? 2'h0 : _GEN_84765; // @[FanCtrl.scala 520:{46,46}]
  wire [1:0] _GEN_85988 = 4'h9 == _T_8397 ? 2'h0 : _GEN_84766; // @[FanCtrl.scala 520:{46,46}]
  wire [1:0] _GEN_85989 = 4'ha == _T_8397 ? 2'h0 : _GEN_84767; // @[FanCtrl.scala 520:{46,46}]
  wire [1:0] _GEN_85990 = 4'hb == _T_8397 ? 2'h0 : _GEN_84768; // @[FanCtrl.scala 520:{46,46}]
  wire [1:0] _GEN_85991 = 4'hc == _T_8397 ? 2'h0 : _GEN_84769; // @[FanCtrl.scala 520:{46,46}]
  wire [1:0] _GEN_85992 = 4'hd == _T_8397 ? 2'h0 : _GEN_84770; // @[FanCtrl.scala 520:{46,46}]
  wire [1:0] _GEN_85993 = 4'he == _T_8397 ? 2'h0 : _GEN_84771; // @[FanCtrl.scala 520:{46,46}]
  wire [1:0] _GEN_85994 = 4'hf == _T_8397 ? 2'h0 : _GEN_84772; // @[FanCtrl.scala 520:{46,46}]
  wire [1:0] _GEN_85995 = 5'h10 == _GEN_97978 ? 2'h0 : _GEN_84773; // @[FanCtrl.scala 520:{46,46}]
  wire [1:0] _GEN_85996 = 5'h11 == _GEN_97978 ? 2'h0 : _GEN_84774; // @[FanCtrl.scala 520:{46,46}]
  wire [1:0] _GEN_85997 = 5'h12 == _GEN_97978 ? 2'h0 : _GEN_84775; // @[FanCtrl.scala 520:{46,46}]
  wire [1:0] _GEN_85998 = 5'h13 == _GEN_97978 ? 2'h0 : _GEN_84776; // @[FanCtrl.scala 520:{46,46}]
  wire [5:0] _T_8540 = _T_8399 + 6'h5; // @[FanCtrl.scala 522:65]
  wire [4:0] _GEN_86034 = 5'h3 == _T_8540[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 522:{45,45}]
  wire [4:0] _GEN_86035 = 5'h4 == _T_8540[4:0] ? w_vn_4 : _GEN_86034; // @[FanCtrl.scala 522:{45,45}]
  wire [4:0] _GEN_86036 = 5'h5 == _T_8540[4:0] ? 5'h0 : _GEN_86035; // @[FanCtrl.scala 522:{45,45}]
  wire [4:0] _GEN_86037 = 5'h6 == _T_8540[4:0] ? 5'h0 : _GEN_86036; // @[FanCtrl.scala 522:{45,45}]
  wire [4:0] _GEN_86038 = 5'h7 == _T_8540[4:0] ? w_vn_7 : _GEN_86037; // @[FanCtrl.scala 522:{45,45}]
  wire [4:0] _GEN_86039 = 5'h8 == _T_8540[4:0] ? w_vn_8 : _GEN_86038; // @[FanCtrl.scala 522:{45,45}]
  wire [4:0] _GEN_86040 = 5'h9 == _T_8540[4:0] ? 5'h0 : _GEN_86039; // @[FanCtrl.scala 522:{45,45}]
  wire [4:0] _GEN_86041 = 5'ha == _T_8540[4:0] ? 5'h0 : _GEN_86040; // @[FanCtrl.scala 522:{45,45}]
  wire [4:0] _GEN_86042 = 5'hb == _T_8540[4:0] ? w_vn_11 : _GEN_86041; // @[FanCtrl.scala 522:{45,45}]
  wire [4:0] _GEN_86043 = 5'hc == _T_8540[4:0] ? w_vn_12 : _GEN_86042; // @[FanCtrl.scala 522:{45,45}]
  wire [4:0] _GEN_86044 = 5'hd == _T_8540[4:0] ? w_vn_13 : _GEN_86043; // @[FanCtrl.scala 522:{45,45}]
  wire [4:0] _GEN_86045 = 5'he == _T_8540[4:0] ? 5'h0 : _GEN_86044; // @[FanCtrl.scala 522:{45,45}]
  wire [4:0] _GEN_86046 = 5'hf == _T_8540[4:0] ? w_vn_15 : _GEN_86045; // @[FanCtrl.scala 522:{45,45}]
  wire [4:0] _GEN_86047 = 5'h10 == _T_8540[4:0] ? w_vn_16 : _GEN_86046; // @[FanCtrl.scala 522:{45,45}]
  wire [4:0] _GEN_86048 = 5'h11 == _T_8540[4:0] ? 5'h0 : _GEN_86047; // @[FanCtrl.scala 522:{45,45}]
  wire [4:0] _GEN_86049 = 5'h12 == _T_8540[4:0] ? w_vn_18 : _GEN_86048; // @[FanCtrl.scala 522:{45,45}]
  wire [4:0] _GEN_86050 = 5'h13 == _T_8540[4:0] ? 5'h0 : _GEN_86049; // @[FanCtrl.scala 522:{45,45}]
  wire [4:0] _GEN_86051 = 5'h14 == _T_8540[4:0] ? 5'h0 : _GEN_86050; // @[FanCtrl.scala 522:{45,45}]
  wire [4:0] _GEN_86052 = 5'h15 == _T_8540[4:0] ? 5'h0 : _GEN_86051; // @[FanCtrl.scala 522:{45,45}]
  wire [4:0] _GEN_86053 = 5'h16 == _T_8540[4:0] ? 5'h0 : _GEN_86052; // @[FanCtrl.scala 522:{45,45}]
  wire [4:0] _GEN_86054 = 5'h17 == _T_8540[4:0] ? w_vn_23 : _GEN_86053; // @[FanCtrl.scala 522:{45,45}]
  wire [4:0] _GEN_86055 = 5'h18 == _T_8540[4:0] ? w_vn_24 : _GEN_86054; // @[FanCtrl.scala 522:{45,45}]
  wire [4:0] _GEN_86056 = 5'h19 == _T_8540[4:0] ? 5'h0 : _GEN_86055; // @[FanCtrl.scala 522:{45,45}]
  wire [4:0] _GEN_86057 = 5'h1a == _T_8540[4:0] ? 5'h0 : _GEN_86056; // @[FanCtrl.scala 522:{45,45}]
  wire [4:0] _GEN_86058 = 5'h1b == _T_8540[4:0] ? 5'h0 : _GEN_86057; // @[FanCtrl.scala 522:{45,45}]
  wire [4:0] _GEN_86059 = 5'h1c == _T_8540[4:0] ? 5'h0 : _GEN_86058; // @[FanCtrl.scala 522:{45,45}]
  wire [4:0] _GEN_86060 = 5'h1d == _T_8540[4:0] ? 5'h0 : _GEN_86059; // @[FanCtrl.scala 522:{45,45}]
  wire [4:0] _GEN_86061 = 5'h1e == _T_8540[4:0] ? 5'h0 : _GEN_86060; // @[FanCtrl.scala 522:{45,45}]
  wire [4:0] _GEN_86062 = 5'h1f == _T_8540[4:0] ? 5'h0 : _GEN_86061; // @[FanCtrl.scala 522:{45,45}]
  wire [1:0] _GEN_86063 = 4'h0 == _T_8397 ? 2'h1 : _GEN_84757; // @[FanCtrl.scala 524:{45,45}]
  wire [1:0] _GEN_86064 = 4'h1 == _T_8397 ? 2'h1 : _GEN_84758; // @[FanCtrl.scala 524:{45,45}]
  wire [1:0] _GEN_86065 = 4'h2 == _T_8397 ? 2'h1 : _GEN_84759; // @[FanCtrl.scala 524:{45,45}]
  wire [1:0] _GEN_86066 = 4'h3 == _T_8397 ? 2'h1 : _GEN_84760; // @[FanCtrl.scala 524:{45,45}]
  wire [1:0] _GEN_86067 = 4'h4 == _T_8397 ? 2'h1 : _GEN_84761; // @[FanCtrl.scala 524:{45,45}]
  wire [1:0] _GEN_86068 = 4'h5 == _T_8397 ? 2'h1 : _GEN_84762; // @[FanCtrl.scala 524:{45,45}]
  wire [1:0] _GEN_86069 = 4'h6 == _T_8397 ? 2'h1 : _GEN_84763; // @[FanCtrl.scala 524:{45,45}]
  wire [1:0] _GEN_86070 = 4'h7 == _T_8397 ? 2'h1 : _GEN_84764; // @[FanCtrl.scala 524:{45,45}]
  wire [1:0] _GEN_86071 = 4'h8 == _T_8397 ? 2'h1 : _GEN_84765; // @[FanCtrl.scala 524:{45,45}]
  wire [1:0] _GEN_86072 = 4'h9 == _T_8397 ? 2'h1 : _GEN_84766; // @[FanCtrl.scala 524:{45,45}]
  wire [1:0] _GEN_86073 = 4'ha == _T_8397 ? 2'h1 : _GEN_84767; // @[FanCtrl.scala 524:{45,45}]
  wire [1:0] _GEN_86074 = 4'hb == _T_8397 ? 2'h1 : _GEN_84768; // @[FanCtrl.scala 524:{45,45}]
  wire [1:0] _GEN_86075 = 4'hc == _T_8397 ? 2'h1 : _GEN_84769; // @[FanCtrl.scala 524:{45,45}]
  wire [1:0] _GEN_86076 = 4'hd == _T_8397 ? 2'h1 : _GEN_84770; // @[FanCtrl.scala 524:{45,45}]
  wire [1:0] _GEN_86077 = 4'he == _T_8397 ? 2'h1 : _GEN_84771; // @[FanCtrl.scala 524:{45,45}]
  wire [1:0] _GEN_86078 = 4'hf == _T_8397 ? 2'h1 : _GEN_84772; // @[FanCtrl.scala 524:{45,45}]
  wire [1:0] _GEN_86079 = 5'h10 == _GEN_97978 ? 2'h1 : _GEN_84773; // @[FanCtrl.scala 524:{45,45}]
  wire [1:0] _GEN_86080 = 5'h11 == _GEN_97978 ? 2'h1 : _GEN_84774; // @[FanCtrl.scala 524:{45,45}]
  wire [1:0] _GEN_86081 = 5'h12 == _GEN_97978 ? 2'h1 : _GEN_84775; // @[FanCtrl.scala 524:{45,45}]
  wire [1:0] _GEN_86082 = 5'h13 == _GEN_97978 ? 2'h1 : _GEN_84776; // @[FanCtrl.scala 524:{45,45}]
  wire [1:0] _GEN_86083 = 4'h0 == _T_8397 ? 2'h2 : _GEN_84757; // @[FanCtrl.scala 528:{46,46}]
  wire [1:0] _GEN_86084 = 4'h1 == _T_8397 ? 2'h2 : _GEN_84758; // @[FanCtrl.scala 528:{46,46}]
  wire [1:0] _GEN_86085 = 4'h2 == _T_8397 ? 2'h2 : _GEN_84759; // @[FanCtrl.scala 528:{46,46}]
  wire [1:0] _GEN_86086 = 4'h3 == _T_8397 ? 2'h2 : _GEN_84760; // @[FanCtrl.scala 528:{46,46}]
  wire [1:0] _GEN_86087 = 4'h4 == _T_8397 ? 2'h2 : _GEN_84761; // @[FanCtrl.scala 528:{46,46}]
  wire [1:0] _GEN_86088 = 4'h5 == _T_8397 ? 2'h2 : _GEN_84762; // @[FanCtrl.scala 528:{46,46}]
  wire [1:0] _GEN_86089 = 4'h6 == _T_8397 ? 2'h2 : _GEN_84763; // @[FanCtrl.scala 528:{46,46}]
  wire [1:0] _GEN_86090 = 4'h7 == _T_8397 ? 2'h2 : _GEN_84764; // @[FanCtrl.scala 528:{46,46}]
  wire [1:0] _GEN_86091 = 4'h8 == _T_8397 ? 2'h2 : _GEN_84765; // @[FanCtrl.scala 528:{46,46}]
  wire [1:0] _GEN_86092 = 4'h9 == _T_8397 ? 2'h2 : _GEN_84766; // @[FanCtrl.scala 528:{46,46}]
  wire [1:0] _GEN_86093 = 4'ha == _T_8397 ? 2'h2 : _GEN_84767; // @[FanCtrl.scala 528:{46,46}]
  wire [1:0] _GEN_86094 = 4'hb == _T_8397 ? 2'h2 : _GEN_84768; // @[FanCtrl.scala 528:{46,46}]
  wire [1:0] _GEN_86095 = 4'hc == _T_8397 ? 2'h2 : _GEN_84769; // @[FanCtrl.scala 528:{46,46}]
  wire [1:0] _GEN_86096 = 4'hd == _T_8397 ? 2'h2 : _GEN_84770; // @[FanCtrl.scala 528:{46,46}]
  wire [1:0] _GEN_86097 = 4'he == _T_8397 ? 2'h2 : _GEN_84771; // @[FanCtrl.scala 528:{46,46}]
  wire [1:0] _GEN_86098 = 4'hf == _T_8397 ? 2'h2 : _GEN_84772; // @[FanCtrl.scala 528:{46,46}]
  wire [1:0] _GEN_86099 = 5'h10 == _GEN_97978 ? 2'h2 : _GEN_84773; // @[FanCtrl.scala 528:{46,46}]
  wire [1:0] _GEN_86100 = 5'h11 == _GEN_97978 ? 2'h2 : _GEN_84774; // @[FanCtrl.scala 528:{46,46}]
  wire [1:0] _GEN_86101 = 5'h12 == _GEN_97978 ? 2'h2 : _GEN_84775; // @[FanCtrl.scala 528:{46,46}]
  wire [1:0] _GEN_86102 = 5'h13 == _GEN_97978 ? 2'h2 : _GEN_84776; // @[FanCtrl.scala 528:{46,46}]
  wire [1:0] _GEN_86103 = _GEN_84808 == _GEN_86062 ? _GEN_86063 : _GEN_86083; // @[FanCtrl.scala 522:74]
  wire [1:0] _GEN_86104 = _GEN_84808 == _GEN_86062 ? _GEN_86064 : _GEN_86084; // @[FanCtrl.scala 522:74]
  wire [1:0] _GEN_86105 = _GEN_84808 == _GEN_86062 ? _GEN_86065 : _GEN_86085; // @[FanCtrl.scala 522:74]
  wire [1:0] _GEN_86106 = _GEN_84808 == _GEN_86062 ? _GEN_86066 : _GEN_86086; // @[FanCtrl.scala 522:74]
  wire [1:0] _GEN_86107 = _GEN_84808 == _GEN_86062 ? _GEN_86067 : _GEN_86087; // @[FanCtrl.scala 522:74]
  wire [1:0] _GEN_86108 = _GEN_84808 == _GEN_86062 ? _GEN_86068 : _GEN_86088; // @[FanCtrl.scala 522:74]
  wire [1:0] _GEN_86109 = _GEN_84808 == _GEN_86062 ? _GEN_86069 : _GEN_86089; // @[FanCtrl.scala 522:74]
  wire [1:0] _GEN_86110 = _GEN_84808 == _GEN_86062 ? _GEN_86070 : _GEN_86090; // @[FanCtrl.scala 522:74]
  wire [1:0] _GEN_86111 = _GEN_84808 == _GEN_86062 ? _GEN_86071 : _GEN_86091; // @[FanCtrl.scala 522:74]
  wire [1:0] _GEN_86112 = _GEN_84808 == _GEN_86062 ? _GEN_86072 : _GEN_86092; // @[FanCtrl.scala 522:74]
  wire [1:0] _GEN_86113 = _GEN_84808 == _GEN_86062 ? _GEN_86073 : _GEN_86093; // @[FanCtrl.scala 522:74]
  wire [1:0] _GEN_86114 = _GEN_84808 == _GEN_86062 ? _GEN_86074 : _GEN_86094; // @[FanCtrl.scala 522:74]
  wire [1:0] _GEN_86115 = _GEN_84808 == _GEN_86062 ? _GEN_86075 : _GEN_86095; // @[FanCtrl.scala 522:74]
  wire [1:0] _GEN_86116 = _GEN_84808 == _GEN_86062 ? _GEN_86076 : _GEN_86096; // @[FanCtrl.scala 522:74]
  wire [1:0] _GEN_86117 = _GEN_84808 == _GEN_86062 ? _GEN_86077 : _GEN_86097; // @[FanCtrl.scala 522:74]
  wire [1:0] _GEN_86118 = _GEN_84808 == _GEN_86062 ? _GEN_86078 : _GEN_86098; // @[FanCtrl.scala 522:74]
  wire [1:0] _GEN_86119 = _GEN_84808 == _GEN_86062 ? _GEN_86079 : _GEN_86099; // @[FanCtrl.scala 522:74]
  wire [1:0] _GEN_86120 = _GEN_84808 == _GEN_86062 ? _GEN_86080 : _GEN_86100; // @[FanCtrl.scala 522:74]
  wire [1:0] _GEN_86121 = _GEN_84808 == _GEN_86062 ? _GEN_86081 : _GEN_86101; // @[FanCtrl.scala 522:74]
  wire [1:0] _GEN_86122 = _GEN_84808 == _GEN_86062 ? _GEN_86082 : _GEN_86102; // @[FanCtrl.scala 522:74]
  wire [1:0] _GEN_86123 = _GEN_84808 == _GEN_84965 ? _GEN_85979 : _GEN_86103; // @[FanCtrl.scala 518:68]
  wire [1:0] _GEN_86124 = _GEN_84808 == _GEN_84965 ? _GEN_85980 : _GEN_86104; // @[FanCtrl.scala 518:68]
  wire [1:0] _GEN_86125 = _GEN_84808 == _GEN_84965 ? _GEN_85981 : _GEN_86105; // @[FanCtrl.scala 518:68]
  wire [1:0] _GEN_86126 = _GEN_84808 == _GEN_84965 ? _GEN_85982 : _GEN_86106; // @[FanCtrl.scala 518:68]
  wire [1:0] _GEN_86127 = _GEN_84808 == _GEN_84965 ? _GEN_85983 : _GEN_86107; // @[FanCtrl.scala 518:68]
  wire [1:0] _GEN_86128 = _GEN_84808 == _GEN_84965 ? _GEN_85984 : _GEN_86108; // @[FanCtrl.scala 518:68]
  wire [1:0] _GEN_86129 = _GEN_84808 == _GEN_84965 ? _GEN_85985 : _GEN_86109; // @[FanCtrl.scala 518:68]
  wire [1:0] _GEN_86130 = _GEN_84808 == _GEN_84965 ? _GEN_85986 : _GEN_86110; // @[FanCtrl.scala 518:68]
  wire [1:0] _GEN_86131 = _GEN_84808 == _GEN_84965 ? _GEN_85987 : _GEN_86111; // @[FanCtrl.scala 518:68]
  wire [1:0] _GEN_86132 = _GEN_84808 == _GEN_84965 ? _GEN_85988 : _GEN_86112; // @[FanCtrl.scala 518:68]
  wire [1:0] _GEN_86133 = _GEN_84808 == _GEN_84965 ? _GEN_85989 : _GEN_86113; // @[FanCtrl.scala 518:68]
  wire [1:0] _GEN_86134 = _GEN_84808 == _GEN_84965 ? _GEN_85990 : _GEN_86114; // @[FanCtrl.scala 518:68]
  wire [1:0] _GEN_86135 = _GEN_84808 == _GEN_84965 ? _GEN_85991 : _GEN_86115; // @[FanCtrl.scala 518:68]
  wire [1:0] _GEN_86136 = _GEN_84808 == _GEN_84965 ? _GEN_85992 : _GEN_86116; // @[FanCtrl.scala 518:68]
  wire [1:0] _GEN_86137 = _GEN_84808 == _GEN_84965 ? _GEN_85993 : _GEN_86117; // @[FanCtrl.scala 518:68]
  wire [1:0] _GEN_86138 = _GEN_84808 == _GEN_84965 ? _GEN_85994 : _GEN_86118; // @[FanCtrl.scala 518:68]
  wire [1:0] _GEN_86139 = _GEN_84808 == _GEN_84965 ? _GEN_85995 : _GEN_86119; // @[FanCtrl.scala 518:68]
  wire [1:0] _GEN_86140 = _GEN_84808 == _GEN_84965 ? _GEN_85996 : _GEN_86120; // @[FanCtrl.scala 518:68]
  wire [1:0] _GEN_86141 = _GEN_84808 == _GEN_84965 ? _GEN_85997 : _GEN_86121; // @[FanCtrl.scala 518:68]
  wire [1:0] _GEN_86142 = _GEN_84808 == _GEN_84965 ? _GEN_85998 : _GEN_86122; // @[FanCtrl.scala 518:68]
  wire [1:0] _GEN_86163 = r_valid_1 ? _GEN_86123 : _GEN_85979; // @[FanCtrl.scala 517:33]
  wire [1:0] _GEN_86164 = r_valid_1 ? _GEN_86124 : _GEN_85980; // @[FanCtrl.scala 517:33]
  wire [1:0] _GEN_86165 = r_valid_1 ? _GEN_86125 : _GEN_85981; // @[FanCtrl.scala 517:33]
  wire [1:0] _GEN_86166 = r_valid_1 ? _GEN_86126 : _GEN_85982; // @[FanCtrl.scala 517:33]
  wire [1:0] _GEN_86167 = r_valid_1 ? _GEN_86127 : _GEN_85983; // @[FanCtrl.scala 517:33]
  wire [1:0] _GEN_86168 = r_valid_1 ? _GEN_86128 : _GEN_85984; // @[FanCtrl.scala 517:33]
  wire [1:0] _GEN_86169 = r_valid_1 ? _GEN_86129 : _GEN_85985; // @[FanCtrl.scala 517:33]
  wire [1:0] _GEN_86170 = r_valid_1 ? _GEN_86130 : _GEN_85986; // @[FanCtrl.scala 517:33]
  wire [1:0] _GEN_86171 = r_valid_1 ? _GEN_86131 : _GEN_85987; // @[FanCtrl.scala 517:33]
  wire [1:0] _GEN_86172 = r_valid_1 ? _GEN_86132 : _GEN_85988; // @[FanCtrl.scala 517:33]
  wire [1:0] _GEN_86173 = r_valid_1 ? _GEN_86133 : _GEN_85989; // @[FanCtrl.scala 517:33]
  wire [1:0] _GEN_86174 = r_valid_1 ? _GEN_86134 : _GEN_85990; // @[FanCtrl.scala 517:33]
  wire [1:0] _GEN_86175 = r_valid_1 ? _GEN_86135 : _GEN_85991; // @[FanCtrl.scala 517:33]
  wire [1:0] _GEN_86176 = r_valid_1 ? _GEN_86136 : _GEN_85992; // @[FanCtrl.scala 517:33]
  wire [1:0] _GEN_86177 = r_valid_1 ? _GEN_86137 : _GEN_85993; // @[FanCtrl.scala 517:33]
  wire [1:0] _GEN_86178 = r_valid_1 ? _GEN_86138 : _GEN_85994; // @[FanCtrl.scala 517:33]
  wire [1:0] _GEN_86179 = r_valid_1 ? _GEN_86139 : _GEN_85995; // @[FanCtrl.scala 517:33]
  wire [1:0] _GEN_86180 = r_valid_1 ? _GEN_86140 : _GEN_85996; // @[FanCtrl.scala 517:33]
  wire [1:0] _GEN_86181 = r_valid_1 ? _GEN_86141 : _GEN_85997; // @[FanCtrl.scala 517:33]
  wire [1:0] _GEN_86182 = r_valid_1 ? _GEN_86142 : _GEN_85998; // @[FanCtrl.scala 517:33]
  wire [3:0] _T_8564 = _T_8395 + 4'ha; // @[FanCtrl.scala 538:39]
  wire [1:0] _GEN_86247 = 4'h0 == _T_8564 ? 2'h2 : _GEN_86163; // @[FanCtrl.scala 538:{47,47}]
  wire [1:0] _GEN_86248 = 4'h1 == _T_8564 ? 2'h2 : _GEN_86164; // @[FanCtrl.scala 538:{47,47}]
  wire [1:0] _GEN_86249 = 4'h2 == _T_8564 ? 2'h2 : _GEN_86165; // @[FanCtrl.scala 538:{47,47}]
  wire [1:0] _GEN_86250 = 4'h3 == _T_8564 ? 2'h2 : _GEN_86166; // @[FanCtrl.scala 538:{47,47}]
  wire [1:0] _GEN_86251 = 4'h4 == _T_8564 ? 2'h2 : _GEN_86167; // @[FanCtrl.scala 538:{47,47}]
  wire [1:0] _GEN_86252 = 4'h5 == _T_8564 ? 2'h2 : _GEN_86168; // @[FanCtrl.scala 538:{47,47}]
  wire [1:0] _GEN_86253 = 4'h6 == _T_8564 ? 2'h2 : _GEN_86169; // @[FanCtrl.scala 538:{47,47}]
  wire [1:0] _GEN_86254 = 4'h7 == _T_8564 ? 2'h2 : _GEN_86170; // @[FanCtrl.scala 538:{47,47}]
  wire [1:0] _GEN_86255 = 4'h8 == _T_8564 ? 2'h2 : _GEN_86171; // @[FanCtrl.scala 538:{47,47}]
  wire [1:0] _GEN_86256 = 4'h9 == _T_8564 ? 2'h2 : _GEN_86172; // @[FanCtrl.scala 538:{47,47}]
  wire [1:0] _GEN_86257 = 4'ha == _T_8564 ? 2'h2 : _GEN_86173; // @[FanCtrl.scala 538:{47,47}]
  wire [1:0] _GEN_86258 = 4'hb == _T_8564 ? 2'h2 : _GEN_86174; // @[FanCtrl.scala 538:{47,47}]
  wire [1:0] _GEN_86259 = 4'hc == _T_8564 ? 2'h2 : _GEN_86175; // @[FanCtrl.scala 538:{47,47}]
  wire [1:0] _GEN_86260 = 4'hd == _T_8564 ? 2'h2 : _GEN_86176; // @[FanCtrl.scala 538:{47,47}]
  wire [1:0] _GEN_86261 = 4'he == _T_8564 ? 2'h2 : _GEN_86177; // @[FanCtrl.scala 538:{47,47}]
  wire [1:0] _GEN_86262 = 4'hf == _T_8564 ? 2'h2 : _GEN_86178; // @[FanCtrl.scala 538:{47,47}]
  wire [4:0] _GEN_97998 = {{1'd0}, _T_8564}; // @[FanCtrl.scala 538:{47,47}]
  wire [1:0] _GEN_86263 = 5'h10 == _GEN_97998 ? 2'h2 : _GEN_86179; // @[FanCtrl.scala 538:{47,47}]
  wire [1:0] _GEN_86264 = 5'h11 == _GEN_97998 ? 2'h2 : _GEN_86180; // @[FanCtrl.scala 538:{47,47}]
  wire [1:0] _GEN_86265 = 5'h12 == _GEN_97998 ? 2'h2 : _GEN_86181; // @[FanCtrl.scala 538:{47,47}]
  wire [1:0] _GEN_86266 = 5'h13 == _GEN_97998 ? 2'h2 : _GEN_86182; // @[FanCtrl.scala 538:{47,47}]
  wire [5:0] _T_8571 = _T_8399 + 6'ha; // @[FanCtrl.scala 540:65]
  wire [4:0] _GEN_86302 = 5'h3 == _T_8571[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 540:{45,45}]
  wire [4:0] _GEN_86303 = 5'h4 == _T_8571[4:0] ? w_vn_4 : _GEN_86302; // @[FanCtrl.scala 540:{45,45}]
  wire [4:0] _GEN_86304 = 5'h5 == _T_8571[4:0] ? 5'h0 : _GEN_86303; // @[FanCtrl.scala 540:{45,45}]
  wire [4:0] _GEN_86305 = 5'h6 == _T_8571[4:0] ? 5'h0 : _GEN_86304; // @[FanCtrl.scala 540:{45,45}]
  wire [4:0] _GEN_86306 = 5'h7 == _T_8571[4:0] ? w_vn_7 : _GEN_86305; // @[FanCtrl.scala 540:{45,45}]
  wire [4:0] _GEN_86307 = 5'h8 == _T_8571[4:0] ? w_vn_8 : _GEN_86306; // @[FanCtrl.scala 540:{45,45}]
  wire [4:0] _GEN_86308 = 5'h9 == _T_8571[4:0] ? 5'h0 : _GEN_86307; // @[FanCtrl.scala 540:{45,45}]
  wire [4:0] _GEN_86309 = 5'ha == _T_8571[4:0] ? 5'h0 : _GEN_86308; // @[FanCtrl.scala 540:{45,45}]
  wire [4:0] _GEN_86310 = 5'hb == _T_8571[4:0] ? w_vn_11 : _GEN_86309; // @[FanCtrl.scala 540:{45,45}]
  wire [4:0] _GEN_86311 = 5'hc == _T_8571[4:0] ? w_vn_12 : _GEN_86310; // @[FanCtrl.scala 540:{45,45}]
  wire [4:0] _GEN_86312 = 5'hd == _T_8571[4:0] ? w_vn_13 : _GEN_86311; // @[FanCtrl.scala 540:{45,45}]
  wire [4:0] _GEN_86313 = 5'he == _T_8571[4:0] ? 5'h0 : _GEN_86312; // @[FanCtrl.scala 540:{45,45}]
  wire [4:0] _GEN_86314 = 5'hf == _T_8571[4:0] ? w_vn_15 : _GEN_86313; // @[FanCtrl.scala 540:{45,45}]
  wire [4:0] _GEN_86315 = 5'h10 == _T_8571[4:0] ? w_vn_16 : _GEN_86314; // @[FanCtrl.scala 540:{45,45}]
  wire [4:0] _GEN_86316 = 5'h11 == _T_8571[4:0] ? 5'h0 : _GEN_86315; // @[FanCtrl.scala 540:{45,45}]
  wire [4:0] _GEN_86317 = 5'h12 == _T_8571[4:0] ? w_vn_18 : _GEN_86316; // @[FanCtrl.scala 540:{45,45}]
  wire [4:0] _GEN_86318 = 5'h13 == _T_8571[4:0] ? 5'h0 : _GEN_86317; // @[FanCtrl.scala 540:{45,45}]
  wire [4:0] _GEN_86319 = 5'h14 == _T_8571[4:0] ? 5'h0 : _GEN_86318; // @[FanCtrl.scala 540:{45,45}]
  wire [4:0] _GEN_86320 = 5'h15 == _T_8571[4:0] ? 5'h0 : _GEN_86319; // @[FanCtrl.scala 540:{45,45}]
  wire [4:0] _GEN_86321 = 5'h16 == _T_8571[4:0] ? 5'h0 : _GEN_86320; // @[FanCtrl.scala 540:{45,45}]
  wire [4:0] _GEN_86322 = 5'h17 == _T_8571[4:0] ? w_vn_23 : _GEN_86321; // @[FanCtrl.scala 540:{45,45}]
  wire [4:0] _GEN_86323 = 5'h18 == _T_8571[4:0] ? w_vn_24 : _GEN_86322; // @[FanCtrl.scala 540:{45,45}]
  wire [4:0] _GEN_86324 = 5'h19 == _T_8571[4:0] ? 5'h0 : _GEN_86323; // @[FanCtrl.scala 540:{45,45}]
  wire [4:0] _GEN_86325 = 5'h1a == _T_8571[4:0] ? 5'h0 : _GEN_86324; // @[FanCtrl.scala 540:{45,45}]
  wire [4:0] _GEN_86326 = 5'h1b == _T_8571[4:0] ? 5'h0 : _GEN_86325; // @[FanCtrl.scala 540:{45,45}]
  wire [4:0] _GEN_86327 = 5'h1c == _T_8571[4:0] ? 5'h0 : _GEN_86326; // @[FanCtrl.scala 540:{45,45}]
  wire [4:0] _GEN_86328 = 5'h1d == _T_8571[4:0] ? 5'h0 : _GEN_86327; // @[FanCtrl.scala 540:{45,45}]
  wire [4:0] _GEN_86329 = 5'h1e == _T_8571[4:0] ? 5'h0 : _GEN_86328; // @[FanCtrl.scala 540:{45,45}]
  wire [4:0] _GEN_86330 = 5'h1f == _T_8571[4:0] ? 5'h0 : _GEN_86329; // @[FanCtrl.scala 540:{45,45}]
  wire [1:0] _GEN_86331 = 4'h0 == _T_8564 ? 2'h1 : _GEN_86163; // @[FanCtrl.scala 542:{47,47}]
  wire [1:0] _GEN_86332 = 4'h1 == _T_8564 ? 2'h1 : _GEN_86164; // @[FanCtrl.scala 542:{47,47}]
  wire [1:0] _GEN_86333 = 4'h2 == _T_8564 ? 2'h1 : _GEN_86165; // @[FanCtrl.scala 542:{47,47}]
  wire [1:0] _GEN_86334 = 4'h3 == _T_8564 ? 2'h1 : _GEN_86166; // @[FanCtrl.scala 542:{47,47}]
  wire [1:0] _GEN_86335 = 4'h4 == _T_8564 ? 2'h1 : _GEN_86167; // @[FanCtrl.scala 542:{47,47}]
  wire [1:0] _GEN_86336 = 4'h5 == _T_8564 ? 2'h1 : _GEN_86168; // @[FanCtrl.scala 542:{47,47}]
  wire [1:0] _GEN_86337 = 4'h6 == _T_8564 ? 2'h1 : _GEN_86169; // @[FanCtrl.scala 542:{47,47}]
  wire [1:0] _GEN_86338 = 4'h7 == _T_8564 ? 2'h1 : _GEN_86170; // @[FanCtrl.scala 542:{47,47}]
  wire [1:0] _GEN_86339 = 4'h8 == _T_8564 ? 2'h1 : _GEN_86171; // @[FanCtrl.scala 542:{47,47}]
  wire [1:0] _GEN_86340 = 4'h9 == _T_8564 ? 2'h1 : _GEN_86172; // @[FanCtrl.scala 542:{47,47}]
  wire [1:0] _GEN_86341 = 4'ha == _T_8564 ? 2'h1 : _GEN_86173; // @[FanCtrl.scala 542:{47,47}]
  wire [1:0] _GEN_86342 = 4'hb == _T_8564 ? 2'h1 : _GEN_86174; // @[FanCtrl.scala 542:{47,47}]
  wire [1:0] _GEN_86343 = 4'hc == _T_8564 ? 2'h1 : _GEN_86175; // @[FanCtrl.scala 542:{47,47}]
  wire [1:0] _GEN_86344 = 4'hd == _T_8564 ? 2'h1 : _GEN_86176; // @[FanCtrl.scala 542:{47,47}]
  wire [1:0] _GEN_86345 = 4'he == _T_8564 ? 2'h1 : _GEN_86177; // @[FanCtrl.scala 542:{47,47}]
  wire [1:0] _GEN_86346 = 4'hf == _T_8564 ? 2'h1 : _GEN_86178; // @[FanCtrl.scala 542:{47,47}]
  wire [1:0] _GEN_86347 = 5'h10 == _GEN_97998 ? 2'h1 : _GEN_86179; // @[FanCtrl.scala 542:{47,47}]
  wire [1:0] _GEN_86348 = 5'h11 == _GEN_97998 ? 2'h1 : _GEN_86180; // @[FanCtrl.scala 542:{47,47}]
  wire [1:0] _GEN_86349 = 5'h12 == _GEN_97998 ? 2'h1 : _GEN_86181; // @[FanCtrl.scala 542:{47,47}]
  wire [1:0] _GEN_86350 = 5'h13 == _GEN_97998 ? 2'h1 : _GEN_86182; // @[FanCtrl.scala 542:{47,47}]
  wire [1:0] _GEN_86351 = 4'h0 == _T_8564 ? 2'h0 : _GEN_86163; // @[FanCtrl.scala 545:{47,47}]
  wire [1:0] _GEN_86352 = 4'h1 == _T_8564 ? 2'h0 : _GEN_86164; // @[FanCtrl.scala 545:{47,47}]
  wire [1:0] _GEN_86353 = 4'h2 == _T_8564 ? 2'h0 : _GEN_86165; // @[FanCtrl.scala 545:{47,47}]
  wire [1:0] _GEN_86354 = 4'h3 == _T_8564 ? 2'h0 : _GEN_86166; // @[FanCtrl.scala 545:{47,47}]
  wire [1:0] _GEN_86355 = 4'h4 == _T_8564 ? 2'h0 : _GEN_86167; // @[FanCtrl.scala 545:{47,47}]
  wire [1:0] _GEN_86356 = 4'h5 == _T_8564 ? 2'h0 : _GEN_86168; // @[FanCtrl.scala 545:{47,47}]
  wire [1:0] _GEN_86357 = 4'h6 == _T_8564 ? 2'h0 : _GEN_86169; // @[FanCtrl.scala 545:{47,47}]
  wire [1:0] _GEN_86358 = 4'h7 == _T_8564 ? 2'h0 : _GEN_86170; // @[FanCtrl.scala 545:{47,47}]
  wire [1:0] _GEN_86359 = 4'h8 == _T_8564 ? 2'h0 : _GEN_86171; // @[FanCtrl.scala 545:{47,47}]
  wire [1:0] _GEN_86360 = 4'h9 == _T_8564 ? 2'h0 : _GEN_86172; // @[FanCtrl.scala 545:{47,47}]
  wire [1:0] _GEN_86361 = 4'ha == _T_8564 ? 2'h0 : _GEN_86173; // @[FanCtrl.scala 545:{47,47}]
  wire [1:0] _GEN_86362 = 4'hb == _T_8564 ? 2'h0 : _GEN_86174; // @[FanCtrl.scala 545:{47,47}]
  wire [1:0] _GEN_86363 = 4'hc == _T_8564 ? 2'h0 : _GEN_86175; // @[FanCtrl.scala 545:{47,47}]
  wire [1:0] _GEN_86364 = 4'hd == _T_8564 ? 2'h0 : _GEN_86176; // @[FanCtrl.scala 545:{47,47}]
  wire [1:0] _GEN_86365 = 4'he == _T_8564 ? 2'h0 : _GEN_86177; // @[FanCtrl.scala 545:{47,47}]
  wire [1:0] _GEN_86366 = 4'hf == _T_8564 ? 2'h0 : _GEN_86178; // @[FanCtrl.scala 545:{47,47}]
  wire [1:0] _GEN_86367 = 5'h10 == _GEN_97998 ? 2'h0 : _GEN_86179; // @[FanCtrl.scala 545:{47,47}]
  wire [1:0] _GEN_86368 = 5'h11 == _GEN_97998 ? 2'h0 : _GEN_86180; // @[FanCtrl.scala 545:{47,47}]
  wire [1:0] _GEN_86369 = 5'h12 == _GEN_97998 ? 2'h0 : _GEN_86181; // @[FanCtrl.scala 545:{47,47}]
  wire [1:0] _GEN_86370 = 5'h13 == _GEN_97998 ? 2'h0 : _GEN_86182; // @[FanCtrl.scala 545:{47,47}]
  wire [1:0] _GEN_86371 = _GEN_84840 == _GEN_86330 ? _GEN_86331 : _GEN_86351; // @[FanCtrl.scala 540:74]
  wire [1:0] _GEN_86372 = _GEN_84840 == _GEN_86330 ? _GEN_86332 : _GEN_86352; // @[FanCtrl.scala 540:74]
  wire [1:0] _GEN_86373 = _GEN_84840 == _GEN_86330 ? _GEN_86333 : _GEN_86353; // @[FanCtrl.scala 540:74]
  wire [1:0] _GEN_86374 = _GEN_84840 == _GEN_86330 ? _GEN_86334 : _GEN_86354; // @[FanCtrl.scala 540:74]
  wire [1:0] _GEN_86375 = _GEN_84840 == _GEN_86330 ? _GEN_86335 : _GEN_86355; // @[FanCtrl.scala 540:74]
  wire [1:0] _GEN_86376 = _GEN_84840 == _GEN_86330 ? _GEN_86336 : _GEN_86356; // @[FanCtrl.scala 540:74]
  wire [1:0] _GEN_86377 = _GEN_84840 == _GEN_86330 ? _GEN_86337 : _GEN_86357; // @[FanCtrl.scala 540:74]
  wire [1:0] _GEN_86378 = _GEN_84840 == _GEN_86330 ? _GEN_86338 : _GEN_86358; // @[FanCtrl.scala 540:74]
  wire [1:0] _GEN_86379 = _GEN_84840 == _GEN_86330 ? _GEN_86339 : _GEN_86359; // @[FanCtrl.scala 540:74]
  wire [1:0] _GEN_86380 = _GEN_84840 == _GEN_86330 ? _GEN_86340 : _GEN_86360; // @[FanCtrl.scala 540:74]
  wire [1:0] _GEN_86381 = _GEN_84840 == _GEN_86330 ? _GEN_86341 : _GEN_86361; // @[FanCtrl.scala 540:74]
  wire [1:0] _GEN_86382 = _GEN_84840 == _GEN_86330 ? _GEN_86342 : _GEN_86362; // @[FanCtrl.scala 540:74]
  wire [1:0] _GEN_86383 = _GEN_84840 == _GEN_86330 ? _GEN_86343 : _GEN_86363; // @[FanCtrl.scala 540:74]
  wire [1:0] _GEN_86384 = _GEN_84840 == _GEN_86330 ? _GEN_86344 : _GEN_86364; // @[FanCtrl.scala 540:74]
  wire [1:0] _GEN_86385 = _GEN_84840 == _GEN_86330 ? _GEN_86345 : _GEN_86365; // @[FanCtrl.scala 540:74]
  wire [1:0] _GEN_86386 = _GEN_84840 == _GEN_86330 ? _GEN_86346 : _GEN_86366; // @[FanCtrl.scala 540:74]
  wire [1:0] _GEN_86387 = _GEN_84840 == _GEN_86330 ? _GEN_86347 : _GEN_86367; // @[FanCtrl.scala 540:74]
  wire [1:0] _GEN_86388 = _GEN_84840 == _GEN_86330 ? _GEN_86348 : _GEN_86368; // @[FanCtrl.scala 540:74]
  wire [1:0] _GEN_86389 = _GEN_84840 == _GEN_86330 ? _GEN_86349 : _GEN_86369; // @[FanCtrl.scala 540:74]
  wire [1:0] _GEN_86390 = _GEN_84840 == _GEN_86330 ? _GEN_86350 : _GEN_86370; // @[FanCtrl.scala 540:74]
  wire [1:0] _GEN_86391 = _GEN_84840 == _GEN_85061 ? _GEN_86247 : _GEN_86371; // @[FanCtrl.scala 536:69]
  wire [1:0] _GEN_86392 = _GEN_84840 == _GEN_85061 ? _GEN_86248 : _GEN_86372; // @[FanCtrl.scala 536:69]
  wire [1:0] _GEN_86393 = _GEN_84840 == _GEN_85061 ? _GEN_86249 : _GEN_86373; // @[FanCtrl.scala 536:69]
  wire [1:0] _GEN_86394 = _GEN_84840 == _GEN_85061 ? _GEN_86250 : _GEN_86374; // @[FanCtrl.scala 536:69]
  wire [1:0] _GEN_86395 = _GEN_84840 == _GEN_85061 ? _GEN_86251 : _GEN_86375; // @[FanCtrl.scala 536:69]
  wire [1:0] _GEN_86396 = _GEN_84840 == _GEN_85061 ? _GEN_86252 : _GEN_86376; // @[FanCtrl.scala 536:69]
  wire [1:0] _GEN_86397 = _GEN_84840 == _GEN_85061 ? _GEN_86253 : _GEN_86377; // @[FanCtrl.scala 536:69]
  wire [1:0] _GEN_86398 = _GEN_84840 == _GEN_85061 ? _GEN_86254 : _GEN_86378; // @[FanCtrl.scala 536:69]
  wire [1:0] _GEN_86399 = _GEN_84840 == _GEN_85061 ? _GEN_86255 : _GEN_86379; // @[FanCtrl.scala 536:69]
  wire [1:0] _GEN_86400 = _GEN_84840 == _GEN_85061 ? _GEN_86256 : _GEN_86380; // @[FanCtrl.scala 536:69]
  wire [1:0] _GEN_86401 = _GEN_84840 == _GEN_85061 ? _GEN_86257 : _GEN_86381; // @[FanCtrl.scala 536:69]
  wire [1:0] _GEN_86402 = _GEN_84840 == _GEN_85061 ? _GEN_86258 : _GEN_86382; // @[FanCtrl.scala 536:69]
  wire [1:0] _GEN_86403 = _GEN_84840 == _GEN_85061 ? _GEN_86259 : _GEN_86383; // @[FanCtrl.scala 536:69]
  wire [1:0] _GEN_86404 = _GEN_84840 == _GEN_85061 ? _GEN_86260 : _GEN_86384; // @[FanCtrl.scala 536:69]
  wire [1:0] _GEN_86405 = _GEN_84840 == _GEN_85061 ? _GEN_86261 : _GEN_86385; // @[FanCtrl.scala 536:69]
  wire [1:0] _GEN_86406 = _GEN_84840 == _GEN_85061 ? _GEN_86262 : _GEN_86386; // @[FanCtrl.scala 536:69]
  wire [1:0] _GEN_86407 = _GEN_84840 == _GEN_85061 ? _GEN_86263 : _GEN_86387; // @[FanCtrl.scala 536:69]
  wire [1:0] _GEN_86408 = _GEN_84840 == _GEN_85061 ? _GEN_86264 : _GEN_86388; // @[FanCtrl.scala 536:69]
  wire [1:0] _GEN_86409 = _GEN_84840 == _GEN_85061 ? _GEN_86265 : _GEN_86389; // @[FanCtrl.scala 536:69]
  wire [1:0] _GEN_86410 = _GEN_84840 == _GEN_85061 ? _GEN_86266 : _GEN_86390; // @[FanCtrl.scala 536:69]
  wire [1:0] _GEN_86411 = 4'h0 == _T_8397 ? 2'h0 : _GEN_86163; // @[FanCtrl.scala 548:{44,44}]
  wire [1:0] _GEN_86412 = 4'h1 == _T_8397 ? 2'h0 : _GEN_86164; // @[FanCtrl.scala 548:{44,44}]
  wire [1:0] _GEN_86413 = 4'h2 == _T_8397 ? 2'h0 : _GEN_86165; // @[FanCtrl.scala 548:{44,44}]
  wire [1:0] _GEN_86414 = 4'h3 == _T_8397 ? 2'h0 : _GEN_86166; // @[FanCtrl.scala 548:{44,44}]
  wire [1:0] _GEN_86415 = 4'h4 == _T_8397 ? 2'h0 : _GEN_86167; // @[FanCtrl.scala 548:{44,44}]
  wire [1:0] _GEN_86416 = 4'h5 == _T_8397 ? 2'h0 : _GEN_86168; // @[FanCtrl.scala 548:{44,44}]
  wire [1:0] _GEN_86417 = 4'h6 == _T_8397 ? 2'h0 : _GEN_86169; // @[FanCtrl.scala 548:{44,44}]
  wire [1:0] _GEN_86418 = 4'h7 == _T_8397 ? 2'h0 : _GEN_86170; // @[FanCtrl.scala 548:{44,44}]
  wire [1:0] _GEN_86419 = 4'h8 == _T_8397 ? 2'h0 : _GEN_86171; // @[FanCtrl.scala 548:{44,44}]
  wire [1:0] _GEN_86420 = 4'h9 == _T_8397 ? 2'h0 : _GEN_86172; // @[FanCtrl.scala 548:{44,44}]
  wire [1:0] _GEN_86421 = 4'ha == _T_8397 ? 2'h0 : _GEN_86173; // @[FanCtrl.scala 548:{44,44}]
  wire [1:0] _GEN_86422 = 4'hb == _T_8397 ? 2'h0 : _GEN_86174; // @[FanCtrl.scala 548:{44,44}]
  wire [1:0] _GEN_86423 = 4'hc == _T_8397 ? 2'h0 : _GEN_86175; // @[FanCtrl.scala 548:{44,44}]
  wire [1:0] _GEN_86424 = 4'hd == _T_8397 ? 2'h0 : _GEN_86176; // @[FanCtrl.scala 548:{44,44}]
  wire [1:0] _GEN_86425 = 4'he == _T_8397 ? 2'h0 : _GEN_86177; // @[FanCtrl.scala 548:{44,44}]
  wire [1:0] _GEN_86426 = 4'hf == _T_8397 ? 2'h0 : _GEN_86178; // @[FanCtrl.scala 548:{44,44}]
  wire [1:0] _GEN_86427 = 5'h10 == _GEN_97978 ? 2'h0 : _GEN_86179; // @[FanCtrl.scala 548:{44,44}]
  wire [1:0] _GEN_86428 = 5'h11 == _GEN_97978 ? 2'h0 : _GEN_86180; // @[FanCtrl.scala 548:{44,44}]
  wire [1:0] _GEN_86429 = 5'h12 == _GEN_97978 ? 2'h0 : _GEN_86181; // @[FanCtrl.scala 548:{44,44}]
  wire [1:0] _GEN_86430 = 5'h13 == _GEN_97978 ? 2'h0 : _GEN_86182; // @[FanCtrl.scala 548:{44,44}]
  wire [1:0] _GEN_86431 = r_valid_1 ? _GEN_86391 : _GEN_86411; // @[FanCtrl.scala 535:33]
  wire [1:0] _GEN_86432 = r_valid_1 ? _GEN_86392 : _GEN_86412; // @[FanCtrl.scala 535:33]
  wire [1:0] _GEN_86433 = r_valid_1 ? _GEN_86393 : _GEN_86413; // @[FanCtrl.scala 535:33]
  wire [1:0] _GEN_86434 = r_valid_1 ? _GEN_86394 : _GEN_86414; // @[FanCtrl.scala 535:33]
  wire [1:0] _GEN_86435 = r_valid_1 ? _GEN_86395 : _GEN_86415; // @[FanCtrl.scala 535:33]
  wire [1:0] _GEN_86436 = r_valid_1 ? _GEN_86396 : _GEN_86416; // @[FanCtrl.scala 535:33]
  wire [1:0] _GEN_86437 = r_valid_1 ? _GEN_86397 : _GEN_86417; // @[FanCtrl.scala 535:33]
  wire [1:0] _GEN_86438 = r_valid_1 ? _GEN_86398 : _GEN_86418; // @[FanCtrl.scala 535:33]
  wire [1:0] _GEN_86439 = r_valid_1 ? _GEN_86399 : _GEN_86419; // @[FanCtrl.scala 535:33]
  wire [1:0] _GEN_86440 = r_valid_1 ? _GEN_86400 : _GEN_86420; // @[FanCtrl.scala 535:33]
  wire [1:0] _GEN_86441 = r_valid_1 ? _GEN_86401 : _GEN_86421; // @[FanCtrl.scala 535:33]
  wire [1:0] _GEN_86442 = r_valid_1 ? _GEN_86402 : _GEN_86422; // @[FanCtrl.scala 535:33]
  wire [1:0] _GEN_86443 = r_valid_1 ? _GEN_86403 : _GEN_86423; // @[FanCtrl.scala 535:33]
  wire [1:0] _GEN_86444 = r_valid_1 ? _GEN_86404 : _GEN_86424; // @[FanCtrl.scala 535:33]
  wire [1:0] _GEN_86445 = r_valid_1 ? _GEN_86405 : _GEN_86425; // @[FanCtrl.scala 535:33]
  wire [1:0] _GEN_86446 = r_valid_1 ? _GEN_86406 : _GEN_86426; // @[FanCtrl.scala 535:33]
  wire [1:0] _GEN_86447 = r_valid_1 ? _GEN_86407 : _GEN_86427; // @[FanCtrl.scala 535:33]
  wire [1:0] _GEN_86448 = r_valid_1 ? _GEN_86408 : _GEN_86428; // @[FanCtrl.scala 535:33]
  wire [1:0] _GEN_86449 = r_valid_1 ? _GEN_86409 : _GEN_86429; // @[FanCtrl.scala 535:33]
  wire [1:0] _GEN_86450 = r_valid_1 ? _GEN_86410 : _GEN_86430; // @[FanCtrl.scala 535:33]
  wire [5:0] _T_8630 = _T_8399 - 6'h1; // @[FanCtrl.scala 567:61]
  wire [4:0] _GEN_86853 = 5'h3 == _T_8630[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 567:{41,41}]
  wire [4:0] _GEN_86854 = 5'h4 == _T_8630[4:0] ? w_vn_4 : _GEN_86853; // @[FanCtrl.scala 567:{41,41}]
  wire [4:0] _GEN_86855 = 5'h5 == _T_8630[4:0] ? 5'h0 : _GEN_86854; // @[FanCtrl.scala 567:{41,41}]
  wire [4:0] _GEN_86856 = 5'h6 == _T_8630[4:0] ? 5'h0 : _GEN_86855; // @[FanCtrl.scala 567:{41,41}]
  wire [4:0] _GEN_86857 = 5'h7 == _T_8630[4:0] ? w_vn_7 : _GEN_86856; // @[FanCtrl.scala 567:{41,41}]
  wire [4:0] _GEN_86858 = 5'h8 == _T_8630[4:0] ? w_vn_8 : _GEN_86857; // @[FanCtrl.scala 567:{41,41}]
  wire [4:0] _GEN_86859 = 5'h9 == _T_8630[4:0] ? 5'h0 : _GEN_86858; // @[FanCtrl.scala 567:{41,41}]
  wire [4:0] _GEN_86860 = 5'ha == _T_8630[4:0] ? 5'h0 : _GEN_86859; // @[FanCtrl.scala 567:{41,41}]
  wire [4:0] _GEN_86861 = 5'hb == _T_8630[4:0] ? w_vn_11 : _GEN_86860; // @[FanCtrl.scala 567:{41,41}]
  wire [4:0] _GEN_86862 = 5'hc == _T_8630[4:0] ? w_vn_12 : _GEN_86861; // @[FanCtrl.scala 567:{41,41}]
  wire [4:0] _GEN_86863 = 5'hd == _T_8630[4:0] ? w_vn_13 : _GEN_86862; // @[FanCtrl.scala 567:{41,41}]
  wire [4:0] _GEN_86864 = 5'he == _T_8630[4:0] ? 5'h0 : _GEN_86863; // @[FanCtrl.scala 567:{41,41}]
  wire [4:0] _GEN_86865 = 5'hf == _T_8630[4:0] ? w_vn_15 : _GEN_86864; // @[FanCtrl.scala 567:{41,41}]
  wire [4:0] _GEN_86866 = 5'h10 == _T_8630[4:0] ? w_vn_16 : _GEN_86865; // @[FanCtrl.scala 567:{41,41}]
  wire [4:0] _GEN_86867 = 5'h11 == _T_8630[4:0] ? 5'h0 : _GEN_86866; // @[FanCtrl.scala 567:{41,41}]
  wire [4:0] _GEN_86868 = 5'h12 == _T_8630[4:0] ? w_vn_18 : _GEN_86867; // @[FanCtrl.scala 567:{41,41}]
  wire [4:0] _GEN_86869 = 5'h13 == _T_8630[4:0] ? 5'h0 : _GEN_86868; // @[FanCtrl.scala 567:{41,41}]
  wire [4:0] _GEN_86870 = 5'h14 == _T_8630[4:0] ? 5'h0 : _GEN_86869; // @[FanCtrl.scala 567:{41,41}]
  wire [4:0] _GEN_86871 = 5'h15 == _T_8630[4:0] ? 5'h0 : _GEN_86870; // @[FanCtrl.scala 567:{41,41}]
  wire [4:0] _GEN_86872 = 5'h16 == _T_8630[4:0] ? 5'h0 : _GEN_86871; // @[FanCtrl.scala 567:{41,41}]
  wire [4:0] _GEN_86873 = 5'h17 == _T_8630[4:0] ? w_vn_23 : _GEN_86872; // @[FanCtrl.scala 567:{41,41}]
  wire [4:0] _GEN_86874 = 5'h18 == _T_8630[4:0] ? w_vn_24 : _GEN_86873; // @[FanCtrl.scala 567:{41,41}]
  wire [4:0] _GEN_86875 = 5'h19 == _T_8630[4:0] ? 5'h0 : _GEN_86874; // @[FanCtrl.scala 567:{41,41}]
  wire [4:0] _GEN_86876 = 5'h1a == _T_8630[4:0] ? 5'h0 : _GEN_86875; // @[FanCtrl.scala 567:{41,41}]
  wire [4:0] _GEN_86877 = 5'h1b == _T_8630[4:0] ? 5'h0 : _GEN_86876; // @[FanCtrl.scala 567:{41,41}]
  wire [4:0] _GEN_86878 = 5'h1c == _T_8630[4:0] ? 5'h0 : _GEN_86877; // @[FanCtrl.scala 567:{41,41}]
  wire [4:0] _GEN_86879 = 5'h1d == _T_8630[4:0] ? 5'h0 : _GEN_86878; // @[FanCtrl.scala 567:{41,41}]
  wire [4:0] _GEN_86880 = 5'h1e == _T_8630[4:0] ? 5'h0 : _GEN_86879; // @[FanCtrl.scala 567:{41,41}]
  wire [4:0] _GEN_86881 = 5'h1f == _T_8630[4:0] ? 5'h0 : _GEN_86880; // @[FanCtrl.scala 567:{41,41}]
  wire  _T_8632 = _GEN_84965 != _GEN_86881; // @[FanCtrl.scala 567:41]
  wire  _T_8633 = _T_8430 & _T_8632; // @[FanCtrl.scala 566:73]
  wire  _T_8643 = _T_8633 & _T_8449; // @[FanCtrl.scala 567:69]
  wire  _T_8653 = _T_8643 & _T_8459; // @[FanCtrl.scala 568:71]
  wire  _T_8674 = _T_8420 & _T_8632; // @[FanCtrl.scala 573:77]
  wire  _T_8683 = _GEN_84840 != _GEN_84997; // @[FanCtrl.scala 575:47]
  wire  _T_8684 = _T_8674 & _T_8683; // @[FanCtrl.scala 574:76]
  wire  _T_8705 = _T_8429 & _T_8459; // @[FanCtrl.scala 579:79]
  wire [2:0] _GEN_87483 = _T_8705 ? 3'h4 : 3'h0; // @[FanCtrl.scala 580:78]
  wire [4:0] _GEN_98086 = {{1'd0}, _T_7797}; // @[FanCtrl.scala 697:35]
  wire [4:0] _T_8995 = _GEN_98086 + 5'h10; // @[FanCtrl.scala 697:35]
  wire [1:0] _GEN_90317 = 5'h0 == _T_8995 ? 2'h0 : _GEN_86431; // @[FanCtrl.scala 697:{43,43}]
  wire [1:0] _GEN_90318 = 5'h1 == _T_8995 ? 2'h0 : _GEN_86432; // @[FanCtrl.scala 697:{43,43}]
  wire [1:0] _GEN_90319 = 5'h2 == _T_8995 ? 2'h0 : _GEN_86433; // @[FanCtrl.scala 697:{43,43}]
  wire [1:0] _GEN_90320 = 5'h3 == _T_8995 ? 2'h0 : _GEN_86434; // @[FanCtrl.scala 697:{43,43}]
  wire [1:0] _GEN_90321 = 5'h4 == _T_8995 ? 2'h0 : _GEN_86435; // @[FanCtrl.scala 697:{43,43}]
  wire [1:0] _GEN_90322 = 5'h5 == _T_8995 ? 2'h0 : _GEN_86436; // @[FanCtrl.scala 697:{43,43}]
  wire [1:0] _GEN_90323 = 5'h6 == _T_8995 ? 2'h0 : _GEN_86437; // @[FanCtrl.scala 697:{43,43}]
  wire [1:0] _GEN_90324 = 5'h7 == _T_8995 ? 2'h0 : _GEN_86438; // @[FanCtrl.scala 697:{43,43}]
  wire [1:0] _GEN_90325 = 5'h8 == _T_8995 ? 2'h0 : _GEN_86439; // @[FanCtrl.scala 697:{43,43}]
  wire [1:0] _GEN_90326 = 5'h9 == _T_8995 ? 2'h0 : _GEN_86440; // @[FanCtrl.scala 697:{43,43}]
  wire [1:0] _GEN_90327 = 5'ha == _T_8995 ? 2'h0 : _GEN_86441; // @[FanCtrl.scala 697:{43,43}]
  wire [1:0] _GEN_90328 = 5'hb == _T_8995 ? 2'h0 : _GEN_86442; // @[FanCtrl.scala 697:{43,43}]
  wire [1:0] _GEN_90329 = 5'hc == _T_8995 ? 2'h0 : _GEN_86443; // @[FanCtrl.scala 697:{43,43}]
  wire [1:0] _GEN_90330 = 5'hd == _T_8995 ? 2'h0 : _GEN_86444; // @[FanCtrl.scala 697:{43,43}]
  wire [1:0] _GEN_90331 = 5'he == _T_8995 ? 2'h0 : _GEN_86445; // @[FanCtrl.scala 697:{43,43}]
  wire [1:0] _GEN_90332 = 5'hf == _T_8995 ? 2'h0 : _GEN_86446; // @[FanCtrl.scala 697:{43,43}]
  wire [1:0] _GEN_90333 = 5'h10 == _T_8995 ? 2'h0 : _GEN_86447; // @[FanCtrl.scala 697:{43,43}]
  wire [1:0] _GEN_90334 = 5'h11 == _T_8995 ? 2'h0 : _GEN_86448; // @[FanCtrl.scala 697:{43,43}]
  wire [1:0] _GEN_90335 = 5'h12 == _T_8995 ? 2'h0 : _GEN_86449; // @[FanCtrl.scala 697:{43,43}]
  wire [1:0] _GEN_90336 = 5'h13 == _T_8995 ? 2'h0 : _GEN_86450; // @[FanCtrl.scala 697:{43,43}]
  wire [6:0] _T_8997 = 6'h20 * 1'h0; // @[FanCtrl.scala 700:25]
  wire [6:0] _T_8999 = _T_8997 + 7'hf; // @[FanCtrl.scala 700:31]
  wire [6:0] _T_9003 = _T_8997 + 7'h10; // @[FanCtrl.scala 700:60]
  wire [4:0] _GEN_90340 = 5'h3 == _T_8999[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 700:{40,40}]
  wire [4:0] _GEN_90341 = 5'h4 == _T_8999[4:0] ? w_vn_4 : _GEN_90340; // @[FanCtrl.scala 700:{40,40}]
  wire [4:0] _GEN_90342 = 5'h5 == _T_8999[4:0] ? 5'h0 : _GEN_90341; // @[FanCtrl.scala 700:{40,40}]
  wire [4:0] _GEN_90343 = 5'h6 == _T_8999[4:0] ? 5'h0 : _GEN_90342; // @[FanCtrl.scala 700:{40,40}]
  wire [4:0] _GEN_90344 = 5'h7 == _T_8999[4:0] ? w_vn_7 : _GEN_90343; // @[FanCtrl.scala 700:{40,40}]
  wire [4:0] _GEN_90345 = 5'h8 == _T_8999[4:0] ? w_vn_8 : _GEN_90344; // @[FanCtrl.scala 700:{40,40}]
  wire [4:0] _GEN_90346 = 5'h9 == _T_8999[4:0] ? 5'h0 : _GEN_90345; // @[FanCtrl.scala 700:{40,40}]
  wire [4:0] _GEN_90347 = 5'ha == _T_8999[4:0] ? 5'h0 : _GEN_90346; // @[FanCtrl.scala 700:{40,40}]
  wire [4:0] _GEN_90348 = 5'hb == _T_8999[4:0] ? w_vn_11 : _GEN_90347; // @[FanCtrl.scala 700:{40,40}]
  wire [4:0] _GEN_90349 = 5'hc == _T_8999[4:0] ? w_vn_12 : _GEN_90348; // @[FanCtrl.scala 700:{40,40}]
  wire [4:0] _GEN_90350 = 5'hd == _T_8999[4:0] ? w_vn_13 : _GEN_90349; // @[FanCtrl.scala 700:{40,40}]
  wire [4:0] _GEN_90351 = 5'he == _T_8999[4:0] ? 5'h0 : _GEN_90350; // @[FanCtrl.scala 700:{40,40}]
  wire [4:0] _GEN_90352 = 5'hf == _T_8999[4:0] ? w_vn_15 : _GEN_90351; // @[FanCtrl.scala 700:{40,40}]
  wire [4:0] _GEN_90353 = 5'h10 == _T_8999[4:0] ? w_vn_16 : _GEN_90352; // @[FanCtrl.scala 700:{40,40}]
  wire [4:0] _GEN_90354 = 5'h11 == _T_8999[4:0] ? 5'h0 : _GEN_90353; // @[FanCtrl.scala 700:{40,40}]
  wire [4:0] _GEN_90355 = 5'h12 == _T_8999[4:0] ? w_vn_18 : _GEN_90354; // @[FanCtrl.scala 700:{40,40}]
  wire [4:0] _GEN_90356 = 5'h13 == _T_8999[4:0] ? 5'h0 : _GEN_90355; // @[FanCtrl.scala 700:{40,40}]
  wire [4:0] _GEN_90357 = 5'h14 == _T_8999[4:0] ? 5'h0 : _GEN_90356; // @[FanCtrl.scala 700:{40,40}]
  wire [4:0] _GEN_90358 = 5'h15 == _T_8999[4:0] ? 5'h0 : _GEN_90357; // @[FanCtrl.scala 700:{40,40}]
  wire [4:0] _GEN_90359 = 5'h16 == _T_8999[4:0] ? 5'h0 : _GEN_90358; // @[FanCtrl.scala 700:{40,40}]
  wire [4:0] _GEN_90360 = 5'h17 == _T_8999[4:0] ? w_vn_23 : _GEN_90359; // @[FanCtrl.scala 700:{40,40}]
  wire [4:0] _GEN_90361 = 5'h18 == _T_8999[4:0] ? w_vn_24 : _GEN_90360; // @[FanCtrl.scala 700:{40,40}]
  wire [4:0] _GEN_90362 = 5'h19 == _T_8999[4:0] ? 5'h0 : _GEN_90361; // @[FanCtrl.scala 700:{40,40}]
  wire [4:0] _GEN_90363 = 5'h1a == _T_8999[4:0] ? 5'h0 : _GEN_90362; // @[FanCtrl.scala 700:{40,40}]
  wire [4:0] _GEN_90364 = 5'h1b == _T_8999[4:0] ? 5'h0 : _GEN_90363; // @[FanCtrl.scala 700:{40,40}]
  wire [4:0] _GEN_90365 = 5'h1c == _T_8999[4:0] ? 5'h0 : _GEN_90364; // @[FanCtrl.scala 700:{40,40}]
  wire [4:0] _GEN_90366 = 5'h1d == _T_8999[4:0] ? 5'h0 : _GEN_90365; // @[FanCtrl.scala 700:{40,40}]
  wire [4:0] _GEN_90367 = 5'h1e == _T_8999[4:0] ? 5'h0 : _GEN_90366; // @[FanCtrl.scala 700:{40,40}]
  wire [4:0] _GEN_90368 = 5'h1f == _T_8999[4:0] ? 5'h0 : _GEN_90367; // @[FanCtrl.scala 700:{40,40}]
  wire [4:0] _GEN_90372 = 5'h3 == _T_9003[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 700:{40,40}]
  wire [4:0] _GEN_90373 = 5'h4 == _T_9003[4:0] ? w_vn_4 : _GEN_90372; // @[FanCtrl.scala 700:{40,40}]
  wire [4:0] _GEN_90374 = 5'h5 == _T_9003[4:0] ? 5'h0 : _GEN_90373; // @[FanCtrl.scala 700:{40,40}]
  wire [4:0] _GEN_90375 = 5'h6 == _T_9003[4:0] ? 5'h0 : _GEN_90374; // @[FanCtrl.scala 700:{40,40}]
  wire [4:0] _GEN_90376 = 5'h7 == _T_9003[4:0] ? w_vn_7 : _GEN_90375; // @[FanCtrl.scala 700:{40,40}]
  wire [4:0] _GEN_90377 = 5'h8 == _T_9003[4:0] ? w_vn_8 : _GEN_90376; // @[FanCtrl.scala 700:{40,40}]
  wire [4:0] _GEN_90378 = 5'h9 == _T_9003[4:0] ? 5'h0 : _GEN_90377; // @[FanCtrl.scala 700:{40,40}]
  wire [4:0] _GEN_90379 = 5'ha == _T_9003[4:0] ? 5'h0 : _GEN_90378; // @[FanCtrl.scala 700:{40,40}]
  wire [4:0] _GEN_90380 = 5'hb == _T_9003[4:0] ? w_vn_11 : _GEN_90379; // @[FanCtrl.scala 700:{40,40}]
  wire [4:0] _GEN_90381 = 5'hc == _T_9003[4:0] ? w_vn_12 : _GEN_90380; // @[FanCtrl.scala 700:{40,40}]
  wire [4:0] _GEN_90382 = 5'hd == _T_9003[4:0] ? w_vn_13 : _GEN_90381; // @[FanCtrl.scala 700:{40,40}]
  wire [4:0] _GEN_90383 = 5'he == _T_9003[4:0] ? 5'h0 : _GEN_90382; // @[FanCtrl.scala 700:{40,40}]
  wire [4:0] _GEN_90384 = 5'hf == _T_9003[4:0] ? w_vn_15 : _GEN_90383; // @[FanCtrl.scala 700:{40,40}]
  wire [4:0] _GEN_90385 = 5'h10 == _T_9003[4:0] ? w_vn_16 : _GEN_90384; // @[FanCtrl.scala 700:{40,40}]
  wire [4:0] _GEN_90386 = 5'h11 == _T_9003[4:0] ? 5'h0 : _GEN_90385; // @[FanCtrl.scala 700:{40,40}]
  wire [4:0] _GEN_90387 = 5'h12 == _T_9003[4:0] ? w_vn_18 : _GEN_90386; // @[FanCtrl.scala 700:{40,40}]
  wire [4:0] _GEN_90388 = 5'h13 == _T_9003[4:0] ? 5'h0 : _GEN_90387; // @[FanCtrl.scala 700:{40,40}]
  wire [4:0] _GEN_90389 = 5'h14 == _T_9003[4:0] ? 5'h0 : _GEN_90388; // @[FanCtrl.scala 700:{40,40}]
  wire [4:0] _GEN_90390 = 5'h15 == _T_9003[4:0] ? 5'h0 : _GEN_90389; // @[FanCtrl.scala 700:{40,40}]
  wire [4:0] _GEN_90391 = 5'h16 == _T_9003[4:0] ? 5'h0 : _GEN_90390; // @[FanCtrl.scala 700:{40,40}]
  wire [4:0] _GEN_90392 = 5'h17 == _T_9003[4:0] ? w_vn_23 : _GEN_90391; // @[FanCtrl.scala 700:{40,40}]
  wire [4:0] _GEN_90393 = 5'h18 == _T_9003[4:0] ? w_vn_24 : _GEN_90392; // @[FanCtrl.scala 700:{40,40}]
  wire [4:0] _GEN_90394 = 5'h19 == _T_9003[4:0] ? 5'h0 : _GEN_90393; // @[FanCtrl.scala 700:{40,40}]
  wire [4:0] _GEN_90395 = 5'h1a == _T_9003[4:0] ? 5'h0 : _GEN_90394; // @[FanCtrl.scala 700:{40,40}]
  wire [4:0] _GEN_90396 = 5'h1b == _T_9003[4:0] ? 5'h0 : _GEN_90395; // @[FanCtrl.scala 700:{40,40}]
  wire [4:0] _GEN_90397 = 5'h1c == _T_9003[4:0] ? 5'h0 : _GEN_90396; // @[FanCtrl.scala 700:{40,40}]
  wire [4:0] _GEN_90398 = 5'h1d == _T_9003[4:0] ? 5'h0 : _GEN_90397; // @[FanCtrl.scala 700:{40,40}]
  wire [4:0] _GEN_90399 = 5'h1e == _T_9003[4:0] ? 5'h0 : _GEN_90398; // @[FanCtrl.scala 700:{40,40}]
  wire [4:0] _GEN_90400 = 5'h1f == _T_9003[4:0] ? 5'h0 : _GEN_90399; // @[FanCtrl.scala 700:{40,40}]
  wire  _T_9005 = _GEN_90368 == _GEN_90400; // @[FanCtrl.scala 700:40]
  wire [6:0] _T_9012 = _T_8997 + 7'h7; // @[FanCtrl.scala 706:32]
  wire [6:0] _T_9016 = _T_8997 + 7'h8; // @[FanCtrl.scala 706:60]
  wire [4:0] _GEN_90497 = 5'h3 == _T_9012[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 706:{40,40}]
  wire [4:0] _GEN_90498 = 5'h4 == _T_9012[4:0] ? w_vn_4 : _GEN_90497; // @[FanCtrl.scala 706:{40,40}]
  wire [4:0] _GEN_90499 = 5'h5 == _T_9012[4:0] ? 5'h0 : _GEN_90498; // @[FanCtrl.scala 706:{40,40}]
  wire [4:0] _GEN_90500 = 5'h6 == _T_9012[4:0] ? 5'h0 : _GEN_90499; // @[FanCtrl.scala 706:{40,40}]
  wire [4:0] _GEN_90501 = 5'h7 == _T_9012[4:0] ? w_vn_7 : _GEN_90500; // @[FanCtrl.scala 706:{40,40}]
  wire [4:0] _GEN_90502 = 5'h8 == _T_9012[4:0] ? w_vn_8 : _GEN_90501; // @[FanCtrl.scala 706:{40,40}]
  wire [4:0] _GEN_90503 = 5'h9 == _T_9012[4:0] ? 5'h0 : _GEN_90502; // @[FanCtrl.scala 706:{40,40}]
  wire [4:0] _GEN_90504 = 5'ha == _T_9012[4:0] ? 5'h0 : _GEN_90503; // @[FanCtrl.scala 706:{40,40}]
  wire [4:0] _GEN_90505 = 5'hb == _T_9012[4:0] ? w_vn_11 : _GEN_90504; // @[FanCtrl.scala 706:{40,40}]
  wire [4:0] _GEN_90506 = 5'hc == _T_9012[4:0] ? w_vn_12 : _GEN_90505; // @[FanCtrl.scala 706:{40,40}]
  wire [4:0] _GEN_90507 = 5'hd == _T_9012[4:0] ? w_vn_13 : _GEN_90506; // @[FanCtrl.scala 706:{40,40}]
  wire [4:0] _GEN_90508 = 5'he == _T_9012[4:0] ? 5'h0 : _GEN_90507; // @[FanCtrl.scala 706:{40,40}]
  wire [4:0] _GEN_90509 = 5'hf == _T_9012[4:0] ? w_vn_15 : _GEN_90508; // @[FanCtrl.scala 706:{40,40}]
  wire [4:0] _GEN_90510 = 5'h10 == _T_9012[4:0] ? w_vn_16 : _GEN_90509; // @[FanCtrl.scala 706:{40,40}]
  wire [4:0] _GEN_90511 = 5'h11 == _T_9012[4:0] ? 5'h0 : _GEN_90510; // @[FanCtrl.scala 706:{40,40}]
  wire [4:0] _GEN_90512 = 5'h12 == _T_9012[4:0] ? w_vn_18 : _GEN_90511; // @[FanCtrl.scala 706:{40,40}]
  wire [4:0] _GEN_90513 = 5'h13 == _T_9012[4:0] ? 5'h0 : _GEN_90512; // @[FanCtrl.scala 706:{40,40}]
  wire [4:0] _GEN_90514 = 5'h14 == _T_9012[4:0] ? 5'h0 : _GEN_90513; // @[FanCtrl.scala 706:{40,40}]
  wire [4:0] _GEN_90515 = 5'h15 == _T_9012[4:0] ? 5'h0 : _GEN_90514; // @[FanCtrl.scala 706:{40,40}]
  wire [4:0] _GEN_90516 = 5'h16 == _T_9012[4:0] ? 5'h0 : _GEN_90515; // @[FanCtrl.scala 706:{40,40}]
  wire [4:0] _GEN_90517 = 5'h17 == _T_9012[4:0] ? w_vn_23 : _GEN_90516; // @[FanCtrl.scala 706:{40,40}]
  wire [4:0] _GEN_90518 = 5'h18 == _T_9012[4:0] ? w_vn_24 : _GEN_90517; // @[FanCtrl.scala 706:{40,40}]
  wire [4:0] _GEN_90519 = 5'h19 == _T_9012[4:0] ? 5'h0 : _GEN_90518; // @[FanCtrl.scala 706:{40,40}]
  wire [4:0] _GEN_90520 = 5'h1a == _T_9012[4:0] ? 5'h0 : _GEN_90519; // @[FanCtrl.scala 706:{40,40}]
  wire [4:0] _GEN_90521 = 5'h1b == _T_9012[4:0] ? 5'h0 : _GEN_90520; // @[FanCtrl.scala 706:{40,40}]
  wire [4:0] _GEN_90522 = 5'h1c == _T_9012[4:0] ? 5'h0 : _GEN_90521; // @[FanCtrl.scala 706:{40,40}]
  wire [4:0] _GEN_90523 = 5'h1d == _T_9012[4:0] ? 5'h0 : _GEN_90522; // @[FanCtrl.scala 706:{40,40}]
  wire [4:0] _GEN_90524 = 5'h1e == _T_9012[4:0] ? 5'h0 : _GEN_90523; // @[FanCtrl.scala 706:{40,40}]
  wire [4:0] _GEN_90525 = 5'h1f == _T_9012[4:0] ? 5'h0 : _GEN_90524; // @[FanCtrl.scala 706:{40,40}]
  wire [4:0] _GEN_90529 = 5'h3 == _T_9016[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 706:{40,40}]
  wire [4:0] _GEN_90530 = 5'h4 == _T_9016[4:0] ? w_vn_4 : _GEN_90529; // @[FanCtrl.scala 706:{40,40}]
  wire [4:0] _GEN_90531 = 5'h5 == _T_9016[4:0] ? 5'h0 : _GEN_90530; // @[FanCtrl.scala 706:{40,40}]
  wire [4:0] _GEN_90532 = 5'h6 == _T_9016[4:0] ? 5'h0 : _GEN_90531; // @[FanCtrl.scala 706:{40,40}]
  wire [4:0] _GEN_90533 = 5'h7 == _T_9016[4:0] ? w_vn_7 : _GEN_90532; // @[FanCtrl.scala 706:{40,40}]
  wire [4:0] _GEN_90534 = 5'h8 == _T_9016[4:0] ? w_vn_8 : _GEN_90533; // @[FanCtrl.scala 706:{40,40}]
  wire [4:0] _GEN_90535 = 5'h9 == _T_9016[4:0] ? 5'h0 : _GEN_90534; // @[FanCtrl.scala 706:{40,40}]
  wire [4:0] _GEN_90536 = 5'ha == _T_9016[4:0] ? 5'h0 : _GEN_90535; // @[FanCtrl.scala 706:{40,40}]
  wire [4:0] _GEN_90537 = 5'hb == _T_9016[4:0] ? w_vn_11 : _GEN_90536; // @[FanCtrl.scala 706:{40,40}]
  wire [4:0] _GEN_90538 = 5'hc == _T_9016[4:0] ? w_vn_12 : _GEN_90537; // @[FanCtrl.scala 706:{40,40}]
  wire [4:0] _GEN_90539 = 5'hd == _T_9016[4:0] ? w_vn_13 : _GEN_90538; // @[FanCtrl.scala 706:{40,40}]
  wire [4:0] _GEN_90540 = 5'he == _T_9016[4:0] ? 5'h0 : _GEN_90539; // @[FanCtrl.scala 706:{40,40}]
  wire [4:0] _GEN_90541 = 5'hf == _T_9016[4:0] ? w_vn_15 : _GEN_90540; // @[FanCtrl.scala 706:{40,40}]
  wire [4:0] _GEN_90542 = 5'h10 == _T_9016[4:0] ? w_vn_16 : _GEN_90541; // @[FanCtrl.scala 706:{40,40}]
  wire [4:0] _GEN_90543 = 5'h11 == _T_9016[4:0] ? 5'h0 : _GEN_90542; // @[FanCtrl.scala 706:{40,40}]
  wire [4:0] _GEN_90544 = 5'h12 == _T_9016[4:0] ? w_vn_18 : _GEN_90543; // @[FanCtrl.scala 706:{40,40}]
  wire [4:0] _GEN_90545 = 5'h13 == _T_9016[4:0] ? 5'h0 : _GEN_90544; // @[FanCtrl.scala 706:{40,40}]
  wire [4:0] _GEN_90546 = 5'h14 == _T_9016[4:0] ? 5'h0 : _GEN_90545; // @[FanCtrl.scala 706:{40,40}]
  wire [4:0] _GEN_90547 = 5'h15 == _T_9016[4:0] ? 5'h0 : _GEN_90546; // @[FanCtrl.scala 706:{40,40}]
  wire [4:0] _GEN_90548 = 5'h16 == _T_9016[4:0] ? 5'h0 : _GEN_90547; // @[FanCtrl.scala 706:{40,40}]
  wire [4:0] _GEN_90549 = 5'h17 == _T_9016[4:0] ? w_vn_23 : _GEN_90548; // @[FanCtrl.scala 706:{40,40}]
  wire [4:0] _GEN_90550 = 5'h18 == _T_9016[4:0] ? w_vn_24 : _GEN_90549; // @[FanCtrl.scala 706:{40,40}]
  wire [4:0] _GEN_90551 = 5'h19 == _T_9016[4:0] ? 5'h0 : _GEN_90550; // @[FanCtrl.scala 706:{40,40}]
  wire [4:0] _GEN_90552 = 5'h1a == _T_9016[4:0] ? 5'h0 : _GEN_90551; // @[FanCtrl.scala 706:{40,40}]
  wire [4:0] _GEN_90553 = 5'h1b == _T_9016[4:0] ? 5'h0 : _GEN_90552; // @[FanCtrl.scala 706:{40,40}]
  wire [4:0] _GEN_90554 = 5'h1c == _T_9016[4:0] ? 5'h0 : _GEN_90553; // @[FanCtrl.scala 706:{40,40}]
  wire [4:0] _GEN_90555 = 5'h1d == _T_9016[4:0] ? 5'h0 : _GEN_90554; // @[FanCtrl.scala 706:{40,40}]
  wire [4:0] _GEN_90556 = 5'h1e == _T_9016[4:0] ? 5'h0 : _GEN_90555; // @[FanCtrl.scala 706:{40,40}]
  wire [4:0] _GEN_90557 = 5'h1f == _T_9016[4:0] ? 5'h0 : _GEN_90556; // @[FanCtrl.scala 706:{40,40}]
  wire  _T_9018 = _GEN_90525 == _GEN_90557; // @[FanCtrl.scala 706:40]
  wire [6:0] _T_9021 = _T_8997 + 7'h17; // @[FanCtrl.scala 707:32]
  wire [6:0] _T_9025 = _T_8997 + 7'h18; // @[FanCtrl.scala 707:60]
  wire [4:0] _GEN_90561 = 5'h3 == _T_9021[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 707:{40,40}]
  wire [4:0] _GEN_90562 = 5'h4 == _T_9021[4:0] ? w_vn_4 : _GEN_90561; // @[FanCtrl.scala 707:{40,40}]
  wire [4:0] _GEN_90563 = 5'h5 == _T_9021[4:0] ? 5'h0 : _GEN_90562; // @[FanCtrl.scala 707:{40,40}]
  wire [4:0] _GEN_90564 = 5'h6 == _T_9021[4:0] ? 5'h0 : _GEN_90563; // @[FanCtrl.scala 707:{40,40}]
  wire [4:0] _GEN_90565 = 5'h7 == _T_9021[4:0] ? w_vn_7 : _GEN_90564; // @[FanCtrl.scala 707:{40,40}]
  wire [4:0] _GEN_90566 = 5'h8 == _T_9021[4:0] ? w_vn_8 : _GEN_90565; // @[FanCtrl.scala 707:{40,40}]
  wire [4:0] _GEN_90567 = 5'h9 == _T_9021[4:0] ? 5'h0 : _GEN_90566; // @[FanCtrl.scala 707:{40,40}]
  wire [4:0] _GEN_90568 = 5'ha == _T_9021[4:0] ? 5'h0 : _GEN_90567; // @[FanCtrl.scala 707:{40,40}]
  wire [4:0] _GEN_90569 = 5'hb == _T_9021[4:0] ? w_vn_11 : _GEN_90568; // @[FanCtrl.scala 707:{40,40}]
  wire [4:0] _GEN_90570 = 5'hc == _T_9021[4:0] ? w_vn_12 : _GEN_90569; // @[FanCtrl.scala 707:{40,40}]
  wire [4:0] _GEN_90571 = 5'hd == _T_9021[4:0] ? w_vn_13 : _GEN_90570; // @[FanCtrl.scala 707:{40,40}]
  wire [4:0] _GEN_90572 = 5'he == _T_9021[4:0] ? 5'h0 : _GEN_90571; // @[FanCtrl.scala 707:{40,40}]
  wire [4:0] _GEN_90573 = 5'hf == _T_9021[4:0] ? w_vn_15 : _GEN_90572; // @[FanCtrl.scala 707:{40,40}]
  wire [4:0] _GEN_90574 = 5'h10 == _T_9021[4:0] ? w_vn_16 : _GEN_90573; // @[FanCtrl.scala 707:{40,40}]
  wire [4:0] _GEN_90575 = 5'h11 == _T_9021[4:0] ? 5'h0 : _GEN_90574; // @[FanCtrl.scala 707:{40,40}]
  wire [4:0] _GEN_90576 = 5'h12 == _T_9021[4:0] ? w_vn_18 : _GEN_90575; // @[FanCtrl.scala 707:{40,40}]
  wire [4:0] _GEN_90577 = 5'h13 == _T_9021[4:0] ? 5'h0 : _GEN_90576; // @[FanCtrl.scala 707:{40,40}]
  wire [4:0] _GEN_90578 = 5'h14 == _T_9021[4:0] ? 5'h0 : _GEN_90577; // @[FanCtrl.scala 707:{40,40}]
  wire [4:0] _GEN_90579 = 5'h15 == _T_9021[4:0] ? 5'h0 : _GEN_90578; // @[FanCtrl.scala 707:{40,40}]
  wire [4:0] _GEN_90580 = 5'h16 == _T_9021[4:0] ? 5'h0 : _GEN_90579; // @[FanCtrl.scala 707:{40,40}]
  wire [4:0] _GEN_90581 = 5'h17 == _T_9021[4:0] ? w_vn_23 : _GEN_90580; // @[FanCtrl.scala 707:{40,40}]
  wire [4:0] _GEN_90582 = 5'h18 == _T_9021[4:0] ? w_vn_24 : _GEN_90581; // @[FanCtrl.scala 707:{40,40}]
  wire [4:0] _GEN_90583 = 5'h19 == _T_9021[4:0] ? 5'h0 : _GEN_90582; // @[FanCtrl.scala 707:{40,40}]
  wire [4:0] _GEN_90584 = 5'h1a == _T_9021[4:0] ? 5'h0 : _GEN_90583; // @[FanCtrl.scala 707:{40,40}]
  wire [4:0] _GEN_90585 = 5'h1b == _T_9021[4:0] ? 5'h0 : _GEN_90584; // @[FanCtrl.scala 707:{40,40}]
  wire [4:0] _GEN_90586 = 5'h1c == _T_9021[4:0] ? 5'h0 : _GEN_90585; // @[FanCtrl.scala 707:{40,40}]
  wire [4:0] _GEN_90587 = 5'h1d == _T_9021[4:0] ? 5'h0 : _GEN_90586; // @[FanCtrl.scala 707:{40,40}]
  wire [4:0] _GEN_90588 = 5'h1e == _T_9021[4:0] ? 5'h0 : _GEN_90587; // @[FanCtrl.scala 707:{40,40}]
  wire [4:0] _GEN_90589 = 5'h1f == _T_9021[4:0] ? 5'h0 : _GEN_90588; // @[FanCtrl.scala 707:{40,40}]
  wire [4:0] _GEN_90593 = 5'h3 == _T_9025[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 707:{40,40}]
  wire [4:0] _GEN_90594 = 5'h4 == _T_9025[4:0] ? w_vn_4 : _GEN_90593; // @[FanCtrl.scala 707:{40,40}]
  wire [4:0] _GEN_90595 = 5'h5 == _T_9025[4:0] ? 5'h0 : _GEN_90594; // @[FanCtrl.scala 707:{40,40}]
  wire [4:0] _GEN_90596 = 5'h6 == _T_9025[4:0] ? 5'h0 : _GEN_90595; // @[FanCtrl.scala 707:{40,40}]
  wire [4:0] _GEN_90597 = 5'h7 == _T_9025[4:0] ? w_vn_7 : _GEN_90596; // @[FanCtrl.scala 707:{40,40}]
  wire [4:0] _GEN_90598 = 5'h8 == _T_9025[4:0] ? w_vn_8 : _GEN_90597; // @[FanCtrl.scala 707:{40,40}]
  wire [4:0] _GEN_90599 = 5'h9 == _T_9025[4:0] ? 5'h0 : _GEN_90598; // @[FanCtrl.scala 707:{40,40}]
  wire [4:0] _GEN_90600 = 5'ha == _T_9025[4:0] ? 5'h0 : _GEN_90599; // @[FanCtrl.scala 707:{40,40}]
  wire [4:0] _GEN_90601 = 5'hb == _T_9025[4:0] ? w_vn_11 : _GEN_90600; // @[FanCtrl.scala 707:{40,40}]
  wire [4:0] _GEN_90602 = 5'hc == _T_9025[4:0] ? w_vn_12 : _GEN_90601; // @[FanCtrl.scala 707:{40,40}]
  wire [4:0] _GEN_90603 = 5'hd == _T_9025[4:0] ? w_vn_13 : _GEN_90602; // @[FanCtrl.scala 707:{40,40}]
  wire [4:0] _GEN_90604 = 5'he == _T_9025[4:0] ? 5'h0 : _GEN_90603; // @[FanCtrl.scala 707:{40,40}]
  wire [4:0] _GEN_90605 = 5'hf == _T_9025[4:0] ? w_vn_15 : _GEN_90604; // @[FanCtrl.scala 707:{40,40}]
  wire [4:0] _GEN_90606 = 5'h10 == _T_9025[4:0] ? w_vn_16 : _GEN_90605; // @[FanCtrl.scala 707:{40,40}]
  wire [4:0] _GEN_90607 = 5'h11 == _T_9025[4:0] ? 5'h0 : _GEN_90606; // @[FanCtrl.scala 707:{40,40}]
  wire [4:0] _GEN_90608 = 5'h12 == _T_9025[4:0] ? w_vn_18 : _GEN_90607; // @[FanCtrl.scala 707:{40,40}]
  wire [4:0] _GEN_90609 = 5'h13 == _T_9025[4:0] ? 5'h0 : _GEN_90608; // @[FanCtrl.scala 707:{40,40}]
  wire [4:0] _GEN_90610 = 5'h14 == _T_9025[4:0] ? 5'h0 : _GEN_90609; // @[FanCtrl.scala 707:{40,40}]
  wire [4:0] _GEN_90611 = 5'h15 == _T_9025[4:0] ? 5'h0 : _GEN_90610; // @[FanCtrl.scala 707:{40,40}]
  wire [4:0] _GEN_90612 = 5'h16 == _T_9025[4:0] ? 5'h0 : _GEN_90611; // @[FanCtrl.scala 707:{40,40}]
  wire [4:0] _GEN_90613 = 5'h17 == _T_9025[4:0] ? w_vn_23 : _GEN_90612; // @[FanCtrl.scala 707:{40,40}]
  wire [4:0] _GEN_90614 = 5'h18 == _T_9025[4:0] ? w_vn_24 : _GEN_90613; // @[FanCtrl.scala 707:{40,40}]
  wire [4:0] _GEN_90615 = 5'h19 == _T_9025[4:0] ? 5'h0 : _GEN_90614; // @[FanCtrl.scala 707:{40,40}]
  wire [4:0] _GEN_90616 = 5'h1a == _T_9025[4:0] ? 5'h0 : _GEN_90615; // @[FanCtrl.scala 707:{40,40}]
  wire [4:0] _GEN_90617 = 5'h1b == _T_9025[4:0] ? 5'h0 : _GEN_90616; // @[FanCtrl.scala 707:{40,40}]
  wire [4:0] _GEN_90618 = 5'h1c == _T_9025[4:0] ? 5'h0 : _GEN_90617; // @[FanCtrl.scala 707:{40,40}]
  wire [4:0] _GEN_90619 = 5'h1d == _T_9025[4:0] ? 5'h0 : _GEN_90618; // @[FanCtrl.scala 707:{40,40}]
  wire [4:0] _GEN_90620 = 5'h1e == _T_9025[4:0] ? 5'h0 : _GEN_90619; // @[FanCtrl.scala 707:{40,40}]
  wire [4:0] _GEN_90621 = 5'h1f == _T_9025[4:0] ? 5'h0 : _GEN_90620; // @[FanCtrl.scala 707:{40,40}]
  wire  _T_9027 = _GEN_90589 == _GEN_90621; // @[FanCtrl.scala 707:40]
  wire  _T_9028 = _GEN_90525 == _GEN_90557 & _T_9027; // @[FanCtrl.scala 706:69]
  wire  _T_9037 = _GEN_90557 != _GEN_90400; // @[FanCtrl.scala 708:39]
  wire  _T_9038 = _T_9028 & _T_9037; // @[FanCtrl.scala 707:69]
  wire  _T_9047 = _GEN_90589 != _GEN_90368; // @[FanCtrl.scala 709:41]
  wire  _T_9048 = _T_9038 & _T_9047; // @[FanCtrl.scala 708:69]
  wire  _T_9069 = _T_9027 & _T_9047; // @[FanCtrl.scala 713:77]
  wire  _T_9089 = _GEN_90400 != _GEN_90557; // @[FanCtrl.scala 719:45]
  wire  _T_9090 = _T_9018 & _T_9089; // @[FanCtrl.scala 718:75]
  wire [2:0] _GEN_91160 = _T_9090 ? 3'h3 : 3'h0; // @[FanCtrl.scala 719:75]
  wire  _GEN_91315 = r_valid_1 & _T_9005; // @[FanCtrl.scala 699:36]
  wire [1:0] _GEN_91411 = 5'h0 == _T_8995 ? 2'h0 : _GEN_90317; // @[FanCtrl.scala 733:{47,47}]
  wire [1:0] _GEN_91412 = 5'h1 == _T_8995 ? 2'h0 : _GEN_90318; // @[FanCtrl.scala 733:{47,47}]
  wire [1:0] _GEN_91413 = 5'h2 == _T_8995 ? 2'h0 : _GEN_90319; // @[FanCtrl.scala 733:{47,47}]
  wire [1:0] _GEN_91414 = 5'h3 == _T_8995 ? 2'h0 : _GEN_90320; // @[FanCtrl.scala 733:{47,47}]
  wire [1:0] _GEN_91415 = 5'h4 == _T_8995 ? 2'h0 : _GEN_90321; // @[FanCtrl.scala 733:{47,47}]
  wire [1:0] _GEN_91416 = 5'h5 == _T_8995 ? 2'h0 : _GEN_90322; // @[FanCtrl.scala 733:{47,47}]
  wire [1:0] _GEN_91417 = 5'h6 == _T_8995 ? 2'h0 : _GEN_90323; // @[FanCtrl.scala 733:{47,47}]
  wire [1:0] _GEN_91418 = 5'h7 == _T_8995 ? 2'h0 : _GEN_90324; // @[FanCtrl.scala 733:{47,47}]
  wire [1:0] _GEN_91419 = 5'h8 == _T_8995 ? 2'h0 : _GEN_90325; // @[FanCtrl.scala 733:{47,47}]
  wire [1:0] _GEN_91420 = 5'h9 == _T_8995 ? 2'h0 : _GEN_90326; // @[FanCtrl.scala 733:{47,47}]
  wire [1:0] _GEN_91421 = 5'ha == _T_8995 ? 2'h0 : _GEN_90327; // @[FanCtrl.scala 733:{47,47}]
  wire [1:0] _GEN_91422 = 5'hb == _T_8995 ? 2'h0 : _GEN_90328; // @[FanCtrl.scala 733:{47,47}]
  wire [1:0] _GEN_91423 = 5'hc == _T_8995 ? 2'h0 : _GEN_90329; // @[FanCtrl.scala 733:{47,47}]
  wire [1:0] _GEN_91424 = 5'hd == _T_8995 ? 2'h0 : _GEN_90330; // @[FanCtrl.scala 733:{47,47}]
  wire [1:0] _GEN_91425 = 5'he == _T_8995 ? 2'h0 : _GEN_90331; // @[FanCtrl.scala 733:{47,47}]
  wire [1:0] _GEN_91426 = 5'hf == _T_8995 ? 2'h0 : _GEN_90332; // @[FanCtrl.scala 733:{47,47}]
  wire [1:0] _GEN_91427 = 5'h10 == _T_8995 ? 2'h0 : _GEN_90333; // @[FanCtrl.scala 733:{47,47}]
  wire [1:0] _GEN_91428 = 5'h11 == _T_8995 ? 2'h0 : _GEN_90334; // @[FanCtrl.scala 733:{47,47}]
  wire [1:0] _GEN_91429 = 5'h12 == _T_8995 ? 2'h0 : _GEN_90335; // @[FanCtrl.scala 733:{47,47}]
  wire [1:0] _GEN_91430 = 5'h13 == _T_8995 ? 2'h0 : _GEN_90336; // @[FanCtrl.scala 733:{47,47}]
  wire [6:0] _T_9118 = _T_8997 + 7'hb; // @[FanCtrl.scala 734:67]
  wire [4:0] _GEN_91466 = 5'h3 == _T_9118[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 734:{47,47}]
  wire [4:0] _GEN_91467 = 5'h4 == _T_9118[4:0] ? w_vn_4 : _GEN_91466; // @[FanCtrl.scala 734:{47,47}]
  wire [4:0] _GEN_91468 = 5'h5 == _T_9118[4:0] ? 5'h0 : _GEN_91467; // @[FanCtrl.scala 734:{47,47}]
  wire [4:0] _GEN_91469 = 5'h6 == _T_9118[4:0] ? 5'h0 : _GEN_91468; // @[FanCtrl.scala 734:{47,47}]
  wire [4:0] _GEN_91470 = 5'h7 == _T_9118[4:0] ? w_vn_7 : _GEN_91469; // @[FanCtrl.scala 734:{47,47}]
  wire [4:0] _GEN_91471 = 5'h8 == _T_9118[4:0] ? w_vn_8 : _GEN_91470; // @[FanCtrl.scala 734:{47,47}]
  wire [4:0] _GEN_91472 = 5'h9 == _T_9118[4:0] ? 5'h0 : _GEN_91471; // @[FanCtrl.scala 734:{47,47}]
  wire [4:0] _GEN_91473 = 5'ha == _T_9118[4:0] ? 5'h0 : _GEN_91472; // @[FanCtrl.scala 734:{47,47}]
  wire [4:0] _GEN_91474 = 5'hb == _T_9118[4:0] ? w_vn_11 : _GEN_91473; // @[FanCtrl.scala 734:{47,47}]
  wire [4:0] _GEN_91475 = 5'hc == _T_9118[4:0] ? w_vn_12 : _GEN_91474; // @[FanCtrl.scala 734:{47,47}]
  wire [4:0] _GEN_91476 = 5'hd == _T_9118[4:0] ? w_vn_13 : _GEN_91475; // @[FanCtrl.scala 734:{47,47}]
  wire [4:0] _GEN_91477 = 5'he == _T_9118[4:0] ? 5'h0 : _GEN_91476; // @[FanCtrl.scala 734:{47,47}]
  wire [4:0] _GEN_91478 = 5'hf == _T_9118[4:0] ? w_vn_15 : _GEN_91477; // @[FanCtrl.scala 734:{47,47}]
  wire [4:0] _GEN_91479 = 5'h10 == _T_9118[4:0] ? w_vn_16 : _GEN_91478; // @[FanCtrl.scala 734:{47,47}]
  wire [4:0] _GEN_91480 = 5'h11 == _T_9118[4:0] ? 5'h0 : _GEN_91479; // @[FanCtrl.scala 734:{47,47}]
  wire [4:0] _GEN_91481 = 5'h12 == _T_9118[4:0] ? w_vn_18 : _GEN_91480; // @[FanCtrl.scala 734:{47,47}]
  wire [4:0] _GEN_91482 = 5'h13 == _T_9118[4:0] ? 5'h0 : _GEN_91481; // @[FanCtrl.scala 734:{47,47}]
  wire [4:0] _GEN_91483 = 5'h14 == _T_9118[4:0] ? 5'h0 : _GEN_91482; // @[FanCtrl.scala 734:{47,47}]
  wire [4:0] _GEN_91484 = 5'h15 == _T_9118[4:0] ? 5'h0 : _GEN_91483; // @[FanCtrl.scala 734:{47,47}]
  wire [4:0] _GEN_91485 = 5'h16 == _T_9118[4:0] ? 5'h0 : _GEN_91484; // @[FanCtrl.scala 734:{47,47}]
  wire [4:0] _GEN_91486 = 5'h17 == _T_9118[4:0] ? w_vn_23 : _GEN_91485; // @[FanCtrl.scala 734:{47,47}]
  wire [4:0] _GEN_91487 = 5'h18 == _T_9118[4:0] ? w_vn_24 : _GEN_91486; // @[FanCtrl.scala 734:{47,47}]
  wire [4:0] _GEN_91488 = 5'h19 == _T_9118[4:0] ? 5'h0 : _GEN_91487; // @[FanCtrl.scala 734:{47,47}]
  wire [4:0] _GEN_91489 = 5'h1a == _T_9118[4:0] ? 5'h0 : _GEN_91488; // @[FanCtrl.scala 734:{47,47}]
  wire [4:0] _GEN_91490 = 5'h1b == _T_9118[4:0] ? 5'h0 : _GEN_91489; // @[FanCtrl.scala 734:{47,47}]
  wire [4:0] _GEN_91491 = 5'h1c == _T_9118[4:0] ? 5'h0 : _GEN_91490; // @[FanCtrl.scala 734:{47,47}]
  wire [4:0] _GEN_91492 = 5'h1d == _T_9118[4:0] ? 5'h0 : _GEN_91491; // @[FanCtrl.scala 734:{47,47}]
  wire [4:0] _GEN_91493 = 5'h1e == _T_9118[4:0] ? 5'h0 : _GEN_91492; // @[FanCtrl.scala 734:{47,47}]
  wire [4:0] _GEN_91494 = 5'h1f == _T_9118[4:0] ? 5'h0 : _GEN_91493; // @[FanCtrl.scala 734:{47,47}]
  wire [1:0] _GEN_91495 = 5'h0 == _T_8995 ? 2'h1 : _GEN_90317; // @[FanCtrl.scala 735:{47,47}]
  wire [1:0] _GEN_91496 = 5'h1 == _T_8995 ? 2'h1 : _GEN_90318; // @[FanCtrl.scala 735:{47,47}]
  wire [1:0] _GEN_91497 = 5'h2 == _T_8995 ? 2'h1 : _GEN_90319; // @[FanCtrl.scala 735:{47,47}]
  wire [1:0] _GEN_91498 = 5'h3 == _T_8995 ? 2'h1 : _GEN_90320; // @[FanCtrl.scala 735:{47,47}]
  wire [1:0] _GEN_91499 = 5'h4 == _T_8995 ? 2'h1 : _GEN_90321; // @[FanCtrl.scala 735:{47,47}]
  wire [1:0] _GEN_91500 = 5'h5 == _T_8995 ? 2'h1 : _GEN_90322; // @[FanCtrl.scala 735:{47,47}]
  wire [1:0] _GEN_91501 = 5'h6 == _T_8995 ? 2'h1 : _GEN_90323; // @[FanCtrl.scala 735:{47,47}]
  wire [1:0] _GEN_91502 = 5'h7 == _T_8995 ? 2'h1 : _GEN_90324; // @[FanCtrl.scala 735:{47,47}]
  wire [1:0] _GEN_91503 = 5'h8 == _T_8995 ? 2'h1 : _GEN_90325; // @[FanCtrl.scala 735:{47,47}]
  wire [1:0] _GEN_91504 = 5'h9 == _T_8995 ? 2'h1 : _GEN_90326; // @[FanCtrl.scala 735:{47,47}]
  wire [1:0] _GEN_91505 = 5'ha == _T_8995 ? 2'h1 : _GEN_90327; // @[FanCtrl.scala 735:{47,47}]
  wire [1:0] _GEN_91506 = 5'hb == _T_8995 ? 2'h1 : _GEN_90328; // @[FanCtrl.scala 735:{47,47}]
  wire [1:0] _GEN_91507 = 5'hc == _T_8995 ? 2'h1 : _GEN_90329; // @[FanCtrl.scala 735:{47,47}]
  wire [1:0] _GEN_91508 = 5'hd == _T_8995 ? 2'h1 : _GEN_90330; // @[FanCtrl.scala 735:{47,47}]
  wire [1:0] _GEN_91509 = 5'he == _T_8995 ? 2'h1 : _GEN_90331; // @[FanCtrl.scala 735:{47,47}]
  wire [1:0] _GEN_91510 = 5'hf == _T_8995 ? 2'h1 : _GEN_90332; // @[FanCtrl.scala 735:{47,47}]
  wire [1:0] _GEN_91511 = 5'h10 == _T_8995 ? 2'h1 : _GEN_90333; // @[FanCtrl.scala 735:{47,47}]
  wire [1:0] _GEN_91512 = 5'h11 == _T_8995 ? 2'h1 : _GEN_90334; // @[FanCtrl.scala 735:{47,47}]
  wire [1:0] _GEN_91513 = 5'h12 == _T_8995 ? 2'h1 : _GEN_90335; // @[FanCtrl.scala 735:{47,47}]
  wire [1:0] _GEN_91514 = 5'h13 == _T_8995 ? 2'h1 : _GEN_90336; // @[FanCtrl.scala 735:{47,47}]
  wire [6:0] _T_9130 = _T_8997 + 7'hd; // @[FanCtrl.scala 736:67]
  wire [4:0] _GEN_91550 = 5'h3 == _T_9130[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 736:{47,47}]
  wire [4:0] _GEN_91551 = 5'h4 == _T_9130[4:0] ? w_vn_4 : _GEN_91550; // @[FanCtrl.scala 736:{47,47}]
  wire [4:0] _GEN_91552 = 5'h5 == _T_9130[4:0] ? 5'h0 : _GEN_91551; // @[FanCtrl.scala 736:{47,47}]
  wire [4:0] _GEN_91553 = 5'h6 == _T_9130[4:0] ? 5'h0 : _GEN_91552; // @[FanCtrl.scala 736:{47,47}]
  wire [4:0] _GEN_91554 = 5'h7 == _T_9130[4:0] ? w_vn_7 : _GEN_91553; // @[FanCtrl.scala 736:{47,47}]
  wire [4:0] _GEN_91555 = 5'h8 == _T_9130[4:0] ? w_vn_8 : _GEN_91554; // @[FanCtrl.scala 736:{47,47}]
  wire [4:0] _GEN_91556 = 5'h9 == _T_9130[4:0] ? 5'h0 : _GEN_91555; // @[FanCtrl.scala 736:{47,47}]
  wire [4:0] _GEN_91557 = 5'ha == _T_9130[4:0] ? 5'h0 : _GEN_91556; // @[FanCtrl.scala 736:{47,47}]
  wire [4:0] _GEN_91558 = 5'hb == _T_9130[4:0] ? w_vn_11 : _GEN_91557; // @[FanCtrl.scala 736:{47,47}]
  wire [4:0] _GEN_91559 = 5'hc == _T_9130[4:0] ? w_vn_12 : _GEN_91558; // @[FanCtrl.scala 736:{47,47}]
  wire [4:0] _GEN_91560 = 5'hd == _T_9130[4:0] ? w_vn_13 : _GEN_91559; // @[FanCtrl.scala 736:{47,47}]
  wire [4:0] _GEN_91561 = 5'he == _T_9130[4:0] ? 5'h0 : _GEN_91560; // @[FanCtrl.scala 736:{47,47}]
  wire [4:0] _GEN_91562 = 5'hf == _T_9130[4:0] ? w_vn_15 : _GEN_91561; // @[FanCtrl.scala 736:{47,47}]
  wire [4:0] _GEN_91563 = 5'h10 == _T_9130[4:0] ? w_vn_16 : _GEN_91562; // @[FanCtrl.scala 736:{47,47}]
  wire [4:0] _GEN_91564 = 5'h11 == _T_9130[4:0] ? 5'h0 : _GEN_91563; // @[FanCtrl.scala 736:{47,47}]
  wire [4:0] _GEN_91565 = 5'h12 == _T_9130[4:0] ? w_vn_18 : _GEN_91564; // @[FanCtrl.scala 736:{47,47}]
  wire [4:0] _GEN_91566 = 5'h13 == _T_9130[4:0] ? 5'h0 : _GEN_91565; // @[FanCtrl.scala 736:{47,47}]
  wire [4:0] _GEN_91567 = 5'h14 == _T_9130[4:0] ? 5'h0 : _GEN_91566; // @[FanCtrl.scala 736:{47,47}]
  wire [4:0] _GEN_91568 = 5'h15 == _T_9130[4:0] ? 5'h0 : _GEN_91567; // @[FanCtrl.scala 736:{47,47}]
  wire [4:0] _GEN_91569 = 5'h16 == _T_9130[4:0] ? 5'h0 : _GEN_91568; // @[FanCtrl.scala 736:{47,47}]
  wire [4:0] _GEN_91570 = 5'h17 == _T_9130[4:0] ? w_vn_23 : _GEN_91569; // @[FanCtrl.scala 736:{47,47}]
  wire [4:0] _GEN_91571 = 5'h18 == _T_9130[4:0] ? w_vn_24 : _GEN_91570; // @[FanCtrl.scala 736:{47,47}]
  wire [4:0] _GEN_91572 = 5'h19 == _T_9130[4:0] ? 5'h0 : _GEN_91571; // @[FanCtrl.scala 736:{47,47}]
  wire [4:0] _GEN_91573 = 5'h1a == _T_9130[4:0] ? 5'h0 : _GEN_91572; // @[FanCtrl.scala 736:{47,47}]
  wire [4:0] _GEN_91574 = 5'h1b == _T_9130[4:0] ? 5'h0 : _GEN_91573; // @[FanCtrl.scala 736:{47,47}]
  wire [4:0] _GEN_91575 = 5'h1c == _T_9130[4:0] ? 5'h0 : _GEN_91574; // @[FanCtrl.scala 736:{47,47}]
  wire [4:0] _GEN_91576 = 5'h1d == _T_9130[4:0] ? 5'h0 : _GEN_91575; // @[FanCtrl.scala 736:{47,47}]
  wire [4:0] _GEN_91577 = 5'h1e == _T_9130[4:0] ? 5'h0 : _GEN_91576; // @[FanCtrl.scala 736:{47,47}]
  wire [4:0] _GEN_91578 = 5'h1f == _T_9130[4:0] ? 5'h0 : _GEN_91577; // @[FanCtrl.scala 736:{47,47}]
  wire [1:0] _GEN_91579 = 5'h0 == _T_8995 ? 2'h2 : _GEN_90317; // @[FanCtrl.scala 737:{47,47}]
  wire [1:0] _GEN_91580 = 5'h1 == _T_8995 ? 2'h2 : _GEN_90318; // @[FanCtrl.scala 737:{47,47}]
  wire [1:0] _GEN_91581 = 5'h2 == _T_8995 ? 2'h2 : _GEN_90319; // @[FanCtrl.scala 737:{47,47}]
  wire [1:0] _GEN_91582 = 5'h3 == _T_8995 ? 2'h2 : _GEN_90320; // @[FanCtrl.scala 737:{47,47}]
  wire [1:0] _GEN_91583 = 5'h4 == _T_8995 ? 2'h2 : _GEN_90321; // @[FanCtrl.scala 737:{47,47}]
  wire [1:0] _GEN_91584 = 5'h5 == _T_8995 ? 2'h2 : _GEN_90322; // @[FanCtrl.scala 737:{47,47}]
  wire [1:0] _GEN_91585 = 5'h6 == _T_8995 ? 2'h2 : _GEN_90323; // @[FanCtrl.scala 737:{47,47}]
  wire [1:0] _GEN_91586 = 5'h7 == _T_8995 ? 2'h2 : _GEN_90324; // @[FanCtrl.scala 737:{47,47}]
  wire [1:0] _GEN_91587 = 5'h8 == _T_8995 ? 2'h2 : _GEN_90325; // @[FanCtrl.scala 737:{47,47}]
  wire [1:0] _GEN_91588 = 5'h9 == _T_8995 ? 2'h2 : _GEN_90326; // @[FanCtrl.scala 737:{47,47}]
  wire [1:0] _GEN_91589 = 5'ha == _T_8995 ? 2'h2 : _GEN_90327; // @[FanCtrl.scala 737:{47,47}]
  wire [1:0] _GEN_91590 = 5'hb == _T_8995 ? 2'h2 : _GEN_90328; // @[FanCtrl.scala 737:{47,47}]
  wire [1:0] _GEN_91591 = 5'hc == _T_8995 ? 2'h2 : _GEN_90329; // @[FanCtrl.scala 737:{47,47}]
  wire [1:0] _GEN_91592 = 5'hd == _T_8995 ? 2'h2 : _GEN_90330; // @[FanCtrl.scala 737:{47,47}]
  wire [1:0] _GEN_91593 = 5'he == _T_8995 ? 2'h2 : _GEN_90331; // @[FanCtrl.scala 737:{47,47}]
  wire [1:0] _GEN_91594 = 5'hf == _T_8995 ? 2'h2 : _GEN_90332; // @[FanCtrl.scala 737:{47,47}]
  wire [1:0] _GEN_91595 = 5'h10 == _T_8995 ? 2'h2 : _GEN_90333; // @[FanCtrl.scala 737:{47,47}]
  wire [1:0] _GEN_91596 = 5'h11 == _T_8995 ? 2'h2 : _GEN_90334; // @[FanCtrl.scala 737:{47,47}]
  wire [1:0] _GEN_91597 = 5'h12 == _T_8995 ? 2'h2 : _GEN_90335; // @[FanCtrl.scala 737:{47,47}]
  wire [1:0] _GEN_91598 = 5'h13 == _T_8995 ? 2'h2 : _GEN_90336; // @[FanCtrl.scala 737:{47,47}]
  wire [1:0] _GEN_91599 = 5'h0 == _T_8995 ? 2'h3 : _GEN_90317; // @[FanCtrl.scala 739:{47,47}]
  wire [1:0] _GEN_91600 = 5'h1 == _T_8995 ? 2'h3 : _GEN_90318; // @[FanCtrl.scala 739:{47,47}]
  wire [1:0] _GEN_91601 = 5'h2 == _T_8995 ? 2'h3 : _GEN_90319; // @[FanCtrl.scala 739:{47,47}]
  wire [1:0] _GEN_91602 = 5'h3 == _T_8995 ? 2'h3 : _GEN_90320; // @[FanCtrl.scala 739:{47,47}]
  wire [1:0] _GEN_91603 = 5'h4 == _T_8995 ? 2'h3 : _GEN_90321; // @[FanCtrl.scala 739:{47,47}]
  wire [1:0] _GEN_91604 = 5'h5 == _T_8995 ? 2'h3 : _GEN_90322; // @[FanCtrl.scala 739:{47,47}]
  wire [1:0] _GEN_91605 = 5'h6 == _T_8995 ? 2'h3 : _GEN_90323; // @[FanCtrl.scala 739:{47,47}]
  wire [1:0] _GEN_91606 = 5'h7 == _T_8995 ? 2'h3 : _GEN_90324; // @[FanCtrl.scala 739:{47,47}]
  wire [1:0] _GEN_91607 = 5'h8 == _T_8995 ? 2'h3 : _GEN_90325; // @[FanCtrl.scala 739:{47,47}]
  wire [1:0] _GEN_91608 = 5'h9 == _T_8995 ? 2'h3 : _GEN_90326; // @[FanCtrl.scala 739:{47,47}]
  wire [1:0] _GEN_91609 = 5'ha == _T_8995 ? 2'h3 : _GEN_90327; // @[FanCtrl.scala 739:{47,47}]
  wire [1:0] _GEN_91610 = 5'hb == _T_8995 ? 2'h3 : _GEN_90328; // @[FanCtrl.scala 739:{47,47}]
  wire [1:0] _GEN_91611 = 5'hc == _T_8995 ? 2'h3 : _GEN_90329; // @[FanCtrl.scala 739:{47,47}]
  wire [1:0] _GEN_91612 = 5'hd == _T_8995 ? 2'h3 : _GEN_90330; // @[FanCtrl.scala 739:{47,47}]
  wire [1:0] _GEN_91613 = 5'he == _T_8995 ? 2'h3 : _GEN_90331; // @[FanCtrl.scala 739:{47,47}]
  wire [1:0] _GEN_91614 = 5'hf == _T_8995 ? 2'h3 : _GEN_90332; // @[FanCtrl.scala 739:{47,47}]
  wire [1:0] _GEN_91615 = 5'h10 == _T_8995 ? 2'h3 : _GEN_90333; // @[FanCtrl.scala 739:{47,47}]
  wire [1:0] _GEN_91616 = 5'h11 == _T_8995 ? 2'h3 : _GEN_90334; // @[FanCtrl.scala 739:{47,47}]
  wire [1:0] _GEN_91617 = 5'h12 == _T_8995 ? 2'h3 : _GEN_90335; // @[FanCtrl.scala 739:{47,47}]
  wire [1:0] _GEN_91618 = 5'h13 == _T_8995 ? 2'h3 : _GEN_90336; // @[FanCtrl.scala 739:{47,47}]
  wire [1:0] _GEN_91619 = _GEN_90368 == _GEN_91578 ? _GEN_91579 : _GEN_91599; // @[FanCtrl.scala 736:76]
  wire [1:0] _GEN_91620 = _GEN_90368 == _GEN_91578 ? _GEN_91580 : _GEN_91600; // @[FanCtrl.scala 736:76]
  wire [1:0] _GEN_91621 = _GEN_90368 == _GEN_91578 ? _GEN_91581 : _GEN_91601; // @[FanCtrl.scala 736:76]
  wire [1:0] _GEN_91622 = _GEN_90368 == _GEN_91578 ? _GEN_91582 : _GEN_91602; // @[FanCtrl.scala 736:76]
  wire [1:0] _GEN_91623 = _GEN_90368 == _GEN_91578 ? _GEN_91583 : _GEN_91603; // @[FanCtrl.scala 736:76]
  wire [1:0] _GEN_91624 = _GEN_90368 == _GEN_91578 ? _GEN_91584 : _GEN_91604; // @[FanCtrl.scala 736:76]
  wire [1:0] _GEN_91625 = _GEN_90368 == _GEN_91578 ? _GEN_91585 : _GEN_91605; // @[FanCtrl.scala 736:76]
  wire [1:0] _GEN_91626 = _GEN_90368 == _GEN_91578 ? _GEN_91586 : _GEN_91606; // @[FanCtrl.scala 736:76]
  wire [1:0] _GEN_91627 = _GEN_90368 == _GEN_91578 ? _GEN_91587 : _GEN_91607; // @[FanCtrl.scala 736:76]
  wire [1:0] _GEN_91628 = _GEN_90368 == _GEN_91578 ? _GEN_91588 : _GEN_91608; // @[FanCtrl.scala 736:76]
  wire [1:0] _GEN_91629 = _GEN_90368 == _GEN_91578 ? _GEN_91589 : _GEN_91609; // @[FanCtrl.scala 736:76]
  wire [1:0] _GEN_91630 = _GEN_90368 == _GEN_91578 ? _GEN_91590 : _GEN_91610; // @[FanCtrl.scala 736:76]
  wire [1:0] _GEN_91631 = _GEN_90368 == _GEN_91578 ? _GEN_91591 : _GEN_91611; // @[FanCtrl.scala 736:76]
  wire [1:0] _GEN_91632 = _GEN_90368 == _GEN_91578 ? _GEN_91592 : _GEN_91612; // @[FanCtrl.scala 736:76]
  wire [1:0] _GEN_91633 = _GEN_90368 == _GEN_91578 ? _GEN_91593 : _GEN_91613; // @[FanCtrl.scala 736:76]
  wire [1:0] _GEN_91634 = _GEN_90368 == _GEN_91578 ? _GEN_91594 : _GEN_91614; // @[FanCtrl.scala 736:76]
  wire [1:0] _GEN_91635 = _GEN_90368 == _GEN_91578 ? _GEN_91595 : _GEN_91615; // @[FanCtrl.scala 736:76]
  wire [1:0] _GEN_91636 = _GEN_90368 == _GEN_91578 ? _GEN_91596 : _GEN_91616; // @[FanCtrl.scala 736:76]
  wire [1:0] _GEN_91637 = _GEN_90368 == _GEN_91578 ? _GEN_91597 : _GEN_91617; // @[FanCtrl.scala 736:76]
  wire [1:0] _GEN_91638 = _GEN_90368 == _GEN_91578 ? _GEN_91598 : _GEN_91618; // @[FanCtrl.scala 736:76]
  wire [1:0] _GEN_91639 = _GEN_90368 == _GEN_91494 ? _GEN_91495 : _GEN_91619; // @[FanCtrl.scala 734:76]
  wire [1:0] _GEN_91640 = _GEN_90368 == _GEN_91494 ? _GEN_91496 : _GEN_91620; // @[FanCtrl.scala 734:76]
  wire [1:0] _GEN_91641 = _GEN_90368 == _GEN_91494 ? _GEN_91497 : _GEN_91621; // @[FanCtrl.scala 734:76]
  wire [1:0] _GEN_91642 = _GEN_90368 == _GEN_91494 ? _GEN_91498 : _GEN_91622; // @[FanCtrl.scala 734:76]
  wire [1:0] _GEN_91643 = _GEN_90368 == _GEN_91494 ? _GEN_91499 : _GEN_91623; // @[FanCtrl.scala 734:76]
  wire [1:0] _GEN_91644 = _GEN_90368 == _GEN_91494 ? _GEN_91500 : _GEN_91624; // @[FanCtrl.scala 734:76]
  wire [1:0] _GEN_91645 = _GEN_90368 == _GEN_91494 ? _GEN_91501 : _GEN_91625; // @[FanCtrl.scala 734:76]
  wire [1:0] _GEN_91646 = _GEN_90368 == _GEN_91494 ? _GEN_91502 : _GEN_91626; // @[FanCtrl.scala 734:76]
  wire [1:0] _GEN_91647 = _GEN_90368 == _GEN_91494 ? _GEN_91503 : _GEN_91627; // @[FanCtrl.scala 734:76]
  wire [1:0] _GEN_91648 = _GEN_90368 == _GEN_91494 ? _GEN_91504 : _GEN_91628; // @[FanCtrl.scala 734:76]
  wire [1:0] _GEN_91649 = _GEN_90368 == _GEN_91494 ? _GEN_91505 : _GEN_91629; // @[FanCtrl.scala 734:76]
  wire [1:0] _GEN_91650 = _GEN_90368 == _GEN_91494 ? _GEN_91506 : _GEN_91630; // @[FanCtrl.scala 734:76]
  wire [1:0] _GEN_91651 = _GEN_90368 == _GEN_91494 ? _GEN_91507 : _GEN_91631; // @[FanCtrl.scala 734:76]
  wire [1:0] _GEN_91652 = _GEN_90368 == _GEN_91494 ? _GEN_91508 : _GEN_91632; // @[FanCtrl.scala 734:76]
  wire [1:0] _GEN_91653 = _GEN_90368 == _GEN_91494 ? _GEN_91509 : _GEN_91633; // @[FanCtrl.scala 734:76]
  wire [1:0] _GEN_91654 = _GEN_90368 == _GEN_91494 ? _GEN_91510 : _GEN_91634; // @[FanCtrl.scala 734:76]
  wire [1:0] _GEN_91655 = _GEN_90368 == _GEN_91494 ? _GEN_91511 : _GEN_91635; // @[FanCtrl.scala 734:76]
  wire [1:0] _GEN_91656 = _GEN_90368 == _GEN_91494 ? _GEN_91512 : _GEN_91636; // @[FanCtrl.scala 734:76]
  wire [1:0] _GEN_91657 = _GEN_90368 == _GEN_91494 ? _GEN_91513 : _GEN_91637; // @[FanCtrl.scala 734:76]
  wire [1:0] _GEN_91658 = _GEN_90368 == _GEN_91494 ? _GEN_91514 : _GEN_91638; // @[FanCtrl.scala 734:76]
  wire [1:0] _GEN_91659 = _GEN_90368 == _GEN_90525 ? _GEN_91411 : _GEN_91639; // @[FanCtrl.scala 732:69]
  wire [1:0] _GEN_91660 = _GEN_90368 == _GEN_90525 ? _GEN_91412 : _GEN_91640; // @[FanCtrl.scala 732:69]
  wire [1:0] _GEN_91661 = _GEN_90368 == _GEN_90525 ? _GEN_91413 : _GEN_91641; // @[FanCtrl.scala 732:69]
  wire [1:0] _GEN_91662 = _GEN_90368 == _GEN_90525 ? _GEN_91414 : _GEN_91642; // @[FanCtrl.scala 732:69]
  wire [1:0] _GEN_91663 = _GEN_90368 == _GEN_90525 ? _GEN_91415 : _GEN_91643; // @[FanCtrl.scala 732:69]
  wire [1:0] _GEN_91664 = _GEN_90368 == _GEN_90525 ? _GEN_91416 : _GEN_91644; // @[FanCtrl.scala 732:69]
  wire [1:0] _GEN_91665 = _GEN_90368 == _GEN_90525 ? _GEN_91417 : _GEN_91645; // @[FanCtrl.scala 732:69]
  wire [1:0] _GEN_91666 = _GEN_90368 == _GEN_90525 ? _GEN_91418 : _GEN_91646; // @[FanCtrl.scala 732:69]
  wire [1:0] _GEN_91667 = _GEN_90368 == _GEN_90525 ? _GEN_91419 : _GEN_91647; // @[FanCtrl.scala 732:69]
  wire [1:0] _GEN_91668 = _GEN_90368 == _GEN_90525 ? _GEN_91420 : _GEN_91648; // @[FanCtrl.scala 732:69]
  wire [1:0] _GEN_91669 = _GEN_90368 == _GEN_90525 ? _GEN_91421 : _GEN_91649; // @[FanCtrl.scala 732:69]
  wire [1:0] _GEN_91670 = _GEN_90368 == _GEN_90525 ? _GEN_91422 : _GEN_91650; // @[FanCtrl.scala 732:69]
  wire [1:0] _GEN_91671 = _GEN_90368 == _GEN_90525 ? _GEN_91423 : _GEN_91651; // @[FanCtrl.scala 732:69]
  wire [1:0] _GEN_91672 = _GEN_90368 == _GEN_90525 ? _GEN_91424 : _GEN_91652; // @[FanCtrl.scala 732:69]
  wire [1:0] _GEN_91673 = _GEN_90368 == _GEN_90525 ? _GEN_91425 : _GEN_91653; // @[FanCtrl.scala 732:69]
  wire [1:0] _GEN_91674 = _GEN_90368 == _GEN_90525 ? _GEN_91426 : _GEN_91654; // @[FanCtrl.scala 732:69]
  wire [1:0] _GEN_91675 = _GEN_90368 == _GEN_90525 ? _GEN_91427 : _GEN_91655; // @[FanCtrl.scala 732:69]
  wire [1:0] _GEN_91676 = _GEN_90368 == _GEN_90525 ? _GEN_91428 : _GEN_91656; // @[FanCtrl.scala 732:69]
  wire [1:0] _GEN_91677 = _GEN_90368 == _GEN_90525 ? _GEN_91429 : _GEN_91657; // @[FanCtrl.scala 732:69]
  wire [1:0] _GEN_91678 = _GEN_90368 == _GEN_90525 ? _GEN_91430 : _GEN_91658; // @[FanCtrl.scala 732:69]
  wire [1:0] _GEN_91699 = r_valid_1 ? _GEN_91659 : _GEN_91411; // @[FanCtrl.scala 731:33]
  wire [1:0] _GEN_91700 = r_valid_1 ? _GEN_91660 : _GEN_91412; // @[FanCtrl.scala 731:33]
  wire [1:0] _GEN_91701 = r_valid_1 ? _GEN_91661 : _GEN_91413; // @[FanCtrl.scala 731:33]
  wire [1:0] _GEN_91702 = r_valid_1 ? _GEN_91662 : _GEN_91414; // @[FanCtrl.scala 731:33]
  wire [1:0] _GEN_91703 = r_valid_1 ? _GEN_91663 : _GEN_91415; // @[FanCtrl.scala 731:33]
  wire [1:0] _GEN_91704 = r_valid_1 ? _GEN_91664 : _GEN_91416; // @[FanCtrl.scala 731:33]
  wire [1:0] _GEN_91705 = r_valid_1 ? _GEN_91665 : _GEN_91417; // @[FanCtrl.scala 731:33]
  wire [1:0] _GEN_91706 = r_valid_1 ? _GEN_91666 : _GEN_91418; // @[FanCtrl.scala 731:33]
  wire [1:0] _GEN_91707 = r_valid_1 ? _GEN_91667 : _GEN_91419; // @[FanCtrl.scala 731:33]
  wire [1:0] _GEN_91708 = r_valid_1 ? _GEN_91668 : _GEN_91420; // @[FanCtrl.scala 731:33]
  wire [1:0] _GEN_91709 = r_valid_1 ? _GEN_91669 : _GEN_91421; // @[FanCtrl.scala 731:33]
  wire [1:0] _GEN_91710 = r_valid_1 ? _GEN_91670 : _GEN_91422; // @[FanCtrl.scala 731:33]
  wire [1:0] _GEN_91711 = r_valid_1 ? _GEN_91671 : _GEN_91423; // @[FanCtrl.scala 731:33]
  wire [1:0] _GEN_91712 = r_valid_1 ? _GEN_91672 : _GEN_91424; // @[FanCtrl.scala 731:33]
  wire [1:0] _GEN_91713 = r_valid_1 ? _GEN_91673 : _GEN_91425; // @[FanCtrl.scala 731:33]
  wire [1:0] _GEN_91714 = r_valid_1 ? _GEN_91674 : _GEN_91426; // @[FanCtrl.scala 731:33]
  wire [1:0] _GEN_91715 = r_valid_1 ? _GEN_91675 : _GEN_91427; // @[FanCtrl.scala 731:33]
  wire [1:0] _GEN_91716 = r_valid_1 ? _GEN_91676 : _GEN_91428; // @[FanCtrl.scala 731:33]
  wire [1:0] _GEN_91717 = r_valid_1 ? _GEN_91677 : _GEN_91429; // @[FanCtrl.scala 731:33]
  wire [1:0] _GEN_91718 = r_valid_1 ? _GEN_91678 : _GEN_91430; // @[FanCtrl.scala 731:33]
  wire [4:0] _T_9154 = _GEN_98086 + 5'h12; // @[FanCtrl.scala 747:39]
  wire [6:0] _T_9161 = _T_8997 + 7'h14; // @[FanCtrl.scala 748:67]
  wire [4:0] _GEN_91838 = 5'h3 == _T_9161[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 748:{47,47}]
  wire [4:0] _GEN_91839 = 5'h4 == _T_9161[4:0] ? w_vn_4 : _GEN_91838; // @[FanCtrl.scala 748:{47,47}]
  wire [4:0] _GEN_91840 = 5'h5 == _T_9161[4:0] ? 5'h0 : _GEN_91839; // @[FanCtrl.scala 748:{47,47}]
  wire [4:0] _GEN_91841 = 5'h6 == _T_9161[4:0] ? 5'h0 : _GEN_91840; // @[FanCtrl.scala 748:{47,47}]
  wire [4:0] _GEN_91842 = 5'h7 == _T_9161[4:0] ? w_vn_7 : _GEN_91841; // @[FanCtrl.scala 748:{47,47}]
  wire [4:0] _GEN_91843 = 5'h8 == _T_9161[4:0] ? w_vn_8 : _GEN_91842; // @[FanCtrl.scala 748:{47,47}]
  wire [4:0] _GEN_91844 = 5'h9 == _T_9161[4:0] ? 5'h0 : _GEN_91843; // @[FanCtrl.scala 748:{47,47}]
  wire [4:0] _GEN_91845 = 5'ha == _T_9161[4:0] ? 5'h0 : _GEN_91844; // @[FanCtrl.scala 748:{47,47}]
  wire [4:0] _GEN_91846 = 5'hb == _T_9161[4:0] ? w_vn_11 : _GEN_91845; // @[FanCtrl.scala 748:{47,47}]
  wire [4:0] _GEN_91847 = 5'hc == _T_9161[4:0] ? w_vn_12 : _GEN_91846; // @[FanCtrl.scala 748:{47,47}]
  wire [4:0] _GEN_91848 = 5'hd == _T_9161[4:0] ? w_vn_13 : _GEN_91847; // @[FanCtrl.scala 748:{47,47}]
  wire [4:0] _GEN_91849 = 5'he == _T_9161[4:0] ? 5'h0 : _GEN_91848; // @[FanCtrl.scala 748:{47,47}]
  wire [4:0] _GEN_91850 = 5'hf == _T_9161[4:0] ? w_vn_15 : _GEN_91849; // @[FanCtrl.scala 748:{47,47}]
  wire [4:0] _GEN_91851 = 5'h10 == _T_9161[4:0] ? w_vn_16 : _GEN_91850; // @[FanCtrl.scala 748:{47,47}]
  wire [4:0] _GEN_91852 = 5'h11 == _T_9161[4:0] ? 5'h0 : _GEN_91851; // @[FanCtrl.scala 748:{47,47}]
  wire [4:0] _GEN_91853 = 5'h12 == _T_9161[4:0] ? w_vn_18 : _GEN_91852; // @[FanCtrl.scala 748:{47,47}]
  wire [4:0] _GEN_91854 = 5'h13 == _T_9161[4:0] ? 5'h0 : _GEN_91853; // @[FanCtrl.scala 748:{47,47}]
  wire [4:0] _GEN_91855 = 5'h14 == _T_9161[4:0] ? 5'h0 : _GEN_91854; // @[FanCtrl.scala 748:{47,47}]
  wire [4:0] _GEN_91856 = 5'h15 == _T_9161[4:0] ? 5'h0 : _GEN_91855; // @[FanCtrl.scala 748:{47,47}]
  wire [4:0] _GEN_91857 = 5'h16 == _T_9161[4:0] ? 5'h0 : _GEN_91856; // @[FanCtrl.scala 748:{47,47}]
  wire [4:0] _GEN_91858 = 5'h17 == _T_9161[4:0] ? w_vn_23 : _GEN_91857; // @[FanCtrl.scala 748:{47,47}]
  wire [4:0] _GEN_91859 = 5'h18 == _T_9161[4:0] ? w_vn_24 : _GEN_91858; // @[FanCtrl.scala 748:{47,47}]
  wire [4:0] _GEN_91860 = 5'h19 == _T_9161[4:0] ? 5'h0 : _GEN_91859; // @[FanCtrl.scala 748:{47,47}]
  wire [4:0] _GEN_91861 = 5'h1a == _T_9161[4:0] ? 5'h0 : _GEN_91860; // @[FanCtrl.scala 748:{47,47}]
  wire [4:0] _GEN_91862 = 5'h1b == _T_9161[4:0] ? 5'h0 : _GEN_91861; // @[FanCtrl.scala 748:{47,47}]
  wire [4:0] _GEN_91863 = 5'h1c == _T_9161[4:0] ? 5'h0 : _GEN_91862; // @[FanCtrl.scala 748:{47,47}]
  wire [4:0] _GEN_91864 = 5'h1d == _T_9161[4:0] ? 5'h0 : _GEN_91863; // @[FanCtrl.scala 748:{47,47}]
  wire [4:0] _GEN_91865 = 5'h1e == _T_9161[4:0] ? 5'h0 : _GEN_91864; // @[FanCtrl.scala 748:{47,47}]
  wire [4:0] _GEN_91866 = 5'h1f == _T_9161[4:0] ? 5'h0 : _GEN_91865; // @[FanCtrl.scala 748:{47,47}]
  wire [1:0] _GEN_91867 = 5'h0 == _T_9154 ? 2'h2 : _GEN_91699; // @[FanCtrl.scala 749:{47,47}]
  wire [1:0] _GEN_91868 = 5'h1 == _T_9154 ? 2'h2 : _GEN_91700; // @[FanCtrl.scala 749:{47,47}]
  wire [1:0] _GEN_91869 = 5'h2 == _T_9154 ? 2'h2 : _GEN_91701; // @[FanCtrl.scala 749:{47,47}]
  wire [1:0] _GEN_91870 = 5'h3 == _T_9154 ? 2'h2 : _GEN_91702; // @[FanCtrl.scala 749:{47,47}]
  wire [1:0] _GEN_91871 = 5'h4 == _T_9154 ? 2'h2 : _GEN_91703; // @[FanCtrl.scala 749:{47,47}]
  wire [1:0] _GEN_91872 = 5'h5 == _T_9154 ? 2'h2 : _GEN_91704; // @[FanCtrl.scala 749:{47,47}]
  wire [1:0] _GEN_91873 = 5'h6 == _T_9154 ? 2'h2 : _GEN_91705; // @[FanCtrl.scala 749:{47,47}]
  wire [1:0] _GEN_91874 = 5'h7 == _T_9154 ? 2'h2 : _GEN_91706; // @[FanCtrl.scala 749:{47,47}]
  wire [1:0] _GEN_91875 = 5'h8 == _T_9154 ? 2'h2 : _GEN_91707; // @[FanCtrl.scala 749:{47,47}]
  wire [1:0] _GEN_91876 = 5'h9 == _T_9154 ? 2'h2 : _GEN_91708; // @[FanCtrl.scala 749:{47,47}]
  wire [1:0] _GEN_91877 = 5'ha == _T_9154 ? 2'h2 : _GEN_91709; // @[FanCtrl.scala 749:{47,47}]
  wire [1:0] _GEN_91878 = 5'hb == _T_9154 ? 2'h2 : _GEN_91710; // @[FanCtrl.scala 749:{47,47}]
  wire [1:0] _GEN_91879 = 5'hc == _T_9154 ? 2'h2 : _GEN_91711; // @[FanCtrl.scala 749:{47,47}]
  wire [1:0] _GEN_91880 = 5'hd == _T_9154 ? 2'h2 : _GEN_91712; // @[FanCtrl.scala 749:{47,47}]
  wire [1:0] _GEN_91881 = 5'he == _T_9154 ? 2'h2 : _GEN_91713; // @[FanCtrl.scala 749:{47,47}]
  wire [1:0] _GEN_91882 = 5'hf == _T_9154 ? 2'h2 : _GEN_91714; // @[FanCtrl.scala 749:{47,47}]
  wire [1:0] _GEN_91883 = 5'h10 == _T_9154 ? 2'h2 : _GEN_91715; // @[FanCtrl.scala 749:{47,47}]
  wire [1:0] _GEN_91884 = 5'h11 == _T_9154 ? 2'h2 : _GEN_91716; // @[FanCtrl.scala 749:{47,47}]
  wire [1:0] _GEN_91885 = 5'h12 == _T_9154 ? 2'h2 : _GEN_91717; // @[FanCtrl.scala 749:{47,47}]
  wire [1:0] _GEN_91886 = 5'h13 == _T_9154 ? 2'h2 : _GEN_91718; // @[FanCtrl.scala 749:{47,47}]
  wire [6:0] _T_9173 = _T_8997 + 7'h12; // @[FanCtrl.scala 750:66]
  wire [4:0] _GEN_91922 = 5'h3 == _T_9173[4:0] ? w_vn_3 : 5'h0; // @[FanCtrl.scala 750:{46,46}]
  wire [4:0] _GEN_91923 = 5'h4 == _T_9173[4:0] ? w_vn_4 : _GEN_91922; // @[FanCtrl.scala 750:{46,46}]
  wire [4:0] _GEN_91924 = 5'h5 == _T_9173[4:0] ? 5'h0 : _GEN_91923; // @[FanCtrl.scala 750:{46,46}]
  wire [4:0] _GEN_91925 = 5'h6 == _T_9173[4:0] ? 5'h0 : _GEN_91924; // @[FanCtrl.scala 750:{46,46}]
  wire [4:0] _GEN_91926 = 5'h7 == _T_9173[4:0] ? w_vn_7 : _GEN_91925; // @[FanCtrl.scala 750:{46,46}]
  wire [4:0] _GEN_91927 = 5'h8 == _T_9173[4:0] ? w_vn_8 : _GEN_91926; // @[FanCtrl.scala 750:{46,46}]
  wire [4:0] _GEN_91928 = 5'h9 == _T_9173[4:0] ? 5'h0 : _GEN_91927; // @[FanCtrl.scala 750:{46,46}]
  wire [4:0] _GEN_91929 = 5'ha == _T_9173[4:0] ? 5'h0 : _GEN_91928; // @[FanCtrl.scala 750:{46,46}]
  wire [4:0] _GEN_91930 = 5'hb == _T_9173[4:0] ? w_vn_11 : _GEN_91929; // @[FanCtrl.scala 750:{46,46}]
  wire [4:0] _GEN_91931 = 5'hc == _T_9173[4:0] ? w_vn_12 : _GEN_91930; // @[FanCtrl.scala 750:{46,46}]
  wire [4:0] _GEN_91932 = 5'hd == _T_9173[4:0] ? w_vn_13 : _GEN_91931; // @[FanCtrl.scala 750:{46,46}]
  wire [4:0] _GEN_91933 = 5'he == _T_9173[4:0] ? 5'h0 : _GEN_91932; // @[FanCtrl.scala 750:{46,46}]
  wire [4:0] _GEN_91934 = 5'hf == _T_9173[4:0] ? w_vn_15 : _GEN_91933; // @[FanCtrl.scala 750:{46,46}]
  wire [4:0] _GEN_91935 = 5'h10 == _T_9173[4:0] ? w_vn_16 : _GEN_91934; // @[FanCtrl.scala 750:{46,46}]
  wire [4:0] _GEN_91936 = 5'h11 == _T_9173[4:0] ? 5'h0 : _GEN_91935; // @[FanCtrl.scala 750:{46,46}]
  wire [4:0] _GEN_91937 = 5'h12 == _T_9173[4:0] ? w_vn_18 : _GEN_91936; // @[FanCtrl.scala 750:{46,46}]
  wire [4:0] _GEN_91938 = 5'h13 == _T_9173[4:0] ? 5'h0 : _GEN_91937; // @[FanCtrl.scala 750:{46,46}]
  wire [4:0] _GEN_91939 = 5'h14 == _T_9173[4:0] ? 5'h0 : _GEN_91938; // @[FanCtrl.scala 750:{46,46}]
  wire [4:0] _GEN_91940 = 5'h15 == _T_9173[4:0] ? 5'h0 : _GEN_91939; // @[FanCtrl.scala 750:{46,46}]
  wire [4:0] _GEN_91941 = 5'h16 == _T_9173[4:0] ? 5'h0 : _GEN_91940; // @[FanCtrl.scala 750:{46,46}]
  wire [4:0] _GEN_91942 = 5'h17 == _T_9173[4:0] ? w_vn_23 : _GEN_91941; // @[FanCtrl.scala 750:{46,46}]
  wire [4:0] _GEN_91943 = 5'h18 == _T_9173[4:0] ? w_vn_24 : _GEN_91942; // @[FanCtrl.scala 750:{46,46}]
  wire [4:0] _GEN_91944 = 5'h19 == _T_9173[4:0] ? 5'h0 : _GEN_91943; // @[FanCtrl.scala 750:{46,46}]
  wire [4:0] _GEN_91945 = 5'h1a == _T_9173[4:0] ? 5'h0 : _GEN_91944; // @[FanCtrl.scala 750:{46,46}]
  wire [4:0] _GEN_91946 = 5'h1b == _T_9173[4:0] ? 5'h0 : _GEN_91945; // @[FanCtrl.scala 750:{46,46}]
  wire [4:0] _GEN_91947 = 5'h1c == _T_9173[4:0] ? 5'h0 : _GEN_91946; // @[FanCtrl.scala 750:{46,46}]
  wire [4:0] _GEN_91948 = 5'h1d == _T_9173[4:0] ? 5'h0 : _GEN_91947; // @[FanCtrl.scala 750:{46,46}]
  wire [4:0] _GEN_91949 = 5'h1e == _T_9173[4:0] ? 5'h0 : _GEN_91948; // @[FanCtrl.scala 750:{46,46}]
  wire [4:0] _GEN_91950 = 5'h1f == _T_9173[4:0] ? 5'h0 : _GEN_91949; // @[FanCtrl.scala 750:{46,46}]
  wire [1:0] _GEN_91951 = 5'h0 == _T_9154 ? 2'h1 : _GEN_91699; // @[FanCtrl.scala 751:{47,47}]
  wire [1:0] _GEN_91952 = 5'h1 == _T_9154 ? 2'h1 : _GEN_91700; // @[FanCtrl.scala 751:{47,47}]
  wire [1:0] _GEN_91953 = 5'h2 == _T_9154 ? 2'h1 : _GEN_91701; // @[FanCtrl.scala 751:{47,47}]
  wire [1:0] _GEN_91954 = 5'h3 == _T_9154 ? 2'h1 : _GEN_91702; // @[FanCtrl.scala 751:{47,47}]
  wire [1:0] _GEN_91955 = 5'h4 == _T_9154 ? 2'h1 : _GEN_91703; // @[FanCtrl.scala 751:{47,47}]
  wire [1:0] _GEN_91956 = 5'h5 == _T_9154 ? 2'h1 : _GEN_91704; // @[FanCtrl.scala 751:{47,47}]
  wire [1:0] _GEN_91957 = 5'h6 == _T_9154 ? 2'h1 : _GEN_91705; // @[FanCtrl.scala 751:{47,47}]
  wire [1:0] _GEN_91958 = 5'h7 == _T_9154 ? 2'h1 : _GEN_91706; // @[FanCtrl.scala 751:{47,47}]
  wire [1:0] _GEN_91959 = 5'h8 == _T_9154 ? 2'h1 : _GEN_91707; // @[FanCtrl.scala 751:{47,47}]
  wire [1:0] _GEN_91960 = 5'h9 == _T_9154 ? 2'h1 : _GEN_91708; // @[FanCtrl.scala 751:{47,47}]
  wire [1:0] _GEN_91961 = 5'ha == _T_9154 ? 2'h1 : _GEN_91709; // @[FanCtrl.scala 751:{47,47}]
  wire [1:0] _GEN_91962 = 5'hb == _T_9154 ? 2'h1 : _GEN_91710; // @[FanCtrl.scala 751:{47,47}]
  wire [1:0] _GEN_91963 = 5'hc == _T_9154 ? 2'h1 : _GEN_91711; // @[FanCtrl.scala 751:{47,47}]
  wire [1:0] _GEN_91964 = 5'hd == _T_9154 ? 2'h1 : _GEN_91712; // @[FanCtrl.scala 751:{47,47}]
  wire [1:0] _GEN_91965 = 5'he == _T_9154 ? 2'h1 : _GEN_91713; // @[FanCtrl.scala 751:{47,47}]
  wire [1:0] _GEN_91966 = 5'hf == _T_9154 ? 2'h1 : _GEN_91714; // @[FanCtrl.scala 751:{47,47}]
  wire [1:0] _GEN_91967 = 5'h10 == _T_9154 ? 2'h1 : _GEN_91715; // @[FanCtrl.scala 751:{47,47}]
  wire [1:0] _GEN_91968 = 5'h11 == _T_9154 ? 2'h1 : _GEN_91716; // @[FanCtrl.scala 751:{47,47}]
  wire [1:0] _GEN_91969 = 5'h12 == _T_9154 ? 2'h1 : _GEN_91717; // @[FanCtrl.scala 751:{47,47}]
  wire [1:0] _GEN_91970 = 5'h13 == _T_9154 ? 2'h1 : _GEN_91718; // @[FanCtrl.scala 751:{47,47}]
  wire [1:0] _GEN_91971 = 5'h0 == _T_9154 ? 2'h0 : _GEN_91699; // @[FanCtrl.scala 753:{46,46}]
  wire [1:0] _GEN_91972 = 5'h1 == _T_9154 ? 2'h0 : _GEN_91700; // @[FanCtrl.scala 753:{46,46}]
  wire [1:0] _GEN_91973 = 5'h2 == _T_9154 ? 2'h0 : _GEN_91701; // @[FanCtrl.scala 753:{46,46}]
  wire [1:0] _GEN_91974 = 5'h3 == _T_9154 ? 2'h0 : _GEN_91702; // @[FanCtrl.scala 753:{46,46}]
  wire [1:0] _GEN_91975 = 5'h4 == _T_9154 ? 2'h0 : _GEN_91703; // @[FanCtrl.scala 753:{46,46}]
  wire [1:0] _GEN_91976 = 5'h5 == _T_9154 ? 2'h0 : _GEN_91704; // @[FanCtrl.scala 753:{46,46}]
  wire [1:0] _GEN_91977 = 5'h6 == _T_9154 ? 2'h0 : _GEN_91705; // @[FanCtrl.scala 753:{46,46}]
  wire [1:0] _GEN_91978 = 5'h7 == _T_9154 ? 2'h0 : _GEN_91706; // @[FanCtrl.scala 753:{46,46}]
  wire [1:0] _GEN_91979 = 5'h8 == _T_9154 ? 2'h0 : _GEN_91707; // @[FanCtrl.scala 753:{46,46}]
  wire [1:0] _GEN_91980 = 5'h9 == _T_9154 ? 2'h0 : _GEN_91708; // @[FanCtrl.scala 753:{46,46}]
  wire [1:0] _GEN_91981 = 5'ha == _T_9154 ? 2'h0 : _GEN_91709; // @[FanCtrl.scala 753:{46,46}]
  wire [1:0] _GEN_91982 = 5'hb == _T_9154 ? 2'h0 : _GEN_91710; // @[FanCtrl.scala 753:{46,46}]
  wire [1:0] _GEN_91983 = 5'hc == _T_9154 ? 2'h0 : _GEN_91711; // @[FanCtrl.scala 753:{46,46}]
  wire [1:0] _GEN_91984 = 5'hd == _T_9154 ? 2'h0 : _GEN_91712; // @[FanCtrl.scala 753:{46,46}]
  wire [1:0] _GEN_91985 = 5'he == _T_9154 ? 2'h0 : _GEN_91713; // @[FanCtrl.scala 753:{46,46}]
  wire [1:0] _GEN_91986 = 5'hf == _T_9154 ? 2'h0 : _GEN_91714; // @[FanCtrl.scala 753:{46,46}]
  wire [1:0] _GEN_91987 = 5'h10 == _T_9154 ? 2'h0 : _GEN_91715; // @[FanCtrl.scala 753:{46,46}]
  wire [1:0] _GEN_91988 = 5'h11 == _T_9154 ? 2'h0 : _GEN_91716; // @[FanCtrl.scala 753:{46,46}]
  wire [1:0] _GEN_91989 = 5'h12 == _T_9154 ? 2'h0 : _GEN_91717; // @[FanCtrl.scala 753:{46,46}]
  wire [1:0] _GEN_91990 = 5'h13 == _T_9154 ? 2'h0 : _GEN_91718; // @[FanCtrl.scala 753:{46,46}]
  wire [1:0] _GEN_91991 = _GEN_90400 == _GEN_91950 ? _GEN_91951 : _GEN_91971; // @[FanCtrl.scala 750:76]
  wire [1:0] _GEN_91992 = _GEN_90400 == _GEN_91950 ? _GEN_91952 : _GEN_91972; // @[FanCtrl.scala 750:76]
  wire [1:0] _GEN_91993 = _GEN_90400 == _GEN_91950 ? _GEN_91953 : _GEN_91973; // @[FanCtrl.scala 750:76]
  wire [1:0] _GEN_91994 = _GEN_90400 == _GEN_91950 ? _GEN_91954 : _GEN_91974; // @[FanCtrl.scala 750:76]
  wire [1:0] _GEN_91995 = _GEN_90400 == _GEN_91950 ? _GEN_91955 : _GEN_91975; // @[FanCtrl.scala 750:76]
  wire [1:0] _GEN_91996 = _GEN_90400 == _GEN_91950 ? _GEN_91956 : _GEN_91976; // @[FanCtrl.scala 750:76]
  wire [1:0] _GEN_91997 = _GEN_90400 == _GEN_91950 ? _GEN_91957 : _GEN_91977; // @[FanCtrl.scala 750:76]
  wire [1:0] _GEN_91998 = _GEN_90400 == _GEN_91950 ? _GEN_91958 : _GEN_91978; // @[FanCtrl.scala 750:76]
  wire [1:0] _GEN_91999 = _GEN_90400 == _GEN_91950 ? _GEN_91959 : _GEN_91979; // @[FanCtrl.scala 750:76]
  wire [1:0] _GEN_92000 = _GEN_90400 == _GEN_91950 ? _GEN_91960 : _GEN_91980; // @[FanCtrl.scala 750:76]
  wire [1:0] _GEN_92001 = _GEN_90400 == _GEN_91950 ? _GEN_91961 : _GEN_91981; // @[FanCtrl.scala 750:76]
  wire [1:0] _GEN_92002 = _GEN_90400 == _GEN_91950 ? _GEN_91962 : _GEN_91982; // @[FanCtrl.scala 750:76]
  wire [1:0] _GEN_92003 = _GEN_90400 == _GEN_91950 ? _GEN_91963 : _GEN_91983; // @[FanCtrl.scala 750:76]
  wire [1:0] _GEN_92004 = _GEN_90400 == _GEN_91950 ? _GEN_91964 : _GEN_91984; // @[FanCtrl.scala 750:76]
  wire [1:0] _GEN_92005 = _GEN_90400 == _GEN_91950 ? _GEN_91965 : _GEN_91985; // @[FanCtrl.scala 750:76]
  wire [1:0] _GEN_92006 = _GEN_90400 == _GEN_91950 ? _GEN_91966 : _GEN_91986; // @[FanCtrl.scala 750:76]
  wire [1:0] _GEN_92007 = _GEN_90400 == _GEN_91950 ? _GEN_91967 : _GEN_91987; // @[FanCtrl.scala 750:76]
  wire [1:0] _GEN_92008 = _GEN_90400 == _GEN_91950 ? _GEN_91968 : _GEN_91988; // @[FanCtrl.scala 750:76]
  wire [1:0] _GEN_92009 = _GEN_90400 == _GEN_91950 ? _GEN_91969 : _GEN_91989; // @[FanCtrl.scala 750:76]
  wire [1:0] _GEN_92010 = _GEN_90400 == _GEN_91950 ? _GEN_91970 : _GEN_91990; // @[FanCtrl.scala 750:76]
  assign io_o_reduction_add_0 = r_add_lvl_4Reg_4; // @[FanCtrl.scala 1011:{35,35}]
  assign io_o_reduction_add_1 = r_add_lvl_3Reg_6; // @[FanCtrl.scala 1011:{35,35}]
  assign io_o_reduction_add_2 = r_add_lvl_3Reg_7; // @[FanCtrl.scala 1011:{35,35}]
  assign io_o_reduction_add_3 = r_add_lvl_2Reg_8; // @[FanCtrl.scala 1011:{35,35}]
  assign io_o_reduction_add_4 = r_add_lvl_2Reg_9; // @[FanCtrl.scala 1011:{35,35}]
  assign io_o_reduction_add_5 = r_add_lvl_2Reg_10; // @[FanCtrl.scala 1011:{35,35}]
  assign io_o_reduction_add_6 = r_add_lvl_2Reg_11; // @[FanCtrl.scala 1011:{35,35}]
  assign io_o_reduction_add_7 = r_add_lvl_1Reg_8; // @[FanCtrl.scala 1011:{35,35}]
  assign io_o_reduction_add_8 = r_add_lvl_1Reg_9; // @[FanCtrl.scala 1011:{35,35}]
  assign io_o_reduction_add_9 = r_add_lvl_1Reg_10; // @[FanCtrl.scala 1011:{35,35}]
  assign io_o_reduction_add_10 = r_add_lvl_1Reg_11; // @[FanCtrl.scala 1011:{35,35}]
  assign io_o_reduction_add_11 = r_add_lvl_1Reg_12; // @[FanCtrl.scala 1011:{35,35}]
  assign io_o_reduction_add_12 = r_add_lvl_1Reg_13; // @[FanCtrl.scala 1011:{35,35}]
  assign io_o_reduction_add_13 = r_add_lvl_1Reg_14; // @[FanCtrl.scala 1011:{35,35}]
  assign io_o_reduction_add_14 = r_add_lvl_1Reg_15; // @[FanCtrl.scala 1011:{35,35}]
  assign io_o_reduction_add_15 = r_add_lvl_0Reg_0; // @[FanCtrl.scala 1011:{35,35}]
  assign io_o_reduction_add_16 = r_add_lvl_0Reg_1; // @[FanCtrl.scala 1011:{35,35}]
  assign io_o_reduction_add_17 = r_add_lvl_0Reg_2; // @[FanCtrl.scala 1011:{35,35}]
  assign io_o_reduction_add_18 = r_add_lvl_0Reg_3; // @[FanCtrl.scala 1011:{35,35}]
  assign io_o_reduction_add_19 = r_add_lvl_0Reg_4; // @[FanCtrl.scala 1011:{35,35}]
  assign io_o_reduction_add_20 = r_add_lvl_0Reg_5; // @[FanCtrl.scala 1011:{35,35}]
  assign io_o_reduction_add_21 = r_add_lvl_0Reg_6; // @[FanCtrl.scala 1011:{35,35}]
  assign io_o_reduction_add_22 = r_add_lvl_0Reg_7; // @[FanCtrl.scala 1011:{35,35}]
  assign io_o_reduction_add_23 = r_add_lvl_0Reg_8; // @[FanCtrl.scala 1011:{35,35}]
  assign io_o_reduction_add_24 = r_add_lvl_0Reg_9; // @[FanCtrl.scala 1011:{35,35}]
  assign io_o_reduction_add_25 = r_add_lvl_0Reg_10; // @[FanCtrl.scala 1011:{35,35}]
  assign io_o_reduction_add_26 = r_add_lvl_0Reg_11; // @[FanCtrl.scala 1011:{35,35}]
  assign io_o_reduction_add_27 = r_add_lvl_0Reg_12; // @[FanCtrl.scala 1011:{35,35}]
  assign io_o_reduction_add_28 = r_add_lvl_0Reg_13; // @[FanCtrl.scala 1011:{35,35}]
  assign io_o_reduction_add_29 = r_add_lvl_0Reg_14; // @[FanCtrl.scala 1011:{35,35}]
  assign io_o_reduction_add_30 = r_add_lvl_0Reg_15; // @[FanCtrl.scala 1011:{35,35}]
  assign io_o_reduction_cmd_0 = r_cmd_lvl_4Reg_4; // @[FanCtrl.scala 1047:{34,34}]
  assign io_o_reduction_cmd_1 = r_cmd_lvl_3Reg_6; // @[FanCtrl.scala 1047:{34,34}]
  assign io_o_reduction_cmd_2 = r_cmd_lvl_3Reg_7; // @[FanCtrl.scala 1047:{34,34}]
  assign io_o_reduction_cmd_3 = r_cmd_lvl_2Reg_8; // @[FanCtrl.scala 1047:{34,34}]
  assign io_o_reduction_cmd_4 = r_cmd_lvl_2Reg_9; // @[FanCtrl.scala 1047:{34,34}]
  assign io_o_reduction_cmd_5 = r_cmd_lvl_2Reg_10; // @[FanCtrl.scala 1047:{34,34}]
  assign io_o_reduction_cmd_6 = r_cmd_lvl_2Reg_11; // @[FanCtrl.scala 1047:{34,34}]
  assign io_o_reduction_cmd_7 = r_cmd_lvl_1Reg_8; // @[FanCtrl.scala 1047:{34,34}]
  assign io_o_reduction_cmd_8 = r_cmd_lvl_1Reg_9; // @[FanCtrl.scala 1047:{34,34}]
  assign io_o_reduction_cmd_9 = r_cmd_lvl_1Reg_10; // @[FanCtrl.scala 1047:{34,34}]
  assign io_o_reduction_cmd_10 = r_cmd_lvl_1Reg_11; // @[FanCtrl.scala 1047:{34,34}]
  assign io_o_reduction_cmd_11 = r_cmd_lvl_1Reg_12; // @[FanCtrl.scala 1047:{34,34}]
  assign io_o_reduction_cmd_12 = r_cmd_lvl_1Reg_13; // @[FanCtrl.scala 1047:{34,34}]
  assign io_o_reduction_cmd_13 = r_cmd_lvl_1Reg_14; // @[FanCtrl.scala 1047:{34,34}]
  assign io_o_reduction_cmd_14 = r_cmd_lvl_1Reg_15; // @[FanCtrl.scala 1047:{34,34}]
  assign io_o_reduction_cmd_15 = r_cmd_lvl_0Reg_0; // @[FanCtrl.scala 1047:{34,34}]
  assign io_o_reduction_cmd_16 = r_cmd_lvl_0Reg_1; // @[FanCtrl.scala 1047:{34,34}]
  assign io_o_reduction_cmd_17 = r_cmd_lvl_0Reg_2; // @[FanCtrl.scala 1047:{34,34}]
  assign io_o_reduction_cmd_18 = r_cmd_lvl_0Reg_3; // @[FanCtrl.scala 1047:{34,34}]
  assign io_o_reduction_cmd_19 = r_cmd_lvl_0Reg_4; // @[FanCtrl.scala 1047:{34,34}]
  assign io_o_reduction_cmd_20 = r_cmd_lvl_0Reg_5; // @[FanCtrl.scala 1047:{34,34}]
  assign io_o_reduction_cmd_21 = r_cmd_lvl_0Reg_6; // @[FanCtrl.scala 1047:{34,34}]
  assign io_o_reduction_cmd_22 = r_cmd_lvl_0Reg_7; // @[FanCtrl.scala 1047:{34,34}]
  assign io_o_reduction_cmd_23 = r_cmd_lvl_0Reg_8; // @[FanCtrl.scala 1047:{34,34}]
  assign io_o_reduction_cmd_24 = r_cmd_lvl_0Reg_9; // @[FanCtrl.scala 1047:{34,34}]
  assign io_o_reduction_cmd_25 = r_cmd_lvl_0Reg_10; // @[FanCtrl.scala 1047:{34,34}]
  assign io_o_reduction_cmd_26 = r_cmd_lvl_0Reg_11; // @[FanCtrl.scala 1047:{34,34}]
  assign io_o_reduction_cmd_27 = r_cmd_lvl_0Reg_12; // @[FanCtrl.scala 1047:{34,34}]
  assign io_o_reduction_cmd_28 = r_cmd_lvl_0Reg_13; // @[FanCtrl.scala 1047:{34,34}]
  assign io_o_reduction_cmd_29 = r_cmd_lvl_0Reg_14; // @[FanCtrl.scala 1047:{34,34}]
  assign io_o_reduction_cmd_30 = r_cmd_lvl_0Reg_15; // @[FanCtrl.scala 1047:{34,34}]
  assign io_o_reduction_sel_0 = r_sel_lvl_4Reg_16; // @[FanCtrl.scala 1082:{34,34}]
  assign io_o_reduction_sel_1 = r_sel_lvl_4Reg_17; // @[FanCtrl.scala 1082:{34,34}]
  assign io_o_reduction_sel_2 = r_sel_lvl_4Reg_18; // @[FanCtrl.scala 1082:{34,34}]
  assign io_o_reduction_sel_3 = r_sel_lvl_4Reg_19; // @[FanCtrl.scala 1082:{34,34}]
  assign io_o_reduction_sel_4 = r_sel_lvl_3Reg_24; // @[FanCtrl.scala 1082:{34,34}]
  assign io_o_reduction_sel_5 = r_sel_lvl_3Reg_25; // @[FanCtrl.scala 1082:{34,34}]
  assign io_o_reduction_sel_6 = r_sel_lvl_3Reg_26; // @[FanCtrl.scala 1082:{34,34}]
  assign io_o_reduction_sel_7 = r_sel_lvl_3Reg_27; // @[FanCtrl.scala 1082:{34,34}]
  assign io_o_reduction_sel_8 = r_sel_lvl_3Reg_28; // @[FanCtrl.scala 1082:{34,34}]
  assign io_o_reduction_sel_9 = r_sel_lvl_3Reg_29; // @[FanCtrl.scala 1082:{34,34}]
  assign io_o_reduction_sel_10 = r_sel_lvl_3Reg_30; // @[FanCtrl.scala 1082:{34,34}]
  assign io_o_reduction_sel_11 = r_sel_lvl_3Reg_31; // @[FanCtrl.scala 1082:{34,34}]
  assign io_o_reduction_sel_12 = r_sel_lvl_2Reg_16; // @[FanCtrl.scala 1082:{34,34}]
  assign io_o_reduction_sel_13 = r_sel_lvl_2Reg_17; // @[FanCtrl.scala 1082:{34,34}]
  assign io_o_reduction_sel_14 = r_sel_lvl_2Reg_18; // @[FanCtrl.scala 1082:{34,34}]
  assign io_o_reduction_sel_15 = r_sel_lvl_2Reg_19; // @[FanCtrl.scala 1082:{34,34}]
  assign io_o_reduction_sel_16 = r_sel_lvl_2Reg_20; // @[FanCtrl.scala 1082:{34,34}]
  assign io_o_reduction_sel_17 = r_sel_lvl_2Reg_21; // @[FanCtrl.scala 1082:{34,34}]
  assign io_o_reduction_sel_18 = r_sel_lvl_2Reg_22; // @[FanCtrl.scala 1082:{34,34}]
  assign io_o_reduction_sel_19 = r_sel_lvl_2Reg_23; // @[FanCtrl.scala 1082:{34,34}]
  assign io_o_reduction_valid = r_valid_3; // @[FanCtrl.scala 1010:26]
  always @(posedge clock) begin
    if (reset) begin // @[FanCtrl.scala 19:34]
      r_reduction_add_0 <= 1'h0; // @[FanCtrl.scala 19:34]
    end else begin
      r_reduction_add_0 <= _GEN_446;
    end
    if (reset) begin // @[FanCtrl.scala 19:34]
      r_reduction_add_1 <= 1'h0; // @[FanCtrl.scala 19:34]
    end else begin
      r_reduction_add_1 <= _GEN_2328;
    end
    if (reset) begin // @[FanCtrl.scala 19:34]
      r_reduction_add_2 <= 1'h0; // @[FanCtrl.scala 19:34]
    end else begin
      r_reduction_add_2 <= _GEN_4211;
    end
    if (reset) begin // @[FanCtrl.scala 19:34]
      r_reduction_add_3 <= 1'h0; // @[FanCtrl.scala 19:34]
    end else begin
      r_reduction_add_3 <= _GEN_6094;
    end
    if (reset) begin // @[FanCtrl.scala 19:34]
      r_reduction_add_4 <= 1'h0; // @[FanCtrl.scala 19:34]
    end else begin
      r_reduction_add_4 <= _GEN_7977;
    end
    if (reset) begin // @[FanCtrl.scala 19:34]
      r_reduction_add_5 <= 1'h0; // @[FanCtrl.scala 19:34]
    end else begin
      r_reduction_add_5 <= _GEN_9860;
    end
    if (reset) begin // @[FanCtrl.scala 19:34]
      r_reduction_add_6 <= 1'h0; // @[FanCtrl.scala 19:34]
    end else begin
      r_reduction_add_6 <= _GEN_11743;
    end
    if (reset) begin // @[FanCtrl.scala 19:34]
      r_reduction_add_7 <= 1'h0; // @[FanCtrl.scala 19:34]
    end else begin
      r_reduction_add_7 <= _GEN_13626;
    end
    if (reset) begin // @[FanCtrl.scala 19:34]
      r_reduction_add_8 <= 1'h0; // @[FanCtrl.scala 19:34]
    end else begin
      r_reduction_add_8 <= _GEN_15509;
    end
    if (reset) begin // @[FanCtrl.scala 19:34]
      r_reduction_add_9 <= 1'h0; // @[FanCtrl.scala 19:34]
    end else begin
      r_reduction_add_9 <= _GEN_17392;
    end
    if (reset) begin // @[FanCtrl.scala 19:34]
      r_reduction_add_10 <= 1'h0; // @[FanCtrl.scala 19:34]
    end else begin
      r_reduction_add_10 <= _GEN_19275;
    end
    if (reset) begin // @[FanCtrl.scala 19:34]
      r_reduction_add_11 <= 1'h0; // @[FanCtrl.scala 19:34]
    end else begin
      r_reduction_add_11 <= _GEN_21158;
    end
    if (reset) begin // @[FanCtrl.scala 19:34]
      r_reduction_add_12 <= 1'h0; // @[FanCtrl.scala 19:34]
    end else begin
      r_reduction_add_12 <= _GEN_23041;
    end
    if (reset) begin // @[FanCtrl.scala 19:34]
      r_reduction_add_13 <= 1'h0; // @[FanCtrl.scala 19:34]
    end else begin
      r_reduction_add_13 <= _GEN_24924;
    end
    if (reset) begin // @[FanCtrl.scala 19:34]
      r_reduction_add_14 <= 1'h0; // @[FanCtrl.scala 19:34]
    end else begin
      r_reduction_add_14 <= _GEN_26807;
    end
    if (reset) begin // @[FanCtrl.scala 19:34]
      r_reduction_add_15 <= 1'h0; // @[FanCtrl.scala 19:34]
    end else begin
      r_reduction_add_15 <= _GEN_28690;
    end
    if (reset) begin // @[FanCtrl.scala 19:34]
      r_reduction_add_16 <= 1'h0; // @[FanCtrl.scala 19:34]
    end else begin
      r_reduction_add_16 <= _GEN_31201;
    end
    if (reset) begin // @[FanCtrl.scala 19:34]
      r_reduction_add_17 <= 1'h0; // @[FanCtrl.scala 19:34]
    end else begin
      r_reduction_add_17 <= _GEN_34862;
    end
    if (reset) begin // @[FanCtrl.scala 19:34]
      r_reduction_add_18 <= 1'h0; // @[FanCtrl.scala 19:34]
    end else begin
      r_reduction_add_18 <= _GEN_38523;
    end
    if (reset) begin // @[FanCtrl.scala 19:34]
      r_reduction_add_19 <= 1'h0; // @[FanCtrl.scala 19:34]
    end else begin
      r_reduction_add_19 <= _GEN_42184;
    end
    if (reset) begin // @[FanCtrl.scala 19:34]
      r_reduction_add_20 <= 1'h0; // @[FanCtrl.scala 19:34]
    end else begin
      r_reduction_add_20 <= _GEN_45845;
    end
    if (reset) begin // @[FanCtrl.scala 19:34]
      r_reduction_add_21 <= 1'h0; // @[FanCtrl.scala 19:34]
    end else begin
      r_reduction_add_21 <= _GEN_49506;
    end
    if (reset) begin // @[FanCtrl.scala 19:34]
      r_reduction_add_22 <= 1'h0; // @[FanCtrl.scala 19:34]
    end else begin
      r_reduction_add_22 <= _GEN_53167;
    end
    if (reset) begin // @[FanCtrl.scala 19:34]
      r_reduction_add_23 <= 1'h0; // @[FanCtrl.scala 19:34]
    end else begin
      r_reduction_add_23 <= _GEN_56828;
    end
    if (reset) begin // @[FanCtrl.scala 19:34]
      r_reduction_add_24 <= 1'h0; // @[FanCtrl.scala 19:34]
    end else begin
      r_reduction_add_24 <= _GEN_60573;
    end
    if (reset) begin // @[FanCtrl.scala 19:34]
      r_reduction_add_25 <= 1'h0; // @[FanCtrl.scala 19:34]
    end else begin
      r_reduction_add_25 <= _GEN_65510;
    end
    if (reset) begin // @[FanCtrl.scala 19:34]
      r_reduction_add_26 <= 1'h0; // @[FanCtrl.scala 19:34]
    end else begin
      r_reduction_add_26 <= _GEN_70447;
    end
    if (reset) begin // @[FanCtrl.scala 19:34]
      r_reduction_add_27 <= 1'h0; // @[FanCtrl.scala 19:34]
    end else begin
      r_reduction_add_27 <= _GEN_75384;
    end
    if (reset) begin // @[FanCtrl.scala 19:34]
      r_reduction_add_28 <= 1'h0; // @[FanCtrl.scala 19:34]
    end else begin
      r_reduction_add_28 <= _GEN_80321;
    end
    if (reset) begin // @[FanCtrl.scala 19:34]
      r_reduction_add_29 <= 1'h0; // @[FanCtrl.scala 19:34]
    end else begin
      r_reduction_add_29 <= _GEN_85882;
    end
    if (reset) begin // @[FanCtrl.scala 19:34]
      r_reduction_add_30 <= 1'h0; // @[FanCtrl.scala 19:34]
    end else begin
      r_reduction_add_30 <= _GEN_91315;
    end
    if (reset) begin // @[FanCtrl.scala 20:34]
      r_reduction_cmd_0 <= 3'h0; // @[FanCtrl.scala 20:34]
    end else if (r_valid_1) begin // @[FanCtrl.scala 340:33]
      if (_T_7505) begin // @[FanCtrl.scala 351:67]
        r_reduction_cmd_0 <= _GEN_477;
      end else if (_T_7536) begin // @[FanCtrl.scala 357:70]
        r_reduction_cmd_0 <= _GEN_477;
      end else begin
        r_reduction_cmd_0 <= _GEN_76750;
      end
    end else begin
      r_reduction_cmd_0 <= _GEN_477;
    end
    if (reset) begin // @[FanCtrl.scala 20:34]
      r_reduction_cmd_1 <= 3'h0; // @[FanCtrl.scala 20:34]
    end else if (r_valid_1) begin // @[FanCtrl.scala 340:33]
      if (_T_7505) begin // @[FanCtrl.scala 351:67]
        r_reduction_cmd_1 <= _GEN_3697;
      end else if (_T_7536) begin // @[FanCtrl.scala 357:70]
        r_reduction_cmd_1 <= _GEN_3697;
      end else begin
        r_reduction_cmd_1 <= _GEN_76751;
      end
    end else begin
      r_reduction_cmd_1 <= _GEN_3697;
    end
    if (reset) begin // @[FanCtrl.scala 20:34]
      r_reduction_cmd_2 <= 3'h0; // @[FanCtrl.scala 20:34]
    end else if (r_valid_1) begin // @[FanCtrl.scala 340:33]
      if (_T_7505) begin // @[FanCtrl.scala 351:67]
        r_reduction_cmd_2 <= _GEN_5579;
      end else if (_T_7536) begin // @[FanCtrl.scala 357:70]
        r_reduction_cmd_2 <= _GEN_5579;
      end else begin
        r_reduction_cmd_2 <= _GEN_76752;
      end
    end else begin
      r_reduction_cmd_2 <= _GEN_5579;
    end
    if (reset) begin // @[FanCtrl.scala 20:34]
      r_reduction_cmd_3 <= 3'h0; // @[FanCtrl.scala 20:34]
    end else if (r_valid_1) begin // @[FanCtrl.scala 340:33]
      if (_T_7505) begin // @[FanCtrl.scala 351:67]
        r_reduction_cmd_3 <= _GEN_7461;
      end else if (_T_7536) begin // @[FanCtrl.scala 357:70]
        r_reduction_cmd_3 <= _GEN_7461;
      end else begin
        r_reduction_cmd_3 <= _GEN_76753;
      end
    end else begin
      r_reduction_cmd_3 <= _GEN_7461;
    end
    if (reset) begin // @[FanCtrl.scala 20:34]
      r_reduction_cmd_4 <= 3'h0; // @[FanCtrl.scala 20:34]
    end else if (r_valid_1) begin // @[FanCtrl.scala 340:33]
      if (_T_7505) begin // @[FanCtrl.scala 351:67]
        r_reduction_cmd_4 <= _GEN_9343;
      end else if (_T_7536) begin // @[FanCtrl.scala 357:70]
        r_reduction_cmd_4 <= _GEN_9343;
      end else begin
        r_reduction_cmd_4 <= _GEN_76754;
      end
    end else begin
      r_reduction_cmd_4 <= _GEN_9343;
    end
    if (reset) begin // @[FanCtrl.scala 20:34]
      r_reduction_cmd_5 <= 3'h0; // @[FanCtrl.scala 20:34]
    end else if (r_valid_1) begin // @[FanCtrl.scala 340:33]
      if (_T_7505) begin // @[FanCtrl.scala 351:67]
        r_reduction_cmd_5 <= _GEN_11225;
      end else if (_T_7536) begin // @[FanCtrl.scala 357:70]
        r_reduction_cmd_5 <= _GEN_11225;
      end else begin
        r_reduction_cmd_5 <= _GEN_76755;
      end
    end else begin
      r_reduction_cmd_5 <= _GEN_11225;
    end
    if (reset) begin // @[FanCtrl.scala 20:34]
      r_reduction_cmd_6 <= 3'h0; // @[FanCtrl.scala 20:34]
    end else if (r_valid_1) begin // @[FanCtrl.scala 340:33]
      if (_T_7505) begin // @[FanCtrl.scala 351:67]
        r_reduction_cmd_6 <= _GEN_13107;
      end else if (_T_7536) begin // @[FanCtrl.scala 357:70]
        r_reduction_cmd_6 <= _GEN_13107;
      end else begin
        r_reduction_cmd_6 <= _GEN_76756;
      end
    end else begin
      r_reduction_cmd_6 <= _GEN_13107;
    end
    if (reset) begin // @[FanCtrl.scala 20:34]
      r_reduction_cmd_7 <= 3'h0; // @[FanCtrl.scala 20:34]
    end else if (r_valid_1) begin // @[FanCtrl.scala 340:33]
      if (_T_7505) begin // @[FanCtrl.scala 351:67]
        r_reduction_cmd_7 <= _GEN_14989;
      end else if (_T_7536) begin // @[FanCtrl.scala 357:70]
        r_reduction_cmd_7 <= _GEN_14989;
      end else begin
        r_reduction_cmd_7 <= _GEN_76757;
      end
    end else begin
      r_reduction_cmd_7 <= _GEN_14989;
    end
    if (reset) begin // @[FanCtrl.scala 20:34]
      r_reduction_cmd_8 <= 3'h0; // @[FanCtrl.scala 20:34]
    end else if (r_valid_1) begin // @[FanCtrl.scala 340:33]
      if (_T_7505) begin // @[FanCtrl.scala 351:67]
        r_reduction_cmd_8 <= _GEN_16871;
      end else if (_T_7536) begin // @[FanCtrl.scala 357:70]
        r_reduction_cmd_8 <= _GEN_16871;
      end else begin
        r_reduction_cmd_8 <= _GEN_76758;
      end
    end else begin
      r_reduction_cmd_8 <= _GEN_16871;
    end
    if (reset) begin // @[FanCtrl.scala 20:34]
      r_reduction_cmd_9 <= 3'h0; // @[FanCtrl.scala 20:34]
    end else if (r_valid_1) begin // @[FanCtrl.scala 340:33]
      if (_T_7505) begin // @[FanCtrl.scala 351:67]
        r_reduction_cmd_9 <= _GEN_18753;
      end else if (_T_7536) begin // @[FanCtrl.scala 357:70]
        r_reduction_cmd_9 <= _GEN_18753;
      end else begin
        r_reduction_cmd_9 <= _GEN_76759;
      end
    end else begin
      r_reduction_cmd_9 <= _GEN_18753;
    end
    if (reset) begin // @[FanCtrl.scala 20:34]
      r_reduction_cmd_10 <= 3'h0; // @[FanCtrl.scala 20:34]
    end else if (r_valid_1) begin // @[FanCtrl.scala 340:33]
      if (_T_7505) begin // @[FanCtrl.scala 351:67]
        r_reduction_cmd_10 <= _GEN_20635;
      end else if (_T_7536) begin // @[FanCtrl.scala 357:70]
        r_reduction_cmd_10 <= _GEN_20635;
      end else begin
        r_reduction_cmd_10 <= _GEN_76760;
      end
    end else begin
      r_reduction_cmd_10 <= _GEN_20635;
    end
    if (reset) begin // @[FanCtrl.scala 20:34]
      r_reduction_cmd_11 <= 3'h0; // @[FanCtrl.scala 20:34]
    end else if (r_valid_1) begin // @[FanCtrl.scala 340:33]
      if (_T_7505) begin // @[FanCtrl.scala 351:67]
        r_reduction_cmd_11 <= _GEN_22517;
      end else if (_T_7536) begin // @[FanCtrl.scala 357:70]
        r_reduction_cmd_11 <= _GEN_22517;
      end else begin
        r_reduction_cmd_11 <= _GEN_76761;
      end
    end else begin
      r_reduction_cmd_11 <= _GEN_22517;
    end
    if (reset) begin // @[FanCtrl.scala 20:34]
      r_reduction_cmd_12 <= 3'h0; // @[FanCtrl.scala 20:34]
    end else if (r_valid_1) begin // @[FanCtrl.scala 340:33]
      if (_T_7505) begin // @[FanCtrl.scala 351:67]
        r_reduction_cmd_12 <= _GEN_24399;
      end else if (_T_7536) begin // @[FanCtrl.scala 357:70]
        r_reduction_cmd_12 <= _GEN_24399;
      end else begin
        r_reduction_cmd_12 <= _GEN_76762;
      end
    end else begin
      r_reduction_cmd_12 <= _GEN_24399;
    end
    if (reset) begin // @[FanCtrl.scala 20:34]
      r_reduction_cmd_13 <= 3'h0; // @[FanCtrl.scala 20:34]
    end else if (r_valid_1) begin // @[FanCtrl.scala 340:33]
      if (_T_7505) begin // @[FanCtrl.scala 351:67]
        r_reduction_cmd_13 <= _GEN_26281;
      end else if (_T_7536) begin // @[FanCtrl.scala 357:70]
        r_reduction_cmd_13 <= _GEN_26281;
      end else begin
        r_reduction_cmd_13 <= _GEN_76763;
      end
    end else begin
      r_reduction_cmd_13 <= _GEN_26281;
    end
    if (reset) begin // @[FanCtrl.scala 20:34]
      r_reduction_cmd_14 <= 3'h0; // @[FanCtrl.scala 20:34]
    end else if (r_valid_1) begin // @[FanCtrl.scala 340:33]
      if (_T_7505) begin // @[FanCtrl.scala 351:67]
        r_reduction_cmd_14 <= _GEN_28163;
      end else if (_T_7536) begin // @[FanCtrl.scala 357:70]
        r_reduction_cmd_14 <= _GEN_28163;
      end else begin
        r_reduction_cmd_14 <= _GEN_76764;
      end
    end else begin
      r_reduction_cmd_14 <= _GEN_28163;
    end
    if (reset) begin // @[FanCtrl.scala 20:34]
      r_reduction_cmd_15 <= 3'h0; // @[FanCtrl.scala 20:34]
    end else if (r_valid_1) begin // @[FanCtrl.scala 340:33]
      if (_T_7505) begin // @[FanCtrl.scala 351:67]
        r_reduction_cmd_15 <= _GEN_29215;
      end else if (_T_7536) begin // @[FanCtrl.scala 357:70]
        r_reduction_cmd_15 <= _GEN_29215;
      end else begin
        r_reduction_cmd_15 <= _GEN_76765;
      end
    end else begin
      r_reduction_cmd_15 <= _GEN_29215;
    end
    if (reset) begin // @[FanCtrl.scala 20:34]
      r_reduction_cmd_16 <= 3'h0; // @[FanCtrl.scala 20:34]
    end else if (r_valid_1) begin // @[FanCtrl.scala 340:33]
      if (_T_7505) begin // @[FanCtrl.scala 351:67]
        r_reduction_cmd_16 <= _GEN_31232;
      end else if (_T_7536) begin // @[FanCtrl.scala 357:70]
        r_reduction_cmd_16 <= _GEN_31232;
      end else begin
        r_reduction_cmd_16 <= _GEN_76766;
      end
    end else begin
      r_reduction_cmd_16 <= _GEN_31232;
    end
    if (reset) begin // @[FanCtrl.scala 20:34]
      r_reduction_cmd_17 <= 3'h0; // @[FanCtrl.scala 20:34]
    end else if (r_valid_1) begin // @[FanCtrl.scala 340:33]
      if (_T_7505) begin // @[FanCtrl.scala 351:67]
        r_reduction_cmd_17 <= _GEN_37293;
      end else if (_T_7536) begin // @[FanCtrl.scala 357:70]
        r_reduction_cmd_17 <= _GEN_37293;
      end else begin
        r_reduction_cmd_17 <= _GEN_76767;
      end
    end else begin
      r_reduction_cmd_17 <= _GEN_37293;
    end
    if (reset) begin // @[FanCtrl.scala 20:34]
      r_reduction_cmd_18 <= 3'h0; // @[FanCtrl.scala 20:34]
    end else if (r_valid_1) begin // @[FanCtrl.scala 340:33]
      if (_T_7505) begin // @[FanCtrl.scala 351:67]
        r_reduction_cmd_18 <= _GEN_40954;
      end else if (_T_7536) begin // @[FanCtrl.scala 357:70]
        r_reduction_cmd_18 <= _GEN_40954;
      end else begin
        r_reduction_cmd_18 <= _GEN_76768;
      end
    end else begin
      r_reduction_cmd_18 <= _GEN_40954;
    end
    if (reset) begin // @[FanCtrl.scala 20:34]
      r_reduction_cmd_19 <= 3'h0; // @[FanCtrl.scala 20:34]
    end else if (r_valid_1) begin // @[FanCtrl.scala 340:33]
      if (_T_7505) begin // @[FanCtrl.scala 351:67]
        r_reduction_cmd_19 <= _GEN_44615;
      end else if (_T_7536) begin // @[FanCtrl.scala 357:70]
        r_reduction_cmd_19 <= _GEN_44615;
      end else begin
        r_reduction_cmd_19 <= _GEN_76769;
      end
    end else begin
      r_reduction_cmd_19 <= _GEN_44615;
    end
    if (reset) begin // @[FanCtrl.scala 20:34]
      r_reduction_cmd_20 <= 3'h0; // @[FanCtrl.scala 20:34]
    end else if (r_valid_1) begin // @[FanCtrl.scala 340:33]
      if (_T_7505) begin // @[FanCtrl.scala 351:67]
        r_reduction_cmd_20 <= _GEN_48276;
      end else if (_T_7536) begin // @[FanCtrl.scala 357:70]
        r_reduction_cmd_20 <= _GEN_48276;
      end else begin
        r_reduction_cmd_20 <= _GEN_76770;
      end
    end else begin
      r_reduction_cmd_20 <= _GEN_48276;
    end
    if (reset) begin // @[FanCtrl.scala 20:34]
      r_reduction_cmd_21 <= 3'h0; // @[FanCtrl.scala 20:34]
    end else if (r_valid_1) begin // @[FanCtrl.scala 340:33]
      if (_T_7505) begin // @[FanCtrl.scala 351:67]
        r_reduction_cmd_21 <= _GEN_51937;
      end else if (_T_7536) begin // @[FanCtrl.scala 357:70]
        r_reduction_cmd_21 <= _GEN_51937;
      end else begin
        r_reduction_cmd_21 <= _GEN_76771;
      end
    end else begin
      r_reduction_cmd_21 <= _GEN_51937;
    end
    if (reset) begin // @[FanCtrl.scala 20:34]
      r_reduction_cmd_22 <= 3'h0; // @[FanCtrl.scala 20:34]
    end else if (r_valid_1) begin // @[FanCtrl.scala 340:33]
      if (_T_7505) begin // @[FanCtrl.scala 351:67]
        r_reduction_cmd_22 <= _GEN_55598;
      end else if (_T_7536) begin // @[FanCtrl.scala 357:70]
        r_reduction_cmd_22 <= _GEN_55598;
      end else begin
        r_reduction_cmd_22 <= _GEN_76772;
      end
    end else begin
      r_reduction_cmd_22 <= _GEN_55598;
    end
    if (reset) begin // @[FanCtrl.scala 20:34]
      r_reduction_cmd_23 <= 3'h0; // @[FanCtrl.scala 20:34]
    end else if (r_valid_1) begin // @[FanCtrl.scala 340:33]
      if (_T_7505) begin // @[FanCtrl.scala 351:67]
        r_reduction_cmd_23 <= _GEN_57995;
      end else if (_T_7536) begin // @[FanCtrl.scala 357:70]
        r_reduction_cmd_23 <= _GEN_57995;
      end else begin
        r_reduction_cmd_23 <= _GEN_76773;
      end
    end else begin
      r_reduction_cmd_23 <= _GEN_57995;
    end
    if (reset) begin // @[FanCtrl.scala 20:34]
      r_reduction_cmd_24 <= 3'h0; // @[FanCtrl.scala 20:34]
    end else if (r_valid_1) begin // @[FanCtrl.scala 340:33]
      if (_T_7505) begin // @[FanCtrl.scala 351:67]
        r_reduction_cmd_24 <= _GEN_60604;
      end else if (_T_7536) begin // @[FanCtrl.scala 357:70]
        r_reduction_cmd_24 <= _GEN_60604;
      end else begin
        r_reduction_cmd_24 <= _GEN_76774;
      end
    end else begin
      r_reduction_cmd_24 <= _GEN_60604;
    end
    if (reset) begin // @[FanCtrl.scala 20:34]
      r_reduction_cmd_25 <= 3'h0; // @[FanCtrl.scala 20:34]
    end else if (r_valid_1) begin // @[FanCtrl.scala 340:33]
      if (_T_7505) begin // @[FanCtrl.scala 351:67]
        r_reduction_cmd_25 <= _GEN_68765;
      end else if (_T_7536) begin // @[FanCtrl.scala 357:70]
        r_reduction_cmd_25 <= _GEN_68765;
      end else begin
        r_reduction_cmd_25 <= _GEN_76775;
      end
    end else begin
      r_reduction_cmd_25 <= _GEN_68765;
    end
    if (reset) begin // @[FanCtrl.scala 20:34]
      r_reduction_cmd_26 <= 3'h0; // @[FanCtrl.scala 20:34]
    end else if (r_valid_1) begin // @[FanCtrl.scala 340:33]
      if (_T_7505) begin // @[FanCtrl.scala 351:67]
        r_reduction_cmd_26 <= _GEN_73702;
      end else if (_T_7536) begin // @[FanCtrl.scala 357:70]
        r_reduction_cmd_26 <= _GEN_73702;
      end else begin
        r_reduction_cmd_26 <= _GEN_76776;
      end
    end else begin
      r_reduction_cmd_26 <= _GEN_73702;
    end
    if (reset) begin // @[FanCtrl.scala 20:34]
      r_reduction_cmd_27 <= 3'h0; // @[FanCtrl.scala 20:34]
    end else if (r_valid_1) begin // @[FanCtrl.scala 340:33]
      if (_T_7505) begin // @[FanCtrl.scala 351:67]
        r_reduction_cmd_27 <= 3'h5;
      end else if (_T_7536) begin // @[FanCtrl.scala 357:70]
        r_reduction_cmd_27 <= 3'h3;
      end else begin
        r_reduction_cmd_27 <= _GEN_76777;
      end
    end else begin
      r_reduction_cmd_27 <= 3'h0;
    end
    if (reset) begin // @[FanCtrl.scala 20:34]
      r_reduction_cmd_28 <= 3'h0; // @[FanCtrl.scala 20:34]
    end else if (r_valid_1) begin // @[FanCtrl.scala 482:33]
      if (_T_7862) begin // @[FanCtrl.scala 493:70]
        r_reduction_cmd_28 <= 3'h5;
      end else if (_T_7893) begin // @[FanCtrl.scala 499:74]
        r_reduction_cmd_28 <= 3'h4;
      end else begin
        r_reduction_cmd_28 <= _GEN_80166;
      end
    end else begin
      r_reduction_cmd_28 <= 3'h0;
    end
    if (reset) begin // @[FanCtrl.scala 20:34]
      r_reduction_cmd_29 <= 3'h0; // @[FanCtrl.scala 20:34]
    end else if (r_valid_1) begin // @[FanCtrl.scala 558:33]
      if (_T_8653) begin // @[FanCtrl.scala 569:73]
        r_reduction_cmd_29 <= 3'h5;
      end else if (_T_8684) begin // @[FanCtrl.scala 575:77]
        r_reduction_cmd_29 <= 3'h3;
      end else begin
        r_reduction_cmd_29 <= _GEN_87483;
      end
    end else begin
      r_reduction_cmd_29 <= 3'h0;
    end
    if (reset) begin // @[FanCtrl.scala 20:34]
      r_reduction_cmd_30 <= 3'h0; // @[FanCtrl.scala 20:34]
    end else if (r_valid_1) begin // @[FanCtrl.scala 699:36]
      if (_T_9048) begin // @[FanCtrl.scala 709:71]
        r_reduction_cmd_30 <= 3'h5;
      end else if (_T_9069) begin // @[FanCtrl.scala 714:76]
        r_reduction_cmd_30 <= 3'h4;
      end else begin
        r_reduction_cmd_30 <= _GEN_91160;
      end
    end else begin
      r_reduction_cmd_30 <= 3'h0;
    end
    if (reset) begin // @[FanCtrl.scala 21:34]
      r_reduction_sel_0 <= 2'h0; // @[FanCtrl.scala 21:34]
    end else if (r_valid_1) begin // @[FanCtrl.scala 745:33]
      if (_GEN_90400 == _GEN_90621) begin // @[FanCtrl.scala 746:70]
        if (5'h0 == _T_9154) begin // @[FanCtrl.scala 747:46]
          r_reduction_sel_0 <= 2'h3; // @[FanCtrl.scala 747:46]
        end else begin
          r_reduction_sel_0 <= _GEN_91699;
        end
      end else if (_GEN_90400 == _GEN_91866) begin // @[FanCtrl.scala 748:77]
        r_reduction_sel_0 <= _GEN_91867;
      end else begin
        r_reduction_sel_0 <= _GEN_91991;
      end
    end else if (5'h0 == _T_9154) begin // @[FanCtrl.scala 753:46]
      r_reduction_sel_0 <= 2'h0; // @[FanCtrl.scala 753:46]
    end else begin
      r_reduction_sel_0 <= _GEN_91699;
    end
    if (reset) begin // @[FanCtrl.scala 21:34]
      r_reduction_sel_1 <= 2'h0; // @[FanCtrl.scala 21:34]
    end else if (r_valid_1) begin // @[FanCtrl.scala 745:33]
      if (_GEN_90400 == _GEN_90621) begin // @[FanCtrl.scala 746:70]
        if (5'h1 == _T_9154) begin // @[FanCtrl.scala 747:46]
          r_reduction_sel_1 <= 2'h3; // @[FanCtrl.scala 747:46]
        end else begin
          r_reduction_sel_1 <= _GEN_91700;
        end
      end else if (_GEN_90400 == _GEN_91866) begin // @[FanCtrl.scala 748:77]
        r_reduction_sel_1 <= _GEN_91868;
      end else begin
        r_reduction_sel_1 <= _GEN_91992;
      end
    end else if (5'h1 == _T_9154) begin // @[FanCtrl.scala 753:46]
      r_reduction_sel_1 <= 2'h0; // @[FanCtrl.scala 753:46]
    end else begin
      r_reduction_sel_1 <= _GEN_91700;
    end
    if (reset) begin // @[FanCtrl.scala 21:34]
      r_reduction_sel_2 <= 2'h0; // @[FanCtrl.scala 21:34]
    end else if (r_valid_1) begin // @[FanCtrl.scala 745:33]
      if (_GEN_90400 == _GEN_90621) begin // @[FanCtrl.scala 746:70]
        if (5'h2 == _T_9154) begin // @[FanCtrl.scala 747:46]
          r_reduction_sel_2 <= 2'h3; // @[FanCtrl.scala 747:46]
        end else begin
          r_reduction_sel_2 <= _GEN_91701;
        end
      end else if (_GEN_90400 == _GEN_91866) begin // @[FanCtrl.scala 748:77]
        r_reduction_sel_2 <= _GEN_91869;
      end else begin
        r_reduction_sel_2 <= _GEN_91993;
      end
    end else if (5'h2 == _T_9154) begin // @[FanCtrl.scala 753:46]
      r_reduction_sel_2 <= 2'h0; // @[FanCtrl.scala 753:46]
    end else begin
      r_reduction_sel_2 <= _GEN_91701;
    end
    if (reset) begin // @[FanCtrl.scala 21:34]
      r_reduction_sel_3 <= 2'h0; // @[FanCtrl.scala 21:34]
    end else if (r_valid_1) begin // @[FanCtrl.scala 745:33]
      if (_GEN_90400 == _GEN_90621) begin // @[FanCtrl.scala 746:70]
        if (5'h3 == _T_9154) begin // @[FanCtrl.scala 747:46]
          r_reduction_sel_3 <= 2'h3; // @[FanCtrl.scala 747:46]
        end else begin
          r_reduction_sel_3 <= _GEN_91702;
        end
      end else if (_GEN_90400 == _GEN_91866) begin // @[FanCtrl.scala 748:77]
        r_reduction_sel_3 <= _GEN_91870;
      end else begin
        r_reduction_sel_3 <= _GEN_91994;
      end
    end else if (5'h3 == _T_9154) begin // @[FanCtrl.scala 753:46]
      r_reduction_sel_3 <= 2'h0; // @[FanCtrl.scala 753:46]
    end else begin
      r_reduction_sel_3 <= _GEN_91702;
    end
    if (reset) begin // @[FanCtrl.scala 21:34]
      r_reduction_sel_4 <= 2'h0; // @[FanCtrl.scala 21:34]
    end else if (r_valid_1) begin // @[FanCtrl.scala 745:33]
      if (_GEN_90400 == _GEN_90621) begin // @[FanCtrl.scala 746:70]
        if (5'h4 == _T_9154) begin // @[FanCtrl.scala 747:46]
          r_reduction_sel_4 <= 2'h3; // @[FanCtrl.scala 747:46]
        end else begin
          r_reduction_sel_4 <= _GEN_91703;
        end
      end else if (_GEN_90400 == _GEN_91866) begin // @[FanCtrl.scala 748:77]
        r_reduction_sel_4 <= _GEN_91871;
      end else begin
        r_reduction_sel_4 <= _GEN_91995;
      end
    end else if (5'h4 == _T_9154) begin // @[FanCtrl.scala 753:46]
      r_reduction_sel_4 <= 2'h0; // @[FanCtrl.scala 753:46]
    end else begin
      r_reduction_sel_4 <= _GEN_91703;
    end
    if (reset) begin // @[FanCtrl.scala 21:34]
      r_reduction_sel_5 <= 2'h0; // @[FanCtrl.scala 21:34]
    end else if (r_valid_1) begin // @[FanCtrl.scala 745:33]
      if (_GEN_90400 == _GEN_90621) begin // @[FanCtrl.scala 746:70]
        if (5'h5 == _T_9154) begin // @[FanCtrl.scala 747:46]
          r_reduction_sel_5 <= 2'h3; // @[FanCtrl.scala 747:46]
        end else begin
          r_reduction_sel_5 <= _GEN_91704;
        end
      end else if (_GEN_90400 == _GEN_91866) begin // @[FanCtrl.scala 748:77]
        r_reduction_sel_5 <= _GEN_91872;
      end else begin
        r_reduction_sel_5 <= _GEN_91996;
      end
    end else if (5'h5 == _T_9154) begin // @[FanCtrl.scala 753:46]
      r_reduction_sel_5 <= 2'h0; // @[FanCtrl.scala 753:46]
    end else begin
      r_reduction_sel_5 <= _GEN_91704;
    end
    if (reset) begin // @[FanCtrl.scala 21:34]
      r_reduction_sel_6 <= 2'h0; // @[FanCtrl.scala 21:34]
    end else if (r_valid_1) begin // @[FanCtrl.scala 745:33]
      if (_GEN_90400 == _GEN_90621) begin // @[FanCtrl.scala 746:70]
        if (5'h6 == _T_9154) begin // @[FanCtrl.scala 747:46]
          r_reduction_sel_6 <= 2'h3; // @[FanCtrl.scala 747:46]
        end else begin
          r_reduction_sel_6 <= _GEN_91705;
        end
      end else if (_GEN_90400 == _GEN_91866) begin // @[FanCtrl.scala 748:77]
        r_reduction_sel_6 <= _GEN_91873;
      end else begin
        r_reduction_sel_6 <= _GEN_91997;
      end
    end else if (5'h6 == _T_9154) begin // @[FanCtrl.scala 753:46]
      r_reduction_sel_6 <= 2'h0; // @[FanCtrl.scala 753:46]
    end else begin
      r_reduction_sel_6 <= _GEN_91705;
    end
    if (reset) begin // @[FanCtrl.scala 21:34]
      r_reduction_sel_7 <= 2'h0; // @[FanCtrl.scala 21:34]
    end else if (r_valid_1) begin // @[FanCtrl.scala 745:33]
      if (_GEN_90400 == _GEN_90621) begin // @[FanCtrl.scala 746:70]
        if (5'h7 == _T_9154) begin // @[FanCtrl.scala 747:46]
          r_reduction_sel_7 <= 2'h3; // @[FanCtrl.scala 747:46]
        end else begin
          r_reduction_sel_7 <= _GEN_91706;
        end
      end else if (_GEN_90400 == _GEN_91866) begin // @[FanCtrl.scala 748:77]
        r_reduction_sel_7 <= _GEN_91874;
      end else begin
        r_reduction_sel_7 <= _GEN_91998;
      end
    end else if (5'h7 == _T_9154) begin // @[FanCtrl.scala 753:46]
      r_reduction_sel_7 <= 2'h0; // @[FanCtrl.scala 753:46]
    end else begin
      r_reduction_sel_7 <= _GEN_91706;
    end
    if (reset) begin // @[FanCtrl.scala 21:34]
      r_reduction_sel_8 <= 2'h0; // @[FanCtrl.scala 21:34]
    end else if (r_valid_1) begin // @[FanCtrl.scala 745:33]
      if (_GEN_90400 == _GEN_90621) begin // @[FanCtrl.scala 746:70]
        if (5'h8 == _T_9154) begin // @[FanCtrl.scala 747:46]
          r_reduction_sel_8 <= 2'h3; // @[FanCtrl.scala 747:46]
        end else begin
          r_reduction_sel_8 <= _GEN_91707;
        end
      end else if (_GEN_90400 == _GEN_91866) begin // @[FanCtrl.scala 748:77]
        r_reduction_sel_8 <= _GEN_91875;
      end else begin
        r_reduction_sel_8 <= _GEN_91999;
      end
    end else if (5'h8 == _T_9154) begin // @[FanCtrl.scala 753:46]
      r_reduction_sel_8 <= 2'h0; // @[FanCtrl.scala 753:46]
    end else begin
      r_reduction_sel_8 <= _GEN_91707;
    end
    if (reset) begin // @[FanCtrl.scala 21:34]
      r_reduction_sel_9 <= 2'h0; // @[FanCtrl.scala 21:34]
    end else if (r_valid_1) begin // @[FanCtrl.scala 745:33]
      if (_GEN_90400 == _GEN_90621) begin // @[FanCtrl.scala 746:70]
        if (5'h9 == _T_9154) begin // @[FanCtrl.scala 747:46]
          r_reduction_sel_9 <= 2'h3; // @[FanCtrl.scala 747:46]
        end else begin
          r_reduction_sel_9 <= _GEN_91708;
        end
      end else if (_GEN_90400 == _GEN_91866) begin // @[FanCtrl.scala 748:77]
        r_reduction_sel_9 <= _GEN_91876;
      end else begin
        r_reduction_sel_9 <= _GEN_92000;
      end
    end else if (5'h9 == _T_9154) begin // @[FanCtrl.scala 753:46]
      r_reduction_sel_9 <= 2'h0; // @[FanCtrl.scala 753:46]
    end else begin
      r_reduction_sel_9 <= _GEN_91708;
    end
    if (reset) begin // @[FanCtrl.scala 21:34]
      r_reduction_sel_10 <= 2'h0; // @[FanCtrl.scala 21:34]
    end else if (r_valid_1) begin // @[FanCtrl.scala 745:33]
      if (_GEN_90400 == _GEN_90621) begin // @[FanCtrl.scala 746:70]
        if (5'ha == _T_9154) begin // @[FanCtrl.scala 747:46]
          r_reduction_sel_10 <= 2'h3; // @[FanCtrl.scala 747:46]
        end else begin
          r_reduction_sel_10 <= _GEN_91709;
        end
      end else if (_GEN_90400 == _GEN_91866) begin // @[FanCtrl.scala 748:77]
        r_reduction_sel_10 <= _GEN_91877;
      end else begin
        r_reduction_sel_10 <= _GEN_92001;
      end
    end else if (5'ha == _T_9154) begin // @[FanCtrl.scala 753:46]
      r_reduction_sel_10 <= 2'h0; // @[FanCtrl.scala 753:46]
    end else begin
      r_reduction_sel_10 <= _GEN_91709;
    end
    if (reset) begin // @[FanCtrl.scala 21:34]
      r_reduction_sel_11 <= 2'h0; // @[FanCtrl.scala 21:34]
    end else if (r_valid_1) begin // @[FanCtrl.scala 745:33]
      if (_GEN_90400 == _GEN_90621) begin // @[FanCtrl.scala 746:70]
        if (5'hb == _T_9154) begin // @[FanCtrl.scala 747:46]
          r_reduction_sel_11 <= 2'h3; // @[FanCtrl.scala 747:46]
        end else begin
          r_reduction_sel_11 <= _GEN_91710;
        end
      end else if (_GEN_90400 == _GEN_91866) begin // @[FanCtrl.scala 748:77]
        r_reduction_sel_11 <= _GEN_91878;
      end else begin
        r_reduction_sel_11 <= _GEN_92002;
      end
    end else if (5'hb == _T_9154) begin // @[FanCtrl.scala 753:46]
      r_reduction_sel_11 <= 2'h0; // @[FanCtrl.scala 753:46]
    end else begin
      r_reduction_sel_11 <= _GEN_91710;
    end
    if (reset) begin // @[FanCtrl.scala 21:34]
      r_reduction_sel_12 <= 2'h0; // @[FanCtrl.scala 21:34]
    end else if (r_valid_1) begin // @[FanCtrl.scala 745:33]
      if (_GEN_90400 == _GEN_90621) begin // @[FanCtrl.scala 746:70]
        if (5'hc == _T_9154) begin // @[FanCtrl.scala 747:46]
          r_reduction_sel_12 <= 2'h3; // @[FanCtrl.scala 747:46]
        end else begin
          r_reduction_sel_12 <= _GEN_91711;
        end
      end else if (_GEN_90400 == _GEN_91866) begin // @[FanCtrl.scala 748:77]
        r_reduction_sel_12 <= _GEN_91879;
      end else begin
        r_reduction_sel_12 <= _GEN_92003;
      end
    end else if (5'hc == _T_9154) begin // @[FanCtrl.scala 753:46]
      r_reduction_sel_12 <= 2'h0; // @[FanCtrl.scala 753:46]
    end else begin
      r_reduction_sel_12 <= _GEN_91711;
    end
    if (reset) begin // @[FanCtrl.scala 21:34]
      r_reduction_sel_13 <= 2'h0; // @[FanCtrl.scala 21:34]
    end else if (r_valid_1) begin // @[FanCtrl.scala 745:33]
      if (_GEN_90400 == _GEN_90621) begin // @[FanCtrl.scala 746:70]
        if (5'hd == _T_9154) begin // @[FanCtrl.scala 747:46]
          r_reduction_sel_13 <= 2'h3; // @[FanCtrl.scala 747:46]
        end else begin
          r_reduction_sel_13 <= _GEN_91712;
        end
      end else if (_GEN_90400 == _GEN_91866) begin // @[FanCtrl.scala 748:77]
        r_reduction_sel_13 <= _GEN_91880;
      end else begin
        r_reduction_sel_13 <= _GEN_92004;
      end
    end else if (5'hd == _T_9154) begin // @[FanCtrl.scala 753:46]
      r_reduction_sel_13 <= 2'h0; // @[FanCtrl.scala 753:46]
    end else begin
      r_reduction_sel_13 <= _GEN_91712;
    end
    if (reset) begin // @[FanCtrl.scala 21:34]
      r_reduction_sel_14 <= 2'h0; // @[FanCtrl.scala 21:34]
    end else if (r_valid_1) begin // @[FanCtrl.scala 745:33]
      if (_GEN_90400 == _GEN_90621) begin // @[FanCtrl.scala 746:70]
        if (5'he == _T_9154) begin // @[FanCtrl.scala 747:46]
          r_reduction_sel_14 <= 2'h3; // @[FanCtrl.scala 747:46]
        end else begin
          r_reduction_sel_14 <= _GEN_91713;
        end
      end else if (_GEN_90400 == _GEN_91866) begin // @[FanCtrl.scala 748:77]
        r_reduction_sel_14 <= _GEN_91881;
      end else begin
        r_reduction_sel_14 <= _GEN_92005;
      end
    end else if (5'he == _T_9154) begin // @[FanCtrl.scala 753:46]
      r_reduction_sel_14 <= 2'h0; // @[FanCtrl.scala 753:46]
    end else begin
      r_reduction_sel_14 <= _GEN_91713;
    end
    if (reset) begin // @[FanCtrl.scala 21:34]
      r_reduction_sel_15 <= 2'h0; // @[FanCtrl.scala 21:34]
    end else if (r_valid_1) begin // @[FanCtrl.scala 745:33]
      if (_GEN_90400 == _GEN_90621) begin // @[FanCtrl.scala 746:70]
        if (5'hf == _T_9154) begin // @[FanCtrl.scala 747:46]
          r_reduction_sel_15 <= 2'h3; // @[FanCtrl.scala 747:46]
        end else begin
          r_reduction_sel_15 <= _GEN_91714;
        end
      end else if (_GEN_90400 == _GEN_91866) begin // @[FanCtrl.scala 748:77]
        r_reduction_sel_15 <= _GEN_91882;
      end else begin
        r_reduction_sel_15 <= _GEN_92006;
      end
    end else if (5'hf == _T_9154) begin // @[FanCtrl.scala 753:46]
      r_reduction_sel_15 <= 2'h0; // @[FanCtrl.scala 753:46]
    end else begin
      r_reduction_sel_15 <= _GEN_91714;
    end
    if (reset) begin // @[FanCtrl.scala 21:34]
      r_reduction_sel_16 <= 2'h0; // @[FanCtrl.scala 21:34]
    end else if (r_valid_1) begin // @[FanCtrl.scala 745:33]
      if (_GEN_90400 == _GEN_90621) begin // @[FanCtrl.scala 746:70]
        if (5'h10 == _T_9154) begin // @[FanCtrl.scala 747:46]
          r_reduction_sel_16 <= 2'h3; // @[FanCtrl.scala 747:46]
        end else begin
          r_reduction_sel_16 <= _GEN_91715;
        end
      end else if (_GEN_90400 == _GEN_91866) begin // @[FanCtrl.scala 748:77]
        r_reduction_sel_16 <= _GEN_91883;
      end else begin
        r_reduction_sel_16 <= _GEN_92007;
      end
    end else if (5'h10 == _T_9154) begin // @[FanCtrl.scala 753:46]
      r_reduction_sel_16 <= 2'h0; // @[FanCtrl.scala 753:46]
    end else begin
      r_reduction_sel_16 <= _GEN_91715;
    end
    if (reset) begin // @[FanCtrl.scala 21:34]
      r_reduction_sel_17 <= 2'h0; // @[FanCtrl.scala 21:34]
    end else if (r_valid_1) begin // @[FanCtrl.scala 745:33]
      if (_GEN_90400 == _GEN_90621) begin // @[FanCtrl.scala 746:70]
        if (5'h11 == _T_9154) begin // @[FanCtrl.scala 747:46]
          r_reduction_sel_17 <= 2'h3; // @[FanCtrl.scala 747:46]
        end else begin
          r_reduction_sel_17 <= _GEN_91716;
        end
      end else if (_GEN_90400 == _GEN_91866) begin // @[FanCtrl.scala 748:77]
        r_reduction_sel_17 <= _GEN_91884;
      end else begin
        r_reduction_sel_17 <= _GEN_92008;
      end
    end else if (5'h11 == _T_9154) begin // @[FanCtrl.scala 753:46]
      r_reduction_sel_17 <= 2'h0; // @[FanCtrl.scala 753:46]
    end else begin
      r_reduction_sel_17 <= _GEN_91716;
    end
    if (reset) begin // @[FanCtrl.scala 21:34]
      r_reduction_sel_18 <= 2'h0; // @[FanCtrl.scala 21:34]
    end else if (r_valid_1) begin // @[FanCtrl.scala 745:33]
      if (_GEN_90400 == _GEN_90621) begin // @[FanCtrl.scala 746:70]
        if (5'h12 == _T_9154) begin // @[FanCtrl.scala 747:46]
          r_reduction_sel_18 <= 2'h3; // @[FanCtrl.scala 747:46]
        end else begin
          r_reduction_sel_18 <= _GEN_91717;
        end
      end else if (_GEN_90400 == _GEN_91866) begin // @[FanCtrl.scala 748:77]
        r_reduction_sel_18 <= _GEN_91885;
      end else begin
        r_reduction_sel_18 <= _GEN_92009;
      end
    end else if (5'h12 == _T_9154) begin // @[FanCtrl.scala 753:46]
      r_reduction_sel_18 <= 2'h0; // @[FanCtrl.scala 753:46]
    end else begin
      r_reduction_sel_18 <= _GEN_91717;
    end
    if (reset) begin // @[FanCtrl.scala 21:34]
      r_reduction_sel_19 <= 2'h0; // @[FanCtrl.scala 21:34]
    end else if (r_valid_1) begin // @[FanCtrl.scala 745:33]
      if (_GEN_90400 == _GEN_90621) begin // @[FanCtrl.scala 746:70]
        if (5'h13 == _T_9154) begin // @[FanCtrl.scala 747:46]
          r_reduction_sel_19 <= 2'h3; // @[FanCtrl.scala 747:46]
        end else begin
          r_reduction_sel_19 <= _GEN_91718;
        end
      end else if (_GEN_90400 == _GEN_91866) begin // @[FanCtrl.scala 748:77]
        r_reduction_sel_19 <= _GEN_91886;
      end else begin
        r_reduction_sel_19 <= _GEN_92010;
      end
    end else if (5'h13 == _T_9154) begin // @[FanCtrl.scala 753:46]
      r_reduction_sel_19 <= 2'h0; // @[FanCtrl.scala 753:46]
    end else begin
      r_reduction_sel_19 <= _GEN_91718;
    end
    if (reset) begin // @[FanCtrl.scala 23:33]
      r_add_lvl_0Reg_0 <= 1'h0; // @[FanCtrl.scala 23:33]
    end else begin
      r_add_lvl_0Reg_0 <= r_reduction_add_0; // @[FanCtrl.scala 762:20]
    end
    if (reset) begin // @[FanCtrl.scala 23:33]
      r_add_lvl_0Reg_1 <= 1'h0; // @[FanCtrl.scala 23:33]
    end else begin
      r_add_lvl_0Reg_1 <= r_reduction_add_1; // @[FanCtrl.scala 762:20]
    end
    if (reset) begin // @[FanCtrl.scala 23:33]
      r_add_lvl_0Reg_2 <= 1'h0; // @[FanCtrl.scala 23:33]
    end else begin
      r_add_lvl_0Reg_2 <= r_reduction_add_2; // @[FanCtrl.scala 762:20]
    end
    if (reset) begin // @[FanCtrl.scala 23:33]
      r_add_lvl_0Reg_3 <= 1'h0; // @[FanCtrl.scala 23:33]
    end else begin
      r_add_lvl_0Reg_3 <= r_reduction_add_3; // @[FanCtrl.scala 762:20]
    end
    if (reset) begin // @[FanCtrl.scala 23:33]
      r_add_lvl_0Reg_4 <= 1'h0; // @[FanCtrl.scala 23:33]
    end else begin
      r_add_lvl_0Reg_4 <= r_reduction_add_4; // @[FanCtrl.scala 762:20]
    end
    if (reset) begin // @[FanCtrl.scala 23:33]
      r_add_lvl_0Reg_5 <= 1'h0; // @[FanCtrl.scala 23:33]
    end else begin
      r_add_lvl_0Reg_5 <= r_reduction_add_5; // @[FanCtrl.scala 762:20]
    end
    if (reset) begin // @[FanCtrl.scala 23:33]
      r_add_lvl_0Reg_6 <= 1'h0; // @[FanCtrl.scala 23:33]
    end else begin
      r_add_lvl_0Reg_6 <= r_reduction_add_6; // @[FanCtrl.scala 762:20]
    end
    if (reset) begin // @[FanCtrl.scala 23:33]
      r_add_lvl_0Reg_7 <= 1'h0; // @[FanCtrl.scala 23:33]
    end else begin
      r_add_lvl_0Reg_7 <= r_reduction_add_7; // @[FanCtrl.scala 762:20]
    end
    if (reset) begin // @[FanCtrl.scala 23:33]
      r_add_lvl_0Reg_8 <= 1'h0; // @[FanCtrl.scala 23:33]
    end else begin
      r_add_lvl_0Reg_8 <= r_reduction_add_8; // @[FanCtrl.scala 762:20]
    end
    if (reset) begin // @[FanCtrl.scala 23:33]
      r_add_lvl_0Reg_9 <= 1'h0; // @[FanCtrl.scala 23:33]
    end else begin
      r_add_lvl_0Reg_9 <= r_reduction_add_9; // @[FanCtrl.scala 762:20]
    end
    if (reset) begin // @[FanCtrl.scala 23:33]
      r_add_lvl_0Reg_10 <= 1'h0; // @[FanCtrl.scala 23:33]
    end else begin
      r_add_lvl_0Reg_10 <= r_reduction_add_10; // @[FanCtrl.scala 762:20]
    end
    if (reset) begin // @[FanCtrl.scala 23:33]
      r_add_lvl_0Reg_11 <= 1'h0; // @[FanCtrl.scala 23:33]
    end else begin
      r_add_lvl_0Reg_11 <= r_reduction_add_11; // @[FanCtrl.scala 762:20]
    end
    if (reset) begin // @[FanCtrl.scala 23:33]
      r_add_lvl_0Reg_12 <= 1'h0; // @[FanCtrl.scala 23:33]
    end else begin
      r_add_lvl_0Reg_12 <= r_reduction_add_12; // @[FanCtrl.scala 762:20]
    end
    if (reset) begin // @[FanCtrl.scala 23:33]
      r_add_lvl_0Reg_13 <= 1'h0; // @[FanCtrl.scala 23:33]
    end else begin
      r_add_lvl_0Reg_13 <= r_reduction_add_13; // @[FanCtrl.scala 762:20]
    end
    if (reset) begin // @[FanCtrl.scala 23:33]
      r_add_lvl_0Reg_14 <= 1'h0; // @[FanCtrl.scala 23:33]
    end else begin
      r_add_lvl_0Reg_14 <= r_reduction_add_14; // @[FanCtrl.scala 762:20]
    end
    if (reset) begin // @[FanCtrl.scala 23:33]
      r_add_lvl_0Reg_15 <= 1'h0; // @[FanCtrl.scala 23:33]
    end else begin
      r_add_lvl_0Reg_15 <= r_reduction_add_15; // @[FanCtrl.scala 762:20]
    end
    if (reset) begin // @[FanCtrl.scala 24:33]
      r_add_lvl_1Reg_8 <= 1'h0; // @[FanCtrl.scala 24:33]
    end else begin
      r_add_lvl_1Reg_8 <= r_reduction_add_16; // @[FanCtrl.scala 781:20]
    end
    if (reset) begin // @[FanCtrl.scala 24:33]
      r_add_lvl_1Reg_9 <= 1'h0; // @[FanCtrl.scala 24:33]
    end else begin
      r_add_lvl_1Reg_9 <= r_reduction_add_17; // @[FanCtrl.scala 781:20]
    end
    if (reset) begin // @[FanCtrl.scala 24:33]
      r_add_lvl_1Reg_10 <= 1'h0; // @[FanCtrl.scala 24:33]
    end else begin
      r_add_lvl_1Reg_10 <= r_reduction_add_18; // @[FanCtrl.scala 781:20]
    end
    if (reset) begin // @[FanCtrl.scala 24:33]
      r_add_lvl_1Reg_11 <= 1'h0; // @[FanCtrl.scala 24:33]
    end else begin
      r_add_lvl_1Reg_11 <= r_reduction_add_19; // @[FanCtrl.scala 781:20]
    end
    if (reset) begin // @[FanCtrl.scala 24:33]
      r_add_lvl_1Reg_12 <= 1'h0; // @[FanCtrl.scala 24:33]
    end else begin
      r_add_lvl_1Reg_12 <= r_reduction_add_20; // @[FanCtrl.scala 781:20]
    end
    if (reset) begin // @[FanCtrl.scala 24:33]
      r_add_lvl_1Reg_13 <= 1'h0; // @[FanCtrl.scala 24:33]
    end else begin
      r_add_lvl_1Reg_13 <= r_reduction_add_21; // @[FanCtrl.scala 781:20]
    end
    if (reset) begin // @[FanCtrl.scala 24:33]
      r_add_lvl_1Reg_14 <= 1'h0; // @[FanCtrl.scala 24:33]
    end else begin
      r_add_lvl_1Reg_14 <= r_reduction_add_22; // @[FanCtrl.scala 781:20]
    end
    if (reset) begin // @[FanCtrl.scala 24:33]
      r_add_lvl_1Reg_15 <= 1'h0; // @[FanCtrl.scala 24:33]
    end else begin
      r_add_lvl_1Reg_15 <= r_reduction_add_23; // @[FanCtrl.scala 781:20]
    end
    if (reset) begin // @[FanCtrl.scala 25:33]
      r_add_lvl_2Reg_8 <= 1'h0; // @[FanCtrl.scala 25:33]
    end else begin
      r_add_lvl_2Reg_8 <= r_reduction_add_24; // @[FanCtrl.scala 802:20]
    end
    if (reset) begin // @[FanCtrl.scala 25:33]
      r_add_lvl_2Reg_9 <= 1'h0; // @[FanCtrl.scala 25:33]
    end else begin
      r_add_lvl_2Reg_9 <= r_reduction_add_25; // @[FanCtrl.scala 802:20]
    end
    if (reset) begin // @[FanCtrl.scala 25:33]
      r_add_lvl_2Reg_10 <= 1'h0; // @[FanCtrl.scala 25:33]
    end else begin
      r_add_lvl_2Reg_10 <= r_reduction_add_26; // @[FanCtrl.scala 802:20]
    end
    if (reset) begin // @[FanCtrl.scala 25:33]
      r_add_lvl_2Reg_11 <= 1'h0; // @[FanCtrl.scala 25:33]
    end else begin
      r_add_lvl_2Reg_11 <= r_reduction_add_27; // @[FanCtrl.scala 802:20]
    end
    if (reset) begin // @[FanCtrl.scala 26:33]
      r_add_lvl_3Reg_6 <= 1'h0; // @[FanCtrl.scala 26:33]
    end else begin
      r_add_lvl_3Reg_6 <= r_reduction_add_28; // @[FanCtrl.scala 817:20]
    end
    if (reset) begin // @[FanCtrl.scala 26:33]
      r_add_lvl_3Reg_7 <= 1'h0; // @[FanCtrl.scala 26:33]
    end else begin
      r_add_lvl_3Reg_7 <= r_reduction_add_29; // @[FanCtrl.scala 817:20]
    end
    if (reset) begin // @[FanCtrl.scala 27:33]
      r_add_lvl_4Reg_4 <= 1'h0; // @[FanCtrl.scala 27:33]
    end else begin
      r_add_lvl_4Reg_4 <= r_reduction_add_30; // @[FanCtrl.scala 829:20]
    end
    if (reset) begin // @[FanCtrl.scala 29:33]
      r_cmd_lvl_0Reg_0 <= 3'h0; // @[FanCtrl.scala 29:33]
    end else begin
      r_cmd_lvl_0Reg_0 <= r_reduction_cmd_0; // @[FanCtrl.scala 838:20]
    end
    if (reset) begin // @[FanCtrl.scala 29:33]
      r_cmd_lvl_0Reg_1 <= 3'h0; // @[FanCtrl.scala 29:33]
    end else begin
      r_cmd_lvl_0Reg_1 <= r_reduction_cmd_1; // @[FanCtrl.scala 838:20]
    end
    if (reset) begin // @[FanCtrl.scala 29:33]
      r_cmd_lvl_0Reg_2 <= 3'h0; // @[FanCtrl.scala 29:33]
    end else begin
      r_cmd_lvl_0Reg_2 <= r_reduction_cmd_2; // @[FanCtrl.scala 838:20]
    end
    if (reset) begin // @[FanCtrl.scala 29:33]
      r_cmd_lvl_0Reg_3 <= 3'h0; // @[FanCtrl.scala 29:33]
    end else begin
      r_cmd_lvl_0Reg_3 <= r_reduction_cmd_3; // @[FanCtrl.scala 838:20]
    end
    if (reset) begin // @[FanCtrl.scala 29:33]
      r_cmd_lvl_0Reg_4 <= 3'h0; // @[FanCtrl.scala 29:33]
    end else begin
      r_cmd_lvl_0Reg_4 <= r_reduction_cmd_4; // @[FanCtrl.scala 838:20]
    end
    if (reset) begin // @[FanCtrl.scala 29:33]
      r_cmd_lvl_0Reg_5 <= 3'h0; // @[FanCtrl.scala 29:33]
    end else begin
      r_cmd_lvl_0Reg_5 <= r_reduction_cmd_5; // @[FanCtrl.scala 838:20]
    end
    if (reset) begin // @[FanCtrl.scala 29:33]
      r_cmd_lvl_0Reg_6 <= 3'h0; // @[FanCtrl.scala 29:33]
    end else begin
      r_cmd_lvl_0Reg_6 <= r_reduction_cmd_6; // @[FanCtrl.scala 838:20]
    end
    if (reset) begin // @[FanCtrl.scala 29:33]
      r_cmd_lvl_0Reg_7 <= 3'h0; // @[FanCtrl.scala 29:33]
    end else begin
      r_cmd_lvl_0Reg_7 <= r_reduction_cmd_7; // @[FanCtrl.scala 838:20]
    end
    if (reset) begin // @[FanCtrl.scala 29:33]
      r_cmd_lvl_0Reg_8 <= 3'h0; // @[FanCtrl.scala 29:33]
    end else begin
      r_cmd_lvl_0Reg_8 <= r_reduction_cmd_8; // @[FanCtrl.scala 838:20]
    end
    if (reset) begin // @[FanCtrl.scala 29:33]
      r_cmd_lvl_0Reg_9 <= 3'h0; // @[FanCtrl.scala 29:33]
    end else begin
      r_cmd_lvl_0Reg_9 <= r_reduction_cmd_9; // @[FanCtrl.scala 838:20]
    end
    if (reset) begin // @[FanCtrl.scala 29:33]
      r_cmd_lvl_0Reg_10 <= 3'h0; // @[FanCtrl.scala 29:33]
    end else begin
      r_cmd_lvl_0Reg_10 <= r_reduction_cmd_10; // @[FanCtrl.scala 838:20]
    end
    if (reset) begin // @[FanCtrl.scala 29:33]
      r_cmd_lvl_0Reg_11 <= 3'h0; // @[FanCtrl.scala 29:33]
    end else begin
      r_cmd_lvl_0Reg_11 <= r_reduction_cmd_11; // @[FanCtrl.scala 838:20]
    end
    if (reset) begin // @[FanCtrl.scala 29:33]
      r_cmd_lvl_0Reg_12 <= 3'h0; // @[FanCtrl.scala 29:33]
    end else begin
      r_cmd_lvl_0Reg_12 <= r_reduction_cmd_12; // @[FanCtrl.scala 838:20]
    end
    if (reset) begin // @[FanCtrl.scala 29:33]
      r_cmd_lvl_0Reg_13 <= 3'h0; // @[FanCtrl.scala 29:33]
    end else begin
      r_cmd_lvl_0Reg_13 <= r_reduction_cmd_13; // @[FanCtrl.scala 838:20]
    end
    if (reset) begin // @[FanCtrl.scala 29:33]
      r_cmd_lvl_0Reg_14 <= 3'h0; // @[FanCtrl.scala 29:33]
    end else begin
      r_cmd_lvl_0Reg_14 <= r_reduction_cmd_14; // @[FanCtrl.scala 838:20]
    end
    if (reset) begin // @[FanCtrl.scala 29:33]
      r_cmd_lvl_0Reg_15 <= 3'h0; // @[FanCtrl.scala 29:33]
    end else begin
      r_cmd_lvl_0Reg_15 <= r_reduction_cmd_15; // @[FanCtrl.scala 838:20]
    end
    if (reset) begin // @[FanCtrl.scala 30:33]
      r_cmd_lvl_1Reg_8 <= 3'h0; // @[FanCtrl.scala 30:33]
    end else begin
      r_cmd_lvl_1Reg_8 <= r_reduction_cmd_16; // @[FanCtrl.scala 859:20]
    end
    if (reset) begin // @[FanCtrl.scala 30:33]
      r_cmd_lvl_1Reg_9 <= 3'h0; // @[FanCtrl.scala 30:33]
    end else begin
      r_cmd_lvl_1Reg_9 <= r_reduction_cmd_17; // @[FanCtrl.scala 859:20]
    end
    if (reset) begin // @[FanCtrl.scala 30:33]
      r_cmd_lvl_1Reg_10 <= 3'h0; // @[FanCtrl.scala 30:33]
    end else begin
      r_cmd_lvl_1Reg_10 <= r_reduction_cmd_18; // @[FanCtrl.scala 859:20]
    end
    if (reset) begin // @[FanCtrl.scala 30:33]
      r_cmd_lvl_1Reg_11 <= 3'h0; // @[FanCtrl.scala 30:33]
    end else begin
      r_cmd_lvl_1Reg_11 <= r_reduction_cmd_19; // @[FanCtrl.scala 859:20]
    end
    if (reset) begin // @[FanCtrl.scala 30:33]
      r_cmd_lvl_1Reg_12 <= 3'h0; // @[FanCtrl.scala 30:33]
    end else begin
      r_cmd_lvl_1Reg_12 <= r_reduction_cmd_20; // @[FanCtrl.scala 859:20]
    end
    if (reset) begin // @[FanCtrl.scala 30:33]
      r_cmd_lvl_1Reg_13 <= 3'h0; // @[FanCtrl.scala 30:33]
    end else begin
      r_cmd_lvl_1Reg_13 <= r_reduction_cmd_21; // @[FanCtrl.scala 859:20]
    end
    if (reset) begin // @[FanCtrl.scala 30:33]
      r_cmd_lvl_1Reg_14 <= 3'h0; // @[FanCtrl.scala 30:33]
    end else begin
      r_cmd_lvl_1Reg_14 <= r_reduction_cmd_22; // @[FanCtrl.scala 859:20]
    end
    if (reset) begin // @[FanCtrl.scala 30:33]
      r_cmd_lvl_1Reg_15 <= 3'h0; // @[FanCtrl.scala 30:33]
    end else begin
      r_cmd_lvl_1Reg_15 <= r_reduction_cmd_23; // @[FanCtrl.scala 859:20]
    end
    if (reset) begin // @[FanCtrl.scala 31:33]
      r_cmd_lvl_2Reg_8 <= 3'h0; // @[FanCtrl.scala 31:33]
    end else begin
      r_cmd_lvl_2Reg_8 <= r_reduction_cmd_24; // @[FanCtrl.scala 878:20]
    end
    if (reset) begin // @[FanCtrl.scala 31:33]
      r_cmd_lvl_2Reg_9 <= 3'h0; // @[FanCtrl.scala 31:33]
    end else begin
      r_cmd_lvl_2Reg_9 <= r_reduction_cmd_25; // @[FanCtrl.scala 878:20]
    end
    if (reset) begin // @[FanCtrl.scala 31:33]
      r_cmd_lvl_2Reg_10 <= 3'h0; // @[FanCtrl.scala 31:33]
    end else begin
      r_cmd_lvl_2Reg_10 <= r_reduction_cmd_26; // @[FanCtrl.scala 878:20]
    end
    if (reset) begin // @[FanCtrl.scala 31:33]
      r_cmd_lvl_2Reg_11 <= 3'h0; // @[FanCtrl.scala 31:33]
    end else begin
      r_cmd_lvl_2Reg_11 <= r_reduction_cmd_27; // @[FanCtrl.scala 878:20]
    end
    if (reset) begin // @[FanCtrl.scala 32:33]
      r_cmd_lvl_3Reg_6 <= 3'h0; // @[FanCtrl.scala 32:33]
    end else begin
      r_cmd_lvl_3Reg_6 <= r_reduction_cmd_28; // @[FanCtrl.scala 893:20]
    end
    if (reset) begin // @[FanCtrl.scala 32:33]
      r_cmd_lvl_3Reg_7 <= 3'h0; // @[FanCtrl.scala 32:33]
    end else begin
      r_cmd_lvl_3Reg_7 <= r_reduction_cmd_29; // @[FanCtrl.scala 893:20]
    end
    if (reset) begin // @[FanCtrl.scala 33:33]
      r_cmd_lvl_4Reg_4 <= 3'h0; // @[FanCtrl.scala 33:33]
    end else begin
      r_cmd_lvl_4Reg_4 <= r_reduction_cmd_30; // @[FanCtrl.scala 904:20]
    end
    if (reset) begin // @[FanCtrl.scala 35:33]
      r_sel_lvl_2Reg_16 <= 2'h0; // @[FanCtrl.scala 35:33]
    end else begin
      r_sel_lvl_2Reg_16 <= r_reduction_sel_0; // @[FanCtrl.scala 912:21]
    end
    if (reset) begin // @[FanCtrl.scala 35:33]
      r_sel_lvl_2Reg_17 <= 2'h0; // @[FanCtrl.scala 35:33]
    end else begin
      r_sel_lvl_2Reg_17 <= r_reduction_sel_1; // @[FanCtrl.scala 912:21]
    end
    if (reset) begin // @[FanCtrl.scala 35:33]
      r_sel_lvl_2Reg_18 <= 2'h0; // @[FanCtrl.scala 35:33]
    end else begin
      r_sel_lvl_2Reg_18 <= r_reduction_sel_2; // @[FanCtrl.scala 912:21]
    end
    if (reset) begin // @[FanCtrl.scala 35:33]
      r_sel_lvl_2Reg_19 <= 2'h0; // @[FanCtrl.scala 35:33]
    end else begin
      r_sel_lvl_2Reg_19 <= r_reduction_sel_3; // @[FanCtrl.scala 912:21]
    end
    if (reset) begin // @[FanCtrl.scala 35:33]
      r_sel_lvl_2Reg_20 <= 2'h0; // @[FanCtrl.scala 35:33]
    end else begin
      r_sel_lvl_2Reg_20 <= r_reduction_sel_4; // @[FanCtrl.scala 912:21]
    end
    if (reset) begin // @[FanCtrl.scala 35:33]
      r_sel_lvl_2Reg_21 <= 2'h0; // @[FanCtrl.scala 35:33]
    end else begin
      r_sel_lvl_2Reg_21 <= r_reduction_sel_5; // @[FanCtrl.scala 912:21]
    end
    if (reset) begin // @[FanCtrl.scala 35:33]
      r_sel_lvl_2Reg_22 <= 2'h0; // @[FanCtrl.scala 35:33]
    end else begin
      r_sel_lvl_2Reg_22 <= r_reduction_sel_6; // @[FanCtrl.scala 912:21]
    end
    if (reset) begin // @[FanCtrl.scala 35:33]
      r_sel_lvl_2Reg_23 <= 2'h0; // @[FanCtrl.scala 35:33]
    end else begin
      r_sel_lvl_2Reg_23 <= r_reduction_sel_7; // @[FanCtrl.scala 912:21]
    end
    if (reset) begin // @[FanCtrl.scala 36:33]
      r_sel_lvl_3Reg_24 <= 2'h0; // @[FanCtrl.scala 36:33]
    end else begin
      r_sel_lvl_3Reg_24 <= r_reduction_sel_8; // @[FanCtrl.scala 940:20]
    end
    if (reset) begin // @[FanCtrl.scala 36:33]
      r_sel_lvl_3Reg_25 <= 2'h0; // @[FanCtrl.scala 36:33]
    end else begin
      r_sel_lvl_3Reg_25 <= r_reduction_sel_9; // @[FanCtrl.scala 940:20]
    end
    if (reset) begin // @[FanCtrl.scala 36:33]
      r_sel_lvl_3Reg_26 <= 2'h0; // @[FanCtrl.scala 36:33]
    end else begin
      r_sel_lvl_3Reg_26 <= r_reduction_sel_10; // @[FanCtrl.scala 940:20]
    end
    if (reset) begin // @[FanCtrl.scala 36:33]
      r_sel_lvl_3Reg_27 <= 2'h0; // @[FanCtrl.scala 36:33]
    end else begin
      r_sel_lvl_3Reg_27 <= r_reduction_sel_11; // @[FanCtrl.scala 940:20]
    end
    if (reset) begin // @[FanCtrl.scala 36:33]
      r_sel_lvl_3Reg_28 <= 2'h0; // @[FanCtrl.scala 36:33]
    end else begin
      r_sel_lvl_3Reg_28 <= r_reduction_sel_12; // @[FanCtrl.scala 940:20]
    end
    if (reset) begin // @[FanCtrl.scala 36:33]
      r_sel_lvl_3Reg_29 <= 2'h0; // @[FanCtrl.scala 36:33]
    end else begin
      r_sel_lvl_3Reg_29 <= r_reduction_sel_13; // @[FanCtrl.scala 940:20]
    end
    if (reset) begin // @[FanCtrl.scala 36:33]
      r_sel_lvl_3Reg_30 <= 2'h0; // @[FanCtrl.scala 36:33]
    end else begin
      r_sel_lvl_3Reg_30 <= r_reduction_sel_14; // @[FanCtrl.scala 940:20]
    end
    if (reset) begin // @[FanCtrl.scala 36:33]
      r_sel_lvl_3Reg_31 <= 2'h0; // @[FanCtrl.scala 36:33]
    end else begin
      r_sel_lvl_3Reg_31 <= r_reduction_sel_15; // @[FanCtrl.scala 940:20]
    end
    if (reset) begin // @[FanCtrl.scala 37:33]
      r_sel_lvl_4Reg_16 <= 2'h0; // @[FanCtrl.scala 37:33]
    end else begin
      r_sel_lvl_4Reg_16 <= r_reduction_sel_16; // @[FanCtrl.scala 974:20]
    end
    if (reset) begin // @[FanCtrl.scala 37:33]
      r_sel_lvl_4Reg_17 <= 2'h0; // @[FanCtrl.scala 37:33]
    end else begin
      r_sel_lvl_4Reg_17 <= r_reduction_sel_17; // @[FanCtrl.scala 974:20]
    end
    if (reset) begin // @[FanCtrl.scala 37:33]
      r_sel_lvl_4Reg_18 <= 2'h0; // @[FanCtrl.scala 37:33]
    end else begin
      r_sel_lvl_4Reg_18 <= r_reduction_sel_18; // @[FanCtrl.scala 974:20]
    end
    if (reset) begin // @[FanCtrl.scala 37:33]
      r_sel_lvl_4Reg_19 <= 2'h0; // @[FanCtrl.scala 37:33]
    end else begin
      r_sel_lvl_4Reg_19 <= r_reduction_sel_19; // @[FanCtrl.scala 974:20]
    end
    if (reset) begin // @[FanCtrl.scala 40:23]
      w_vn_3 <= 5'h0; // @[FanCtrl.scala 40:23]
    end else begin
      w_vn_3 <= 5'h1d; // @[FanCtrl.scala 43:10]
    end
    if (reset) begin // @[FanCtrl.scala 40:23]
      w_vn_4 <= 5'h0; // @[FanCtrl.scala 40:23]
    end else begin
      w_vn_4 <= 5'h1d; // @[FanCtrl.scala 43:10]
    end
    if (reset) begin // @[FanCtrl.scala 40:23]
      w_vn_7 <= 5'h0; // @[FanCtrl.scala 40:23]
    end else begin
      w_vn_7 <= 5'h17; // @[FanCtrl.scala 43:10]
    end
    if (reset) begin // @[FanCtrl.scala 40:23]
      w_vn_8 <= 5'h0; // @[FanCtrl.scala 40:23]
    end else begin
      w_vn_8 <= 5'h17; // @[FanCtrl.scala 43:10]
    end
    if (reset) begin // @[FanCtrl.scala 40:23]
      w_vn_11 <= 5'h0; // @[FanCtrl.scala 40:23]
    end else begin
      w_vn_11 <= 5'hf; // @[FanCtrl.scala 43:10]
    end
    if (reset) begin // @[FanCtrl.scala 40:23]
      w_vn_12 <= 5'h0; // @[FanCtrl.scala 40:23]
    end else begin
      w_vn_12 <= 5'hf; // @[FanCtrl.scala 43:10]
    end
    if (reset) begin // @[FanCtrl.scala 40:23]
      w_vn_13 <= 5'h0; // @[FanCtrl.scala 40:23]
    end else begin
      w_vn_13 <= 5'h18; // @[FanCtrl.scala 43:10]
    end
    if (reset) begin // @[FanCtrl.scala 40:23]
      w_vn_15 <= 5'h0; // @[FanCtrl.scala 40:23]
    end else begin
      w_vn_15 <= 5'h1e; // @[FanCtrl.scala 43:10]
    end
    if (reset) begin // @[FanCtrl.scala 40:23]
      w_vn_16 <= 5'h0; // @[FanCtrl.scala 40:23]
    end else begin
      w_vn_16 <= 5'h1e; // @[FanCtrl.scala 43:10]
    end
    if (reset) begin // @[FanCtrl.scala 40:23]
      w_vn_18 <= 5'h0; // @[FanCtrl.scala 40:23]
    end else begin
      w_vn_18 <= 5'h1f; // @[FanCtrl.scala 43:10]
    end
    if (reset) begin // @[FanCtrl.scala 40:23]
      w_vn_23 <= 5'h0; // @[FanCtrl.scala 40:23]
    end else begin
      w_vn_23 <= 5'h1f; // @[FanCtrl.scala 43:10]
    end
    if (reset) begin // @[FanCtrl.scala 40:23]
      w_vn_24 <= 5'h0; // @[FanCtrl.scala 40:23]
    end else begin
      w_vn_24 <= 5'h1f; // @[FanCtrl.scala 43:10]
    end
    if (reset) begin // @[FanCtrl.scala 41:26]
      r_valid_0 <= 1'h0; // @[FanCtrl.scala 41:26]
    end else begin
      r_valid_0 <= 1'h1;
    end
    if (reset) begin // @[FanCtrl.scala 41:26]
      r_valid_1 <= 1'h0; // @[FanCtrl.scala 41:26]
    end else begin
      r_valid_1 <= r_valid_0; // @[FanCtrl.scala 1006:24]
    end
    if (reset) begin // @[FanCtrl.scala 41:26]
      r_valid_2 <= 1'h0; // @[FanCtrl.scala 41:26]
    end else begin
      r_valid_2 <= r_valid_1; // @[FanCtrl.scala 1006:24]
    end
    if (reset) begin // @[FanCtrl.scala 41:26]
      r_valid_3 <= 1'h0; // @[FanCtrl.scala 41:26]
    end else begin
      r_valid_3 <= r_valid_2; // @[FanCtrl.scala 1006:24]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_reduction_add_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  r_reduction_add_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  r_reduction_add_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  r_reduction_add_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  r_reduction_add_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  r_reduction_add_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  r_reduction_add_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  r_reduction_add_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  r_reduction_add_8 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  r_reduction_add_9 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  r_reduction_add_10 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  r_reduction_add_11 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  r_reduction_add_12 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  r_reduction_add_13 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  r_reduction_add_14 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  r_reduction_add_15 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  r_reduction_add_16 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  r_reduction_add_17 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  r_reduction_add_18 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  r_reduction_add_19 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  r_reduction_add_20 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  r_reduction_add_21 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  r_reduction_add_22 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  r_reduction_add_23 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  r_reduction_add_24 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  r_reduction_add_25 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  r_reduction_add_26 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  r_reduction_add_27 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  r_reduction_add_28 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  r_reduction_add_29 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  r_reduction_add_30 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  r_reduction_cmd_0 = _RAND_31[2:0];
  _RAND_32 = {1{`RANDOM}};
  r_reduction_cmd_1 = _RAND_32[2:0];
  _RAND_33 = {1{`RANDOM}};
  r_reduction_cmd_2 = _RAND_33[2:0];
  _RAND_34 = {1{`RANDOM}};
  r_reduction_cmd_3 = _RAND_34[2:0];
  _RAND_35 = {1{`RANDOM}};
  r_reduction_cmd_4 = _RAND_35[2:0];
  _RAND_36 = {1{`RANDOM}};
  r_reduction_cmd_5 = _RAND_36[2:0];
  _RAND_37 = {1{`RANDOM}};
  r_reduction_cmd_6 = _RAND_37[2:0];
  _RAND_38 = {1{`RANDOM}};
  r_reduction_cmd_7 = _RAND_38[2:0];
  _RAND_39 = {1{`RANDOM}};
  r_reduction_cmd_8 = _RAND_39[2:0];
  _RAND_40 = {1{`RANDOM}};
  r_reduction_cmd_9 = _RAND_40[2:0];
  _RAND_41 = {1{`RANDOM}};
  r_reduction_cmd_10 = _RAND_41[2:0];
  _RAND_42 = {1{`RANDOM}};
  r_reduction_cmd_11 = _RAND_42[2:0];
  _RAND_43 = {1{`RANDOM}};
  r_reduction_cmd_12 = _RAND_43[2:0];
  _RAND_44 = {1{`RANDOM}};
  r_reduction_cmd_13 = _RAND_44[2:0];
  _RAND_45 = {1{`RANDOM}};
  r_reduction_cmd_14 = _RAND_45[2:0];
  _RAND_46 = {1{`RANDOM}};
  r_reduction_cmd_15 = _RAND_46[2:0];
  _RAND_47 = {1{`RANDOM}};
  r_reduction_cmd_16 = _RAND_47[2:0];
  _RAND_48 = {1{`RANDOM}};
  r_reduction_cmd_17 = _RAND_48[2:0];
  _RAND_49 = {1{`RANDOM}};
  r_reduction_cmd_18 = _RAND_49[2:0];
  _RAND_50 = {1{`RANDOM}};
  r_reduction_cmd_19 = _RAND_50[2:0];
  _RAND_51 = {1{`RANDOM}};
  r_reduction_cmd_20 = _RAND_51[2:0];
  _RAND_52 = {1{`RANDOM}};
  r_reduction_cmd_21 = _RAND_52[2:0];
  _RAND_53 = {1{`RANDOM}};
  r_reduction_cmd_22 = _RAND_53[2:0];
  _RAND_54 = {1{`RANDOM}};
  r_reduction_cmd_23 = _RAND_54[2:0];
  _RAND_55 = {1{`RANDOM}};
  r_reduction_cmd_24 = _RAND_55[2:0];
  _RAND_56 = {1{`RANDOM}};
  r_reduction_cmd_25 = _RAND_56[2:0];
  _RAND_57 = {1{`RANDOM}};
  r_reduction_cmd_26 = _RAND_57[2:0];
  _RAND_58 = {1{`RANDOM}};
  r_reduction_cmd_27 = _RAND_58[2:0];
  _RAND_59 = {1{`RANDOM}};
  r_reduction_cmd_28 = _RAND_59[2:0];
  _RAND_60 = {1{`RANDOM}};
  r_reduction_cmd_29 = _RAND_60[2:0];
  _RAND_61 = {1{`RANDOM}};
  r_reduction_cmd_30 = _RAND_61[2:0];
  _RAND_62 = {1{`RANDOM}};
  r_reduction_sel_0 = _RAND_62[1:0];
  _RAND_63 = {1{`RANDOM}};
  r_reduction_sel_1 = _RAND_63[1:0];
  _RAND_64 = {1{`RANDOM}};
  r_reduction_sel_2 = _RAND_64[1:0];
  _RAND_65 = {1{`RANDOM}};
  r_reduction_sel_3 = _RAND_65[1:0];
  _RAND_66 = {1{`RANDOM}};
  r_reduction_sel_4 = _RAND_66[1:0];
  _RAND_67 = {1{`RANDOM}};
  r_reduction_sel_5 = _RAND_67[1:0];
  _RAND_68 = {1{`RANDOM}};
  r_reduction_sel_6 = _RAND_68[1:0];
  _RAND_69 = {1{`RANDOM}};
  r_reduction_sel_7 = _RAND_69[1:0];
  _RAND_70 = {1{`RANDOM}};
  r_reduction_sel_8 = _RAND_70[1:0];
  _RAND_71 = {1{`RANDOM}};
  r_reduction_sel_9 = _RAND_71[1:0];
  _RAND_72 = {1{`RANDOM}};
  r_reduction_sel_10 = _RAND_72[1:0];
  _RAND_73 = {1{`RANDOM}};
  r_reduction_sel_11 = _RAND_73[1:0];
  _RAND_74 = {1{`RANDOM}};
  r_reduction_sel_12 = _RAND_74[1:0];
  _RAND_75 = {1{`RANDOM}};
  r_reduction_sel_13 = _RAND_75[1:0];
  _RAND_76 = {1{`RANDOM}};
  r_reduction_sel_14 = _RAND_76[1:0];
  _RAND_77 = {1{`RANDOM}};
  r_reduction_sel_15 = _RAND_77[1:0];
  _RAND_78 = {1{`RANDOM}};
  r_reduction_sel_16 = _RAND_78[1:0];
  _RAND_79 = {1{`RANDOM}};
  r_reduction_sel_17 = _RAND_79[1:0];
  _RAND_80 = {1{`RANDOM}};
  r_reduction_sel_18 = _RAND_80[1:0];
  _RAND_81 = {1{`RANDOM}};
  r_reduction_sel_19 = _RAND_81[1:0];
  _RAND_82 = {1{`RANDOM}};
  r_add_lvl_0Reg_0 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  r_add_lvl_0Reg_1 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  r_add_lvl_0Reg_2 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  r_add_lvl_0Reg_3 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  r_add_lvl_0Reg_4 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  r_add_lvl_0Reg_5 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  r_add_lvl_0Reg_6 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  r_add_lvl_0Reg_7 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  r_add_lvl_0Reg_8 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  r_add_lvl_0Reg_9 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  r_add_lvl_0Reg_10 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  r_add_lvl_0Reg_11 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  r_add_lvl_0Reg_12 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  r_add_lvl_0Reg_13 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  r_add_lvl_0Reg_14 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  r_add_lvl_0Reg_15 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  r_add_lvl_1Reg_8 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  r_add_lvl_1Reg_9 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  r_add_lvl_1Reg_10 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  r_add_lvl_1Reg_11 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  r_add_lvl_1Reg_12 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  r_add_lvl_1Reg_13 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  r_add_lvl_1Reg_14 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  r_add_lvl_1Reg_15 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  r_add_lvl_2Reg_8 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  r_add_lvl_2Reg_9 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  r_add_lvl_2Reg_10 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  r_add_lvl_2Reg_11 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  r_add_lvl_3Reg_6 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  r_add_lvl_3Reg_7 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  r_add_lvl_4Reg_4 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  r_cmd_lvl_0Reg_0 = _RAND_113[2:0];
  _RAND_114 = {1{`RANDOM}};
  r_cmd_lvl_0Reg_1 = _RAND_114[2:0];
  _RAND_115 = {1{`RANDOM}};
  r_cmd_lvl_0Reg_2 = _RAND_115[2:0];
  _RAND_116 = {1{`RANDOM}};
  r_cmd_lvl_0Reg_3 = _RAND_116[2:0];
  _RAND_117 = {1{`RANDOM}};
  r_cmd_lvl_0Reg_4 = _RAND_117[2:0];
  _RAND_118 = {1{`RANDOM}};
  r_cmd_lvl_0Reg_5 = _RAND_118[2:0];
  _RAND_119 = {1{`RANDOM}};
  r_cmd_lvl_0Reg_6 = _RAND_119[2:0];
  _RAND_120 = {1{`RANDOM}};
  r_cmd_lvl_0Reg_7 = _RAND_120[2:0];
  _RAND_121 = {1{`RANDOM}};
  r_cmd_lvl_0Reg_8 = _RAND_121[2:0];
  _RAND_122 = {1{`RANDOM}};
  r_cmd_lvl_0Reg_9 = _RAND_122[2:0];
  _RAND_123 = {1{`RANDOM}};
  r_cmd_lvl_0Reg_10 = _RAND_123[2:0];
  _RAND_124 = {1{`RANDOM}};
  r_cmd_lvl_0Reg_11 = _RAND_124[2:0];
  _RAND_125 = {1{`RANDOM}};
  r_cmd_lvl_0Reg_12 = _RAND_125[2:0];
  _RAND_126 = {1{`RANDOM}};
  r_cmd_lvl_0Reg_13 = _RAND_126[2:0];
  _RAND_127 = {1{`RANDOM}};
  r_cmd_lvl_0Reg_14 = _RAND_127[2:0];
  _RAND_128 = {1{`RANDOM}};
  r_cmd_lvl_0Reg_15 = _RAND_128[2:0];
  _RAND_129 = {1{`RANDOM}};
  r_cmd_lvl_1Reg_8 = _RAND_129[2:0];
  _RAND_130 = {1{`RANDOM}};
  r_cmd_lvl_1Reg_9 = _RAND_130[2:0];
  _RAND_131 = {1{`RANDOM}};
  r_cmd_lvl_1Reg_10 = _RAND_131[2:0];
  _RAND_132 = {1{`RANDOM}};
  r_cmd_lvl_1Reg_11 = _RAND_132[2:0];
  _RAND_133 = {1{`RANDOM}};
  r_cmd_lvl_1Reg_12 = _RAND_133[2:0];
  _RAND_134 = {1{`RANDOM}};
  r_cmd_lvl_1Reg_13 = _RAND_134[2:0];
  _RAND_135 = {1{`RANDOM}};
  r_cmd_lvl_1Reg_14 = _RAND_135[2:0];
  _RAND_136 = {1{`RANDOM}};
  r_cmd_lvl_1Reg_15 = _RAND_136[2:0];
  _RAND_137 = {1{`RANDOM}};
  r_cmd_lvl_2Reg_8 = _RAND_137[2:0];
  _RAND_138 = {1{`RANDOM}};
  r_cmd_lvl_2Reg_9 = _RAND_138[2:0];
  _RAND_139 = {1{`RANDOM}};
  r_cmd_lvl_2Reg_10 = _RAND_139[2:0];
  _RAND_140 = {1{`RANDOM}};
  r_cmd_lvl_2Reg_11 = _RAND_140[2:0];
  _RAND_141 = {1{`RANDOM}};
  r_cmd_lvl_3Reg_6 = _RAND_141[2:0];
  _RAND_142 = {1{`RANDOM}};
  r_cmd_lvl_3Reg_7 = _RAND_142[2:0];
  _RAND_143 = {1{`RANDOM}};
  r_cmd_lvl_4Reg_4 = _RAND_143[2:0];
  _RAND_144 = {1{`RANDOM}};
  r_sel_lvl_2Reg_16 = _RAND_144[1:0];
  _RAND_145 = {1{`RANDOM}};
  r_sel_lvl_2Reg_17 = _RAND_145[1:0];
  _RAND_146 = {1{`RANDOM}};
  r_sel_lvl_2Reg_18 = _RAND_146[1:0];
  _RAND_147 = {1{`RANDOM}};
  r_sel_lvl_2Reg_19 = _RAND_147[1:0];
  _RAND_148 = {1{`RANDOM}};
  r_sel_lvl_2Reg_20 = _RAND_148[1:0];
  _RAND_149 = {1{`RANDOM}};
  r_sel_lvl_2Reg_21 = _RAND_149[1:0];
  _RAND_150 = {1{`RANDOM}};
  r_sel_lvl_2Reg_22 = _RAND_150[1:0];
  _RAND_151 = {1{`RANDOM}};
  r_sel_lvl_2Reg_23 = _RAND_151[1:0];
  _RAND_152 = {1{`RANDOM}};
  r_sel_lvl_3Reg_24 = _RAND_152[1:0];
  _RAND_153 = {1{`RANDOM}};
  r_sel_lvl_3Reg_25 = _RAND_153[1:0];
  _RAND_154 = {1{`RANDOM}};
  r_sel_lvl_3Reg_26 = _RAND_154[1:0];
  _RAND_155 = {1{`RANDOM}};
  r_sel_lvl_3Reg_27 = _RAND_155[1:0];
  _RAND_156 = {1{`RANDOM}};
  r_sel_lvl_3Reg_28 = _RAND_156[1:0];
  _RAND_157 = {1{`RANDOM}};
  r_sel_lvl_3Reg_29 = _RAND_157[1:0];
  _RAND_158 = {1{`RANDOM}};
  r_sel_lvl_3Reg_30 = _RAND_158[1:0];
  _RAND_159 = {1{`RANDOM}};
  r_sel_lvl_3Reg_31 = _RAND_159[1:0];
  _RAND_160 = {1{`RANDOM}};
  r_sel_lvl_4Reg_16 = _RAND_160[1:0];
  _RAND_161 = {1{`RANDOM}};
  r_sel_lvl_4Reg_17 = _RAND_161[1:0];
  _RAND_162 = {1{`RANDOM}};
  r_sel_lvl_4Reg_18 = _RAND_162[1:0];
  _RAND_163 = {1{`RANDOM}};
  r_sel_lvl_4Reg_19 = _RAND_163[1:0];
  _RAND_164 = {1{`RANDOM}};
  w_vn_3 = _RAND_164[4:0];
  _RAND_165 = {1{`RANDOM}};
  w_vn_4 = _RAND_165[4:0];
  _RAND_166 = {1{`RANDOM}};
  w_vn_7 = _RAND_166[4:0];
  _RAND_167 = {1{`RANDOM}};
  w_vn_8 = _RAND_167[4:0];
  _RAND_168 = {1{`RANDOM}};
  w_vn_11 = _RAND_168[4:0];
  _RAND_169 = {1{`RANDOM}};
  w_vn_12 = _RAND_169[4:0];
  _RAND_170 = {1{`RANDOM}};
  w_vn_13 = _RAND_170[4:0];
  _RAND_171 = {1{`RANDOM}};
  w_vn_15 = _RAND_171[4:0];
  _RAND_172 = {1{`RANDOM}};
  w_vn_16 = _RAND_172[4:0];
  _RAND_173 = {1{`RANDOM}};
  w_vn_18 = _RAND_173[4:0];
  _RAND_174 = {1{`RANDOM}};
  w_vn_23 = _RAND_174[4:0];
  _RAND_175 = {1{`RANDOM}};
  w_vn_24 = _RAND_175[4:0];
  _RAND_176 = {1{`RANDOM}};
  r_valid_0 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  r_valid_1 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  r_valid_2 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  r_valid_3 = _RAND_179[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module InputSwitch(
  output [15:0] io_y,
  output [15:0] io_z,
  input  [15:0] io_in
);
  assign io_y = io_in; // @[Switches.scala 13:8]
  assign io_z = io_in; // @[Switches.scala 14:8]
endmodule
module BenesMux(
  output [15:0] io_o,
  input  [15:0] io_a
);
  assign io_o = io_a; // @[Switches.scala 65:14]
endmodule
module OutputSwitch(
  output [15:0] io_y,
  input  [15:0] io_in0
);
  wire [15:0] mux0_io_o; // @[Switches.scala 26:20]
  wire [15:0] mux0_io_a; // @[Switches.scala 26:20]
  BenesMux mux0 ( // @[Switches.scala 26:20]
    .io_o(mux0_io_o),
    .io_a(mux0_io_a)
  );
  assign io_y = mux0_io_o; // @[Switches.scala 30:8]
  assign mux0_io_a = io_in0; // @[Switches.scala 27:13]
endmodule
module Switch(
  output [15:0] io_y,
  output [15:0] io_z,
  input  [15:0] io_in0
);
  wire [15:0] mux0_io_o; // @[Switches.scala 44:20]
  wire [15:0] mux0_io_a; // @[Switches.scala 44:20]
  wire [15:0] mux1_io_o; // @[Switches.scala 45:20]
  wire [15:0] mux1_io_a; // @[Switches.scala 45:20]
  BenesMux mux0 ( // @[Switches.scala 44:20]
    .io_o(mux0_io_o),
    .io_a(mux0_io_a)
  );
  BenesMux mux1 ( // @[Switches.scala 45:20]
    .io_o(mux1_io_o),
    .io_a(mux1_io_a)
  );
  assign io_y = mux0_io_o; // @[Switches.scala 52:8]
  assign io_z = mux1_io_o; // @[Switches.scala 53:8]
  assign mux0_io_a = io_in0; // @[Switches.scala 46:13]
  assign mux1_io_a = io_in0; // @[Switches.scala 49:13]
endmodule
module Benes(
  input         clock,
  input         reset,
  output [15:0] io_o_dist_bus2_0,
  output [15:0] io_o_dist_bus2_1,
  output [15:0] io_o_dist_bus2_2,
  output [15:0] io_o_dist_bus2_3,
  output [15:0] io_o_dist_bus2_4,
  output [15:0] io_o_dist_bus2_5,
  output [15:0] io_o_dist_bus2_6,
  output [15:0] io_o_dist_bus2_7,
  output [15:0] io_o_dist_bus2_8,
  output [15:0] io_o_dist_bus2_9,
  output [15:0] io_o_dist_bus2_10,
  output [15:0] io_o_dist_bus2_11,
  output [15:0] io_o_dist_bus2_12,
  output [15:0] io_o_dist_bus2_13,
  output [15:0] io_o_dist_bus2_14,
  output [15:0] io_o_dist_bus2_15,
  output [15:0] io_o_dist_bus2_16,
  output [15:0] io_o_dist_bus2_17,
  output [15:0] io_o_dist_bus2_18,
  output [15:0] io_o_dist_bus2_19,
  output [15:0] io_o_dist_bus2_20,
  output [15:0] io_o_dist_bus2_21,
  output [15:0] io_o_dist_bus2_22,
  output [15:0] io_o_dist_bus2_23,
  output [15:0] io_o_dist_bus2_24,
  output [15:0] io_o_dist_bus2_25,
  output [15:0] io_o_dist_bus2_26,
  output [15:0] io_o_dist_bus2_27,
  output [15:0] io_o_dist_bus2_28,
  output [15:0] io_o_dist_bus2_29,
  output [15:0] io_o_dist_bus2_30,
  output [15:0] io_o_dist_bus2_31
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] in_switch_io_y; // @[Benes.scala 90:27]
  wire [15:0] in_switch_io_z; // @[Benes.scala 90:27]
  wire [15:0] in_switch_io_in; // @[Benes.scala 90:27]
  wire [15:0] in_switch_1_io_y; // @[Benes.scala 90:27]
  wire [15:0] in_switch_1_io_z; // @[Benes.scala 90:27]
  wire [15:0] in_switch_1_io_in; // @[Benes.scala 90:27]
  wire [15:0] in_switch_2_io_y; // @[Benes.scala 90:27]
  wire [15:0] in_switch_2_io_z; // @[Benes.scala 90:27]
  wire [15:0] in_switch_2_io_in; // @[Benes.scala 90:27]
  wire [15:0] in_switch_3_io_y; // @[Benes.scala 90:27]
  wire [15:0] in_switch_3_io_z; // @[Benes.scala 90:27]
  wire [15:0] in_switch_3_io_in; // @[Benes.scala 90:27]
  wire [15:0] in_switch_4_io_y; // @[Benes.scala 90:27]
  wire [15:0] in_switch_4_io_z; // @[Benes.scala 90:27]
  wire [15:0] in_switch_4_io_in; // @[Benes.scala 90:27]
  wire [15:0] in_switch_5_io_y; // @[Benes.scala 90:27]
  wire [15:0] in_switch_5_io_z; // @[Benes.scala 90:27]
  wire [15:0] in_switch_5_io_in; // @[Benes.scala 90:27]
  wire [15:0] in_switch_6_io_y; // @[Benes.scala 90:27]
  wire [15:0] in_switch_6_io_z; // @[Benes.scala 90:27]
  wire [15:0] in_switch_6_io_in; // @[Benes.scala 90:27]
  wire [15:0] in_switch_7_io_y; // @[Benes.scala 90:27]
  wire [15:0] in_switch_7_io_z; // @[Benes.scala 90:27]
  wire [15:0] in_switch_7_io_in; // @[Benes.scala 90:27]
  wire [15:0] in_switch_8_io_y; // @[Benes.scala 90:27]
  wire [15:0] in_switch_8_io_z; // @[Benes.scala 90:27]
  wire [15:0] in_switch_8_io_in; // @[Benes.scala 90:27]
  wire [15:0] in_switch_9_io_y; // @[Benes.scala 90:27]
  wire [15:0] in_switch_9_io_z; // @[Benes.scala 90:27]
  wire [15:0] in_switch_9_io_in; // @[Benes.scala 90:27]
  wire [15:0] in_switch_10_io_y; // @[Benes.scala 90:27]
  wire [15:0] in_switch_10_io_z; // @[Benes.scala 90:27]
  wire [15:0] in_switch_10_io_in; // @[Benes.scala 90:27]
  wire [15:0] in_switch_11_io_y; // @[Benes.scala 90:27]
  wire [15:0] in_switch_11_io_z; // @[Benes.scala 90:27]
  wire [15:0] in_switch_11_io_in; // @[Benes.scala 90:27]
  wire [15:0] in_switch_12_io_y; // @[Benes.scala 90:27]
  wire [15:0] in_switch_12_io_z; // @[Benes.scala 90:27]
  wire [15:0] in_switch_12_io_in; // @[Benes.scala 90:27]
  wire [15:0] in_switch_13_io_y; // @[Benes.scala 90:27]
  wire [15:0] in_switch_13_io_z; // @[Benes.scala 90:27]
  wire [15:0] in_switch_13_io_in; // @[Benes.scala 90:27]
  wire [15:0] in_switch_14_io_y; // @[Benes.scala 90:27]
  wire [15:0] in_switch_14_io_z; // @[Benes.scala 90:27]
  wire [15:0] in_switch_14_io_in; // @[Benes.scala 90:27]
  wire [15:0] in_switch_15_io_y; // @[Benes.scala 90:27]
  wire [15:0] in_switch_15_io_z; // @[Benes.scala 90:27]
  wire [15:0] in_switch_15_io_in; // @[Benes.scala 90:27]
  wire [15:0] in_switch_16_io_y; // @[Benes.scala 90:27]
  wire [15:0] in_switch_16_io_z; // @[Benes.scala 90:27]
  wire [15:0] in_switch_16_io_in; // @[Benes.scala 90:27]
  wire [15:0] in_switch_17_io_y; // @[Benes.scala 90:27]
  wire [15:0] in_switch_17_io_z; // @[Benes.scala 90:27]
  wire [15:0] in_switch_17_io_in; // @[Benes.scala 90:27]
  wire [15:0] in_switch_18_io_y; // @[Benes.scala 90:27]
  wire [15:0] in_switch_18_io_z; // @[Benes.scala 90:27]
  wire [15:0] in_switch_18_io_in; // @[Benes.scala 90:27]
  wire [15:0] in_switch_19_io_y; // @[Benes.scala 90:27]
  wire [15:0] in_switch_19_io_z; // @[Benes.scala 90:27]
  wire [15:0] in_switch_19_io_in; // @[Benes.scala 90:27]
  wire [15:0] in_switch_20_io_y; // @[Benes.scala 90:27]
  wire [15:0] in_switch_20_io_z; // @[Benes.scala 90:27]
  wire [15:0] in_switch_20_io_in; // @[Benes.scala 90:27]
  wire [15:0] in_switch_21_io_y; // @[Benes.scala 90:27]
  wire [15:0] in_switch_21_io_z; // @[Benes.scala 90:27]
  wire [15:0] in_switch_21_io_in; // @[Benes.scala 90:27]
  wire [15:0] in_switch_22_io_y; // @[Benes.scala 90:27]
  wire [15:0] in_switch_22_io_z; // @[Benes.scala 90:27]
  wire [15:0] in_switch_22_io_in; // @[Benes.scala 90:27]
  wire [15:0] in_switch_23_io_y; // @[Benes.scala 90:27]
  wire [15:0] in_switch_23_io_z; // @[Benes.scala 90:27]
  wire [15:0] in_switch_23_io_in; // @[Benes.scala 90:27]
  wire [15:0] in_switch_24_io_y; // @[Benes.scala 90:27]
  wire [15:0] in_switch_24_io_z; // @[Benes.scala 90:27]
  wire [15:0] in_switch_24_io_in; // @[Benes.scala 90:27]
  wire [15:0] in_switch_25_io_y; // @[Benes.scala 90:27]
  wire [15:0] in_switch_25_io_z; // @[Benes.scala 90:27]
  wire [15:0] in_switch_25_io_in; // @[Benes.scala 90:27]
  wire [15:0] in_switch_26_io_y; // @[Benes.scala 90:27]
  wire [15:0] in_switch_26_io_z; // @[Benes.scala 90:27]
  wire [15:0] in_switch_26_io_in; // @[Benes.scala 90:27]
  wire [15:0] in_switch_27_io_y; // @[Benes.scala 90:27]
  wire [15:0] in_switch_27_io_z; // @[Benes.scala 90:27]
  wire [15:0] in_switch_27_io_in; // @[Benes.scala 90:27]
  wire [15:0] in_switch_28_io_y; // @[Benes.scala 90:27]
  wire [15:0] in_switch_28_io_z; // @[Benes.scala 90:27]
  wire [15:0] in_switch_28_io_in; // @[Benes.scala 90:27]
  wire [15:0] in_switch_29_io_y; // @[Benes.scala 90:27]
  wire [15:0] in_switch_29_io_z; // @[Benes.scala 90:27]
  wire [15:0] in_switch_29_io_in; // @[Benes.scala 90:27]
  wire [15:0] in_switch_30_io_y; // @[Benes.scala 90:27]
  wire [15:0] in_switch_30_io_z; // @[Benes.scala 90:27]
  wire [15:0] in_switch_30_io_in; // @[Benes.scala 90:27]
  wire [15:0] in_switch_31_io_y; // @[Benes.scala 90:27]
  wire [15:0] in_switch_31_io_z; // @[Benes.scala 90:27]
  wire [15:0] in_switch_31_io_in; // @[Benes.scala 90:27]
  wire [15:0] out_switch_io_y; // @[Benes.scala 99:28]
  wire [15:0] out_switch_io_in0; // @[Benes.scala 99:28]
  wire [15:0] out_switch_1_io_y; // @[Benes.scala 99:28]
  wire [15:0] out_switch_1_io_in0; // @[Benes.scala 99:28]
  wire [15:0] out_switch_2_io_y; // @[Benes.scala 99:28]
  wire [15:0] out_switch_2_io_in0; // @[Benes.scala 99:28]
  wire [15:0] out_switch_3_io_y; // @[Benes.scala 99:28]
  wire [15:0] out_switch_3_io_in0; // @[Benes.scala 99:28]
  wire [15:0] out_switch_4_io_y; // @[Benes.scala 99:28]
  wire [15:0] out_switch_4_io_in0; // @[Benes.scala 99:28]
  wire [15:0] out_switch_5_io_y; // @[Benes.scala 99:28]
  wire [15:0] out_switch_5_io_in0; // @[Benes.scala 99:28]
  wire [15:0] out_switch_6_io_y; // @[Benes.scala 99:28]
  wire [15:0] out_switch_6_io_in0; // @[Benes.scala 99:28]
  wire [15:0] out_switch_7_io_y; // @[Benes.scala 99:28]
  wire [15:0] out_switch_7_io_in0; // @[Benes.scala 99:28]
  wire [15:0] out_switch_8_io_y; // @[Benes.scala 99:28]
  wire [15:0] out_switch_8_io_in0; // @[Benes.scala 99:28]
  wire [15:0] out_switch_9_io_y; // @[Benes.scala 99:28]
  wire [15:0] out_switch_9_io_in0; // @[Benes.scala 99:28]
  wire [15:0] out_switch_10_io_y; // @[Benes.scala 99:28]
  wire [15:0] out_switch_10_io_in0; // @[Benes.scala 99:28]
  wire [15:0] out_switch_11_io_y; // @[Benes.scala 99:28]
  wire [15:0] out_switch_11_io_in0; // @[Benes.scala 99:28]
  wire [15:0] out_switch_12_io_y; // @[Benes.scala 99:28]
  wire [15:0] out_switch_12_io_in0; // @[Benes.scala 99:28]
  wire [15:0] out_switch_13_io_y; // @[Benes.scala 99:28]
  wire [15:0] out_switch_13_io_in0; // @[Benes.scala 99:28]
  wire [15:0] out_switch_14_io_y; // @[Benes.scala 99:28]
  wire [15:0] out_switch_14_io_in0; // @[Benes.scala 99:28]
  wire [15:0] out_switch_15_io_y; // @[Benes.scala 99:28]
  wire [15:0] out_switch_15_io_in0; // @[Benes.scala 99:28]
  wire [15:0] out_switch_16_io_y; // @[Benes.scala 99:28]
  wire [15:0] out_switch_16_io_in0; // @[Benes.scala 99:28]
  wire [15:0] out_switch_17_io_y; // @[Benes.scala 99:28]
  wire [15:0] out_switch_17_io_in0; // @[Benes.scala 99:28]
  wire [15:0] out_switch_18_io_y; // @[Benes.scala 99:28]
  wire [15:0] out_switch_18_io_in0; // @[Benes.scala 99:28]
  wire [15:0] out_switch_19_io_y; // @[Benes.scala 99:28]
  wire [15:0] out_switch_19_io_in0; // @[Benes.scala 99:28]
  wire [15:0] out_switch_20_io_y; // @[Benes.scala 99:28]
  wire [15:0] out_switch_20_io_in0; // @[Benes.scala 99:28]
  wire [15:0] out_switch_21_io_y; // @[Benes.scala 99:28]
  wire [15:0] out_switch_21_io_in0; // @[Benes.scala 99:28]
  wire [15:0] out_switch_22_io_y; // @[Benes.scala 99:28]
  wire [15:0] out_switch_22_io_in0; // @[Benes.scala 99:28]
  wire [15:0] out_switch_23_io_y; // @[Benes.scala 99:28]
  wire [15:0] out_switch_23_io_in0; // @[Benes.scala 99:28]
  wire [15:0] out_switch_24_io_y; // @[Benes.scala 99:28]
  wire [15:0] out_switch_24_io_in0; // @[Benes.scala 99:28]
  wire [15:0] out_switch_25_io_y; // @[Benes.scala 99:28]
  wire [15:0] out_switch_25_io_in0; // @[Benes.scala 99:28]
  wire [15:0] out_switch_26_io_y; // @[Benes.scala 99:28]
  wire [15:0] out_switch_26_io_in0; // @[Benes.scala 99:28]
  wire [15:0] out_switch_27_io_y; // @[Benes.scala 99:28]
  wire [15:0] out_switch_27_io_in0; // @[Benes.scala 99:28]
  wire [15:0] out_switch_28_io_y; // @[Benes.scala 99:28]
  wire [15:0] out_switch_28_io_in0; // @[Benes.scala 99:28]
  wire [15:0] out_switch_29_io_y; // @[Benes.scala 99:28]
  wire [15:0] out_switch_29_io_in0; // @[Benes.scala 99:28]
  wire [15:0] out_switch_30_io_y; // @[Benes.scala 99:28]
  wire [15:0] out_switch_30_io_in0; // @[Benes.scala 99:28]
  wire [15:0] out_switch_31_io_y; // @[Benes.scala 99:28]
  wire [15:0] out_switch_31_io_in0; // @[Benes.scala 99:28]
  wire [15:0] imm_switch_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_1_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_1_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_1_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_2_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_2_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_2_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_3_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_3_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_3_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_4_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_4_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_4_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_5_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_5_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_5_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_6_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_6_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_6_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_7_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_7_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_7_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_8_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_8_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_8_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_9_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_9_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_9_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_10_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_10_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_10_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_11_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_11_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_11_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_12_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_12_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_12_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_13_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_13_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_13_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_14_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_14_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_14_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_15_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_15_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_15_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_16_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_16_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_16_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_17_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_17_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_17_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_18_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_18_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_18_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_19_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_19_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_19_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_20_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_20_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_20_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_21_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_21_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_21_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_22_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_22_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_22_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_23_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_23_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_23_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_24_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_24_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_24_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_25_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_25_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_25_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_26_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_26_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_26_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_27_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_27_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_27_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_28_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_28_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_28_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_29_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_29_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_29_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_30_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_30_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_30_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_31_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_31_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_31_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_32_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_32_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_32_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_33_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_33_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_33_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_34_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_34_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_34_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_35_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_35_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_35_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_36_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_36_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_36_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_37_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_37_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_37_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_38_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_38_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_38_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_39_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_39_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_39_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_40_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_40_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_40_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_41_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_41_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_41_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_42_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_42_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_42_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_43_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_43_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_43_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_44_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_44_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_44_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_45_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_45_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_45_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_46_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_46_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_46_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_47_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_47_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_47_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_48_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_48_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_48_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_49_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_49_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_49_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_50_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_50_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_50_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_51_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_51_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_51_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_52_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_52_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_52_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_53_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_53_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_53_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_54_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_54_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_54_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_55_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_55_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_55_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_56_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_56_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_56_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_57_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_57_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_57_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_58_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_58_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_58_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_59_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_59_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_59_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_60_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_60_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_60_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_61_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_61_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_61_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_62_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_62_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_62_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_63_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_63_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_63_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_64_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_64_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_64_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_65_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_65_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_65_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_66_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_66_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_66_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_67_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_67_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_67_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_68_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_68_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_68_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_69_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_69_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_69_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_70_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_70_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_70_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_71_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_71_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_71_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_72_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_72_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_72_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_73_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_73_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_73_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_74_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_74_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_74_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_75_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_75_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_75_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_76_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_76_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_76_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_77_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_77_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_77_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_78_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_78_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_78_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_79_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_79_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_79_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_80_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_80_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_80_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_81_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_81_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_81_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_82_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_82_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_82_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_83_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_83_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_83_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_84_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_84_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_84_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_85_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_85_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_85_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_86_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_86_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_86_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_87_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_87_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_87_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_88_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_88_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_88_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_89_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_89_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_89_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_90_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_90_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_90_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_91_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_91_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_91_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_92_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_92_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_92_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_93_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_93_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_93_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_94_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_94_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_94_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_95_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_95_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_95_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_96_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_96_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_96_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_97_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_97_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_97_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_98_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_98_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_98_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_99_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_99_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_99_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_100_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_100_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_100_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_101_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_101_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_101_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_102_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_102_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_102_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_103_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_103_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_103_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_104_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_104_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_104_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_105_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_105_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_105_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_106_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_106_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_106_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_107_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_107_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_107_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_108_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_108_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_108_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_109_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_109_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_109_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_110_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_110_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_110_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_111_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_111_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_111_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_112_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_112_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_112_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_113_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_113_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_113_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_114_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_114_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_114_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_115_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_115_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_115_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_116_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_116_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_116_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_117_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_117_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_117_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_118_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_118_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_118_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_119_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_119_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_119_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_120_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_120_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_120_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_121_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_121_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_121_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_122_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_122_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_122_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_123_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_123_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_123_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_124_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_124_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_124_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_125_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_125_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_125_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_126_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_126_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_126_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_127_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_127_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_127_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_128_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_128_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_128_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_129_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_129_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_129_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_130_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_130_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_130_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_131_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_131_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_131_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_132_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_132_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_132_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_133_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_133_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_133_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_134_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_134_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_134_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_135_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_135_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_135_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_136_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_136_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_136_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_137_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_137_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_137_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_138_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_138_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_138_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_139_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_139_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_139_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_140_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_140_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_140_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_141_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_141_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_141_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_142_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_142_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_142_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_143_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_143_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_143_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_144_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_144_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_144_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_145_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_145_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_145_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_146_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_146_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_146_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_147_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_147_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_147_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_148_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_148_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_148_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_149_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_149_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_149_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_150_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_150_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_150_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_151_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_151_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_151_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_152_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_152_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_152_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_153_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_153_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_153_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_154_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_154_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_154_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_155_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_155_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_155_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_156_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_156_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_156_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_157_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_157_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_157_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_158_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_158_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_158_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_159_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_159_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_159_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_160_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_160_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_160_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_161_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_161_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_161_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_162_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_162_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_162_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_163_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_163_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_163_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_164_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_164_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_164_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_165_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_165_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_165_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_166_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_166_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_166_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_167_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_167_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_167_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_168_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_168_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_168_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_169_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_169_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_169_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_170_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_170_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_170_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_171_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_171_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_171_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_172_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_172_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_172_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_173_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_173_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_173_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_174_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_174_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_174_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_175_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_175_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_175_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_176_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_176_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_176_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_177_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_177_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_177_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_178_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_178_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_178_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_179_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_179_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_179_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_180_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_180_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_180_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_181_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_181_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_181_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_182_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_182_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_182_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_183_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_183_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_183_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_184_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_184_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_184_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_185_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_185_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_185_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_186_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_186_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_186_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_187_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_187_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_187_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_188_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_188_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_188_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_189_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_189_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_189_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_190_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_190_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_190_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_191_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_191_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_191_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_192_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_192_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_192_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_193_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_193_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_193_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_194_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_194_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_194_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_195_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_195_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_195_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_196_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_196_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_196_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_197_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_197_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_197_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_198_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_198_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_198_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_199_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_199_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_199_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_200_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_200_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_200_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_201_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_201_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_201_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_202_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_202_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_202_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_203_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_203_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_203_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_204_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_204_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_204_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_205_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_205_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_205_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_206_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_206_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_206_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_207_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_207_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_207_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_208_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_208_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_208_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_209_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_209_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_209_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_210_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_210_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_210_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_211_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_211_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_211_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_212_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_212_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_212_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_213_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_213_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_213_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_214_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_214_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_214_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_215_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_215_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_215_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_216_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_216_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_216_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_217_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_217_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_217_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_218_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_218_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_218_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_219_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_219_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_219_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_220_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_220_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_220_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_221_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_221_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_221_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_222_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_222_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_222_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_223_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_223_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_223_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_224_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_224_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_224_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_225_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_225_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_225_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_226_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_226_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_226_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_227_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_227_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_227_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_228_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_228_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_228_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_229_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_229_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_229_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_230_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_230_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_230_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_231_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_231_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_231_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_232_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_232_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_232_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_233_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_233_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_233_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_234_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_234_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_234_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_235_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_235_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_235_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_236_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_236_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_236_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_237_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_237_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_237_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_238_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_238_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_238_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_239_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_239_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_239_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_240_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_240_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_240_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_241_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_241_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_241_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_242_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_242_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_242_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_243_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_243_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_243_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_244_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_244_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_244_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_245_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_245_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_245_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_246_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_246_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_246_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_247_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_247_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_247_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_248_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_248_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_248_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_249_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_249_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_249_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_250_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_250_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_250_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_251_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_251_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_251_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_252_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_252_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_252_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_253_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_253_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_253_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_254_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_254_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_254_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_255_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_255_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_255_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_256_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_256_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_256_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_257_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_257_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_257_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_258_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_258_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_258_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_259_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_259_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_259_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_260_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_260_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_260_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_261_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_261_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_261_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_262_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_262_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_262_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_263_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_263_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_263_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_264_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_264_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_264_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_265_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_265_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_265_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_266_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_266_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_266_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_267_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_267_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_267_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_268_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_268_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_268_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_269_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_269_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_269_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_270_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_270_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_270_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_271_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_271_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_271_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_272_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_272_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_272_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_273_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_273_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_273_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_274_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_274_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_274_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_275_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_275_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_275_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_276_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_276_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_276_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_277_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_277_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_277_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_278_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_278_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_278_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_279_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_279_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_279_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_280_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_280_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_280_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_281_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_281_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_281_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_282_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_282_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_282_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_283_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_283_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_283_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_284_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_284_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_284_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_285_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_285_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_285_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_286_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_286_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_286_io_in0; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_287_io_y; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_287_io_z; // @[Benes.scala 109:30]
  wire [15:0] imm_switch_287_io_in0; // @[Benes.scala 109:30]
  reg [15:0] r_data_bus_ff_0; // @[Benes.scala 77:32]
  reg [15:0] r_data_bus_ff_1; // @[Benes.scala 77:32]
  reg [15:0] r_data_bus_ff_2; // @[Benes.scala 77:32]
  reg [15:0] r_data_bus_ff_3; // @[Benes.scala 77:32]
  reg [15:0] r_data_bus_ff_4; // @[Benes.scala 77:32]
  reg [15:0] r_data_bus_ff_5; // @[Benes.scala 77:32]
  reg [15:0] r_data_bus_ff_6; // @[Benes.scala 77:32]
  reg [15:0] r_data_bus_ff_7; // @[Benes.scala 77:32]
  reg [15:0] r_data_bus_ff_8; // @[Benes.scala 77:32]
  reg [15:0] r_data_bus_ff_9; // @[Benes.scala 77:32]
  reg [15:0] r_data_bus_ff_10; // @[Benes.scala 77:32]
  reg [15:0] r_data_bus_ff_11; // @[Benes.scala 77:32]
  reg [15:0] r_data_bus_ff_12; // @[Benes.scala 77:32]
  reg [15:0] r_data_bus_ff_13; // @[Benes.scala 77:32]
  reg [15:0] r_data_bus_ff_14; // @[Benes.scala 77:32]
  reg [15:0] r_data_bus_ff_15; // @[Benes.scala 77:32]
  reg [15:0] r_data_bus_ff_16; // @[Benes.scala 77:32]
  reg [15:0] r_data_bus_ff_17; // @[Benes.scala 77:32]
  reg [15:0] r_data_bus_ff_18; // @[Benes.scala 77:32]
  reg [15:0] r_data_bus_ff_19; // @[Benes.scala 77:32]
  reg [15:0] r_data_bus_ff_20; // @[Benes.scala 77:32]
  reg [15:0] r_data_bus_ff_21; // @[Benes.scala 77:32]
  reg [15:0] r_data_bus_ff_22; // @[Benes.scala 77:32]
  reg [15:0] r_data_bus_ff_23; // @[Benes.scala 77:32]
  reg [15:0] r_data_bus_ff_24; // @[Benes.scala 77:32]
  reg [15:0] r_data_bus_ff_25; // @[Benes.scala 77:32]
  reg [15:0] r_data_bus_ff_26; // @[Benes.scala 77:32]
  reg [15:0] r_data_bus_ff_27; // @[Benes.scala 77:32]
  reg [15:0] r_data_bus_ff_28; // @[Benes.scala 77:32]
  reg [15:0] r_data_bus_ff_29; // @[Benes.scala 77:32]
  reg [15:0] r_data_bus_ff_30; // @[Benes.scala 77:32]
  reg [15:0] r_data_bus_ff_31; // @[Benes.scala 77:32]
  wire [15:0] w_dist_bus_0 = out_switch_io_y; // @[Benes.scala 103:23 79:29]
  wire [15:0] w_dist_bus_1 = out_switch_1_io_y; // @[Benes.scala 103:23 79:29]
  wire [15:0] w_dist_bus_2 = out_switch_2_io_y; // @[Benes.scala 103:23 79:29]
  wire [15:0] w_dist_bus_3 = out_switch_3_io_y; // @[Benes.scala 103:23 79:29]
  wire [15:0] w_dist_bus_4 = out_switch_4_io_y; // @[Benes.scala 103:23 79:29]
  wire [15:0] w_dist_bus_5 = out_switch_5_io_y; // @[Benes.scala 103:23 79:29]
  wire [15:0] w_dist_bus_6 = out_switch_6_io_y; // @[Benes.scala 103:23 79:29]
  wire [15:0] w_dist_bus_7 = out_switch_7_io_y; // @[Benes.scala 103:23 79:29]
  wire [15:0] w_dist_bus_8 = out_switch_8_io_y; // @[Benes.scala 103:23 79:29]
  wire [15:0] w_dist_bus_9 = out_switch_9_io_y; // @[Benes.scala 103:23 79:29]
  wire [15:0] w_dist_bus_10 = out_switch_10_io_y; // @[Benes.scala 103:23 79:29]
  wire [15:0] w_dist_bus_11 = out_switch_11_io_y; // @[Benes.scala 103:23 79:29]
  wire [15:0] w_dist_bus_12 = out_switch_12_io_y; // @[Benes.scala 103:23 79:29]
  wire [15:0] w_dist_bus_13 = out_switch_13_io_y; // @[Benes.scala 103:23 79:29]
  wire [15:0] w_dist_bus_14 = out_switch_14_io_y; // @[Benes.scala 103:23 79:29]
  wire [15:0] w_dist_bus_15 = out_switch_15_io_y; // @[Benes.scala 103:23 79:29]
  wire [15:0] w_dist_bus_16 = out_switch_16_io_y; // @[Benes.scala 103:23 79:29]
  wire [15:0] w_dist_bus_17 = out_switch_17_io_y; // @[Benes.scala 103:23 79:29]
  wire [15:0] w_dist_bus_18 = out_switch_18_io_y; // @[Benes.scala 103:23 79:29]
  wire [15:0] w_dist_bus_19 = out_switch_19_io_y; // @[Benes.scala 103:23 79:29]
  wire [15:0] w_dist_bus_20 = out_switch_20_io_y; // @[Benes.scala 103:23 79:29]
  wire [15:0] w_dist_bus_21 = out_switch_21_io_y; // @[Benes.scala 103:23 79:29]
  wire [15:0] w_dist_bus_22 = out_switch_22_io_y; // @[Benes.scala 103:23 79:29]
  wire [15:0] w_dist_bus_23 = out_switch_23_io_y; // @[Benes.scala 103:23 79:29]
  wire [15:0] w_dist_bus_24 = out_switch_24_io_y; // @[Benes.scala 103:23 79:29]
  wire [15:0] w_dist_bus_25 = out_switch_25_io_y; // @[Benes.scala 103:23 79:29]
  wire [15:0] w_dist_bus_26 = out_switch_26_io_y; // @[Benes.scala 103:23 79:29]
  wire [15:0] w_dist_bus_27 = out_switch_27_io_y; // @[Benes.scala 103:23 79:29]
  wire [15:0] w_dist_bus_28 = out_switch_28_io_y; // @[Benes.scala 103:23 79:29]
  wire [15:0] w_dist_bus_29 = out_switch_29_io_y; // @[Benes.scala 103:23 79:29]
  wire [15:0] w_dist_bus_30 = out_switch_30_io_y; // @[Benes.scala 103:23 79:29]
  wire [15:0] w_dist_bus_31 = out_switch_31_io_y; // @[Benes.scala 103:23 79:29]
  wire [15:0] w_internal_0 = in_switch_io_y; // @[Benes.scala 80:29 92:43]
  wire [15:0] w_internal_1 = in_switch_io_z; // @[Benes.scala 80:29 93:43]
  wire [15:0] w_internal_2 = imm_switch_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_3 = imm_switch_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_4 = imm_switch_1_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_5 = imm_switch_1_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_6 = imm_switch_2_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_7 = imm_switch_2_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_8 = imm_switch_3_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_9 = imm_switch_3_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_10 = imm_switch_4_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_11 = imm_switch_4_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_12 = imm_switch_5_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_13 = imm_switch_5_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_14 = imm_switch_6_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_15 = imm_switch_6_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_16 = imm_switch_7_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_17 = imm_switch_7_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_18 = imm_switch_8_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_19 = imm_switch_8_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_20 = in_switch_1_io_y; // @[Benes.scala 80:29 92:43]
  wire [15:0] w_internal_21 = in_switch_1_io_z; // @[Benes.scala 80:29 93:43]
  wire [15:0] w_internal_22 = imm_switch_9_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_23 = imm_switch_9_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_24 = imm_switch_10_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_25 = imm_switch_10_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_26 = imm_switch_11_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_27 = imm_switch_11_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_28 = imm_switch_12_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_29 = imm_switch_12_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_30 = imm_switch_13_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_31 = imm_switch_13_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_32 = imm_switch_14_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_33 = imm_switch_14_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_34 = imm_switch_15_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_35 = imm_switch_15_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_36 = imm_switch_16_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_37 = imm_switch_16_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_38 = imm_switch_17_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_39 = imm_switch_17_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_40 = in_switch_2_io_y; // @[Benes.scala 80:29 92:43]
  wire [15:0] w_internal_41 = in_switch_2_io_z; // @[Benes.scala 80:29 93:43]
  wire [15:0] w_internal_42 = imm_switch_18_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_43 = imm_switch_18_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_44 = imm_switch_19_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_45 = imm_switch_19_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_46 = imm_switch_20_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_47 = imm_switch_20_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_48 = imm_switch_21_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_49 = imm_switch_21_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_50 = imm_switch_22_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_51 = imm_switch_22_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_52 = imm_switch_23_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_53 = imm_switch_23_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_54 = imm_switch_24_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_55 = imm_switch_24_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_56 = imm_switch_25_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_57 = imm_switch_25_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_58 = imm_switch_26_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_59 = imm_switch_26_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_60 = in_switch_3_io_y; // @[Benes.scala 80:29 92:43]
  wire [15:0] w_internal_61 = in_switch_3_io_z; // @[Benes.scala 80:29 93:43]
  wire [15:0] w_internal_62 = imm_switch_27_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_63 = imm_switch_27_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_64 = imm_switch_28_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_65 = imm_switch_28_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_66 = imm_switch_29_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_67 = imm_switch_29_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_68 = imm_switch_30_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_69 = imm_switch_30_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_70 = imm_switch_31_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_71 = imm_switch_31_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_72 = imm_switch_32_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_73 = imm_switch_32_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_74 = imm_switch_33_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_75 = imm_switch_33_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_76 = imm_switch_34_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_77 = imm_switch_34_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_78 = imm_switch_35_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_79 = imm_switch_35_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_80 = in_switch_4_io_y; // @[Benes.scala 80:29 92:43]
  wire [15:0] w_internal_81 = in_switch_4_io_z; // @[Benes.scala 80:29 93:43]
  wire [15:0] w_internal_82 = imm_switch_36_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_83 = imm_switch_36_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_84 = imm_switch_37_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_85 = imm_switch_37_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_86 = imm_switch_38_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_87 = imm_switch_38_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_88 = imm_switch_39_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_89 = imm_switch_39_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_90 = imm_switch_40_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_91 = imm_switch_40_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_92 = imm_switch_41_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_93 = imm_switch_41_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_94 = imm_switch_42_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_95 = imm_switch_42_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_96 = imm_switch_43_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_97 = imm_switch_43_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_98 = imm_switch_44_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_99 = imm_switch_44_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_100 = in_switch_5_io_y; // @[Benes.scala 80:29 92:43]
  wire [15:0] w_internal_101 = in_switch_5_io_z; // @[Benes.scala 80:29 93:43]
  wire [15:0] w_internal_102 = imm_switch_45_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_103 = imm_switch_45_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_104 = imm_switch_46_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_105 = imm_switch_46_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_106 = imm_switch_47_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_107 = imm_switch_47_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_108 = imm_switch_48_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_109 = imm_switch_48_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_110 = imm_switch_49_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_111 = imm_switch_49_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_112 = imm_switch_50_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_113 = imm_switch_50_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_114 = imm_switch_51_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_115 = imm_switch_51_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_116 = imm_switch_52_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_117 = imm_switch_52_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_118 = imm_switch_53_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_119 = imm_switch_53_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_120 = in_switch_6_io_y; // @[Benes.scala 80:29 92:43]
  wire [15:0] w_internal_121 = in_switch_6_io_z; // @[Benes.scala 80:29 93:43]
  wire [15:0] w_internal_122 = imm_switch_54_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_123 = imm_switch_54_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_124 = imm_switch_55_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_125 = imm_switch_55_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_126 = imm_switch_56_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_127 = imm_switch_56_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_128 = imm_switch_57_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_129 = imm_switch_57_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_130 = imm_switch_58_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_131 = imm_switch_58_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_132 = imm_switch_59_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_133 = imm_switch_59_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_134 = imm_switch_60_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_135 = imm_switch_60_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_136 = imm_switch_61_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_137 = imm_switch_61_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_138 = imm_switch_62_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_139 = imm_switch_62_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_140 = in_switch_7_io_y; // @[Benes.scala 80:29 92:43]
  wire [15:0] w_internal_141 = in_switch_7_io_z; // @[Benes.scala 80:29 93:43]
  wire [15:0] w_internal_142 = imm_switch_63_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_143 = imm_switch_63_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_144 = imm_switch_64_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_145 = imm_switch_64_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_146 = imm_switch_65_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_147 = imm_switch_65_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_148 = imm_switch_66_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_149 = imm_switch_66_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_150 = imm_switch_67_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_151 = imm_switch_67_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_152 = imm_switch_68_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_153 = imm_switch_68_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_154 = imm_switch_69_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_155 = imm_switch_69_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_156 = imm_switch_70_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_157 = imm_switch_70_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_158 = imm_switch_71_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_159 = imm_switch_71_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_160 = in_switch_8_io_y; // @[Benes.scala 80:29 92:43]
  wire [15:0] w_internal_161 = in_switch_8_io_z; // @[Benes.scala 80:29 93:43]
  wire [15:0] w_internal_162 = imm_switch_72_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_163 = imm_switch_72_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_164 = imm_switch_73_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_165 = imm_switch_73_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_166 = imm_switch_74_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_167 = imm_switch_74_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_168 = imm_switch_75_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_169 = imm_switch_75_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_170 = imm_switch_76_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_171 = imm_switch_76_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_172 = imm_switch_77_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_173 = imm_switch_77_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_174 = imm_switch_78_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_175 = imm_switch_78_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_176 = imm_switch_79_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_177 = imm_switch_79_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_178 = imm_switch_80_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_179 = imm_switch_80_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_180 = in_switch_9_io_y; // @[Benes.scala 80:29 92:43]
  wire [15:0] w_internal_181 = in_switch_9_io_z; // @[Benes.scala 80:29 93:43]
  wire [15:0] w_internal_182 = imm_switch_81_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_183 = imm_switch_81_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_184 = imm_switch_82_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_185 = imm_switch_82_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_186 = imm_switch_83_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_187 = imm_switch_83_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_188 = imm_switch_84_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_189 = imm_switch_84_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_190 = imm_switch_85_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_191 = imm_switch_85_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_192 = imm_switch_86_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_193 = imm_switch_86_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_194 = imm_switch_87_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_195 = imm_switch_87_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_196 = imm_switch_88_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_197 = imm_switch_88_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_198 = imm_switch_89_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_199 = imm_switch_89_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_200 = in_switch_10_io_y; // @[Benes.scala 80:29 92:43]
  wire [15:0] w_internal_201 = in_switch_10_io_z; // @[Benes.scala 80:29 93:43]
  wire [15:0] w_internal_202 = imm_switch_90_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_203 = imm_switch_90_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_204 = imm_switch_91_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_205 = imm_switch_91_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_206 = imm_switch_92_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_207 = imm_switch_92_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_208 = imm_switch_93_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_209 = imm_switch_93_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_210 = imm_switch_94_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_211 = imm_switch_94_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_212 = imm_switch_95_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_213 = imm_switch_95_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_214 = imm_switch_96_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_215 = imm_switch_96_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_216 = imm_switch_97_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_217 = imm_switch_97_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_218 = imm_switch_98_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_219 = imm_switch_98_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_220 = in_switch_11_io_y; // @[Benes.scala 80:29 92:43]
  wire [15:0] w_internal_221 = in_switch_11_io_z; // @[Benes.scala 80:29 93:43]
  wire [15:0] w_internal_222 = imm_switch_99_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_223 = imm_switch_99_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_224 = imm_switch_100_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_225 = imm_switch_100_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_226 = imm_switch_101_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_227 = imm_switch_101_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_228 = imm_switch_102_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_229 = imm_switch_102_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_230 = imm_switch_103_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_231 = imm_switch_103_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_232 = imm_switch_104_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_233 = imm_switch_104_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_234 = imm_switch_105_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_235 = imm_switch_105_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_236 = imm_switch_106_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_237 = imm_switch_106_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_238 = imm_switch_107_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_239 = imm_switch_107_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_240 = in_switch_12_io_y; // @[Benes.scala 80:29 92:43]
  wire [15:0] w_internal_241 = in_switch_12_io_z; // @[Benes.scala 80:29 93:43]
  wire [15:0] w_internal_242 = imm_switch_108_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_243 = imm_switch_108_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_244 = imm_switch_109_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_245 = imm_switch_109_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_246 = imm_switch_110_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_247 = imm_switch_110_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_248 = imm_switch_111_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_249 = imm_switch_111_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_250 = imm_switch_112_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_251 = imm_switch_112_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_252 = imm_switch_113_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_253 = imm_switch_113_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_254 = imm_switch_114_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_255 = imm_switch_114_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_256 = imm_switch_115_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_257 = imm_switch_115_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_258 = imm_switch_116_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_259 = imm_switch_116_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_260 = in_switch_13_io_y; // @[Benes.scala 80:29 92:43]
  wire [15:0] w_internal_261 = in_switch_13_io_z; // @[Benes.scala 80:29 93:43]
  wire [15:0] w_internal_262 = imm_switch_117_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_263 = imm_switch_117_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_264 = imm_switch_118_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_265 = imm_switch_118_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_266 = imm_switch_119_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_267 = imm_switch_119_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_268 = imm_switch_120_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_269 = imm_switch_120_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_270 = imm_switch_121_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_271 = imm_switch_121_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_272 = imm_switch_122_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_273 = imm_switch_122_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_274 = imm_switch_123_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_275 = imm_switch_123_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_276 = imm_switch_124_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_277 = imm_switch_124_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_278 = imm_switch_125_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_279 = imm_switch_125_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_280 = in_switch_14_io_y; // @[Benes.scala 80:29 92:43]
  wire [15:0] w_internal_281 = in_switch_14_io_z; // @[Benes.scala 80:29 93:43]
  wire [15:0] w_internal_282 = imm_switch_126_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_283 = imm_switch_126_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_284 = imm_switch_127_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_285 = imm_switch_127_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_286 = imm_switch_128_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_287 = imm_switch_128_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_288 = imm_switch_129_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_289 = imm_switch_129_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_290 = imm_switch_130_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_291 = imm_switch_130_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_292 = imm_switch_131_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_293 = imm_switch_131_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_294 = imm_switch_132_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_295 = imm_switch_132_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_296 = imm_switch_133_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_297 = imm_switch_133_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_298 = imm_switch_134_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_299 = imm_switch_134_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_300 = in_switch_15_io_y; // @[Benes.scala 80:29 92:43]
  wire [15:0] w_internal_301 = in_switch_15_io_z; // @[Benes.scala 80:29 93:43]
  wire [15:0] w_internal_302 = imm_switch_135_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_303 = imm_switch_135_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_304 = imm_switch_136_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_305 = imm_switch_136_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_306 = imm_switch_137_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_307 = imm_switch_137_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_308 = imm_switch_138_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_309 = imm_switch_138_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_310 = imm_switch_139_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_311 = imm_switch_139_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_312 = imm_switch_140_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_313 = imm_switch_140_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_314 = imm_switch_141_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_315 = imm_switch_141_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_316 = imm_switch_142_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_317 = imm_switch_142_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_318 = imm_switch_143_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_319 = imm_switch_143_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_320 = in_switch_16_io_y; // @[Benes.scala 80:29 92:43]
  wire [15:0] w_internal_321 = in_switch_16_io_z; // @[Benes.scala 80:29 93:43]
  wire [15:0] w_internal_322 = imm_switch_144_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_323 = imm_switch_144_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_324 = imm_switch_145_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_325 = imm_switch_145_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_326 = imm_switch_146_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_327 = imm_switch_146_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_328 = imm_switch_147_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_329 = imm_switch_147_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_330 = imm_switch_148_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_331 = imm_switch_148_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_332 = imm_switch_149_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_333 = imm_switch_149_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_334 = imm_switch_150_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_335 = imm_switch_150_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_336 = imm_switch_151_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_337 = imm_switch_151_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_338 = imm_switch_152_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_339 = imm_switch_152_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_340 = in_switch_17_io_y; // @[Benes.scala 80:29 92:43]
  wire [15:0] w_internal_341 = in_switch_17_io_z; // @[Benes.scala 80:29 93:43]
  wire [15:0] w_internal_342 = imm_switch_153_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_343 = imm_switch_153_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_344 = imm_switch_154_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_345 = imm_switch_154_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_346 = imm_switch_155_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_347 = imm_switch_155_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_348 = imm_switch_156_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_349 = imm_switch_156_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_350 = imm_switch_157_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_351 = imm_switch_157_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_352 = imm_switch_158_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_353 = imm_switch_158_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_354 = imm_switch_159_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_355 = imm_switch_159_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_356 = imm_switch_160_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_357 = imm_switch_160_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_358 = imm_switch_161_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_359 = imm_switch_161_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_360 = in_switch_18_io_y; // @[Benes.scala 80:29 92:43]
  wire [15:0] w_internal_361 = in_switch_18_io_z; // @[Benes.scala 80:29 93:43]
  wire [15:0] w_internal_362 = imm_switch_162_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_363 = imm_switch_162_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_364 = imm_switch_163_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_365 = imm_switch_163_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_366 = imm_switch_164_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_367 = imm_switch_164_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_368 = imm_switch_165_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_369 = imm_switch_165_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_370 = imm_switch_166_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_371 = imm_switch_166_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_372 = imm_switch_167_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_373 = imm_switch_167_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_374 = imm_switch_168_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_375 = imm_switch_168_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_376 = imm_switch_169_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_377 = imm_switch_169_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_378 = imm_switch_170_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_379 = imm_switch_170_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_380 = in_switch_19_io_y; // @[Benes.scala 80:29 92:43]
  wire [15:0] w_internal_381 = in_switch_19_io_z; // @[Benes.scala 80:29 93:43]
  wire [15:0] w_internal_382 = imm_switch_171_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_383 = imm_switch_171_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_384 = imm_switch_172_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_385 = imm_switch_172_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_386 = imm_switch_173_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_387 = imm_switch_173_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_388 = imm_switch_174_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_389 = imm_switch_174_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_390 = imm_switch_175_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_391 = imm_switch_175_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_392 = imm_switch_176_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_393 = imm_switch_176_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_394 = imm_switch_177_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_395 = imm_switch_177_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_396 = imm_switch_178_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_397 = imm_switch_178_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_398 = imm_switch_179_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_399 = imm_switch_179_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_400 = in_switch_20_io_y; // @[Benes.scala 80:29 92:43]
  wire [15:0] w_internal_401 = in_switch_20_io_z; // @[Benes.scala 80:29 93:43]
  wire [15:0] w_internal_402 = imm_switch_180_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_403 = imm_switch_180_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_404 = imm_switch_181_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_405 = imm_switch_181_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_406 = imm_switch_182_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_407 = imm_switch_182_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_408 = imm_switch_183_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_409 = imm_switch_183_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_410 = imm_switch_184_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_411 = imm_switch_184_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_412 = imm_switch_185_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_413 = imm_switch_185_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_414 = imm_switch_186_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_415 = imm_switch_186_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_416 = imm_switch_187_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_417 = imm_switch_187_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_418 = imm_switch_188_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_419 = imm_switch_188_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_420 = in_switch_21_io_y; // @[Benes.scala 80:29 92:43]
  wire [15:0] w_internal_421 = in_switch_21_io_z; // @[Benes.scala 80:29 93:43]
  wire [15:0] w_internal_422 = imm_switch_189_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_423 = imm_switch_189_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_424 = imm_switch_190_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_425 = imm_switch_190_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_426 = imm_switch_191_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_427 = imm_switch_191_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_428 = imm_switch_192_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_429 = imm_switch_192_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_430 = imm_switch_193_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_431 = imm_switch_193_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_432 = imm_switch_194_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_433 = imm_switch_194_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_434 = imm_switch_195_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_435 = imm_switch_195_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_436 = imm_switch_196_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_437 = imm_switch_196_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_438 = imm_switch_197_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_439 = imm_switch_197_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_440 = in_switch_22_io_y; // @[Benes.scala 80:29 92:43]
  wire [15:0] w_internal_441 = in_switch_22_io_z; // @[Benes.scala 80:29 93:43]
  wire [15:0] w_internal_442 = imm_switch_198_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_443 = imm_switch_198_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_444 = imm_switch_199_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_445 = imm_switch_199_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_446 = imm_switch_200_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_447 = imm_switch_200_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_448 = imm_switch_201_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_449 = imm_switch_201_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_450 = imm_switch_202_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_451 = imm_switch_202_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_452 = imm_switch_203_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_453 = imm_switch_203_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_454 = imm_switch_204_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_455 = imm_switch_204_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_456 = imm_switch_205_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_457 = imm_switch_205_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_458 = imm_switch_206_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_459 = imm_switch_206_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_460 = in_switch_23_io_y; // @[Benes.scala 80:29 92:43]
  wire [15:0] w_internal_461 = in_switch_23_io_z; // @[Benes.scala 80:29 93:43]
  wire [15:0] w_internal_462 = imm_switch_207_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_463 = imm_switch_207_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_464 = imm_switch_208_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_465 = imm_switch_208_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_466 = imm_switch_209_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_467 = imm_switch_209_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_468 = imm_switch_210_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_469 = imm_switch_210_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_470 = imm_switch_211_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_471 = imm_switch_211_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_472 = imm_switch_212_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_473 = imm_switch_212_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_474 = imm_switch_213_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_475 = imm_switch_213_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_476 = imm_switch_214_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_477 = imm_switch_214_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_478 = imm_switch_215_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_479 = imm_switch_215_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_480 = in_switch_24_io_y; // @[Benes.scala 80:29 92:43]
  wire [15:0] w_internal_481 = in_switch_24_io_z; // @[Benes.scala 80:29 93:43]
  wire [15:0] w_internal_482 = imm_switch_216_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_483 = imm_switch_216_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_484 = imm_switch_217_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_485 = imm_switch_217_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_486 = imm_switch_218_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_487 = imm_switch_218_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_488 = imm_switch_219_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_489 = imm_switch_219_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_490 = imm_switch_220_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_491 = imm_switch_220_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_492 = imm_switch_221_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_493 = imm_switch_221_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_494 = imm_switch_222_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_495 = imm_switch_222_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_496 = imm_switch_223_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_497 = imm_switch_223_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_498 = imm_switch_224_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_499 = imm_switch_224_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_500 = in_switch_25_io_y; // @[Benes.scala 80:29 92:43]
  wire [15:0] w_internal_501 = in_switch_25_io_z; // @[Benes.scala 80:29 93:43]
  wire [15:0] w_internal_502 = imm_switch_225_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_503 = imm_switch_225_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_504 = imm_switch_226_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_505 = imm_switch_226_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_506 = imm_switch_227_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_507 = imm_switch_227_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_508 = imm_switch_228_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_509 = imm_switch_228_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_510 = imm_switch_229_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_511 = imm_switch_229_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_512 = imm_switch_230_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_513 = imm_switch_230_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_514 = imm_switch_231_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_515 = imm_switch_231_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_516 = imm_switch_232_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_517 = imm_switch_232_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_518 = imm_switch_233_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_519 = imm_switch_233_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_520 = in_switch_26_io_y; // @[Benes.scala 80:29 92:43]
  wire [15:0] w_internal_521 = in_switch_26_io_z; // @[Benes.scala 80:29 93:43]
  wire [15:0] w_internal_522 = imm_switch_234_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_523 = imm_switch_234_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_524 = imm_switch_235_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_525 = imm_switch_235_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_526 = imm_switch_236_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_527 = imm_switch_236_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_528 = imm_switch_237_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_529 = imm_switch_237_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_530 = imm_switch_238_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_531 = imm_switch_238_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_532 = imm_switch_239_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_533 = imm_switch_239_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_534 = imm_switch_240_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_535 = imm_switch_240_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_536 = imm_switch_241_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_537 = imm_switch_241_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_538 = imm_switch_242_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_539 = imm_switch_242_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_540 = in_switch_27_io_y; // @[Benes.scala 80:29 92:43]
  wire [15:0] w_internal_541 = in_switch_27_io_z; // @[Benes.scala 80:29 93:43]
  wire [15:0] w_internal_542 = imm_switch_243_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_543 = imm_switch_243_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_544 = imm_switch_244_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_545 = imm_switch_244_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_546 = imm_switch_245_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_547 = imm_switch_245_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_548 = imm_switch_246_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_549 = imm_switch_246_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_550 = imm_switch_247_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_551 = imm_switch_247_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_552 = imm_switch_248_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_553 = imm_switch_248_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_554 = imm_switch_249_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_555 = imm_switch_249_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_556 = imm_switch_250_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_557 = imm_switch_250_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_558 = imm_switch_251_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_559 = imm_switch_251_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_560 = in_switch_28_io_y; // @[Benes.scala 80:29 92:43]
  wire [15:0] w_internal_561 = in_switch_28_io_z; // @[Benes.scala 80:29 93:43]
  wire [15:0] w_internal_562 = imm_switch_252_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_563 = imm_switch_252_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_564 = imm_switch_253_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_565 = imm_switch_253_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_566 = imm_switch_254_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_567 = imm_switch_254_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_568 = imm_switch_255_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_569 = imm_switch_255_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_570 = imm_switch_256_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_571 = imm_switch_256_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_572 = imm_switch_257_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_573 = imm_switch_257_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_574 = imm_switch_258_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_575 = imm_switch_258_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_576 = imm_switch_259_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_577 = imm_switch_259_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_578 = imm_switch_260_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_579 = imm_switch_260_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_580 = in_switch_29_io_y; // @[Benes.scala 80:29 92:43]
  wire [15:0] w_internal_581 = in_switch_29_io_z; // @[Benes.scala 80:29 93:43]
  wire [15:0] w_internal_582 = imm_switch_261_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_583 = imm_switch_261_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_584 = imm_switch_262_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_585 = imm_switch_262_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_586 = imm_switch_263_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_587 = imm_switch_263_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_588 = imm_switch_264_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_589 = imm_switch_264_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_590 = imm_switch_265_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_591 = imm_switch_265_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_592 = imm_switch_266_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_593 = imm_switch_266_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_594 = imm_switch_267_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_595 = imm_switch_267_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_596 = imm_switch_268_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_597 = imm_switch_268_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_598 = imm_switch_269_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_599 = imm_switch_269_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_600 = in_switch_30_io_y; // @[Benes.scala 80:29 92:43]
  wire [15:0] w_internal_601 = in_switch_30_io_z; // @[Benes.scala 80:29 93:43]
  wire [15:0] w_internal_602 = imm_switch_270_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_603 = imm_switch_270_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_604 = imm_switch_271_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_605 = imm_switch_271_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_606 = imm_switch_272_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_607 = imm_switch_272_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_608 = imm_switch_273_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_609 = imm_switch_273_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_610 = imm_switch_274_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_611 = imm_switch_274_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_612 = imm_switch_275_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_613 = imm_switch_275_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_614 = imm_switch_276_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_615 = imm_switch_276_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_616 = imm_switch_277_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_617 = imm_switch_277_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_618 = imm_switch_278_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_619 = imm_switch_278_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_620 = in_switch_31_io_y; // @[Benes.scala 80:29 92:43]
  wire [15:0] w_internal_621 = in_switch_31_io_z; // @[Benes.scala 80:29 93:43]
  wire [15:0] w_internal_622 = imm_switch_279_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_623 = imm_switch_279_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_624 = imm_switch_280_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_625 = imm_switch_280_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_626 = imm_switch_281_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_627 = imm_switch_281_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_628 = imm_switch_282_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_629 = imm_switch_282_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_630 = imm_switch_283_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_631 = imm_switch_283_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_632 = imm_switch_284_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_633 = imm_switch_284_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_634 = imm_switch_285_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_635 = imm_switch_285_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_636 = imm_switch_286_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_637 = imm_switch_286_io_z; // @[Benes.scala 80:29 127:53]
  wire [15:0] w_internal_638 = imm_switch_287_io_y; // @[Benes.scala 80:29 126:53]
  wire [15:0] w_internal_639 = imm_switch_287_io_z; // @[Benes.scala 80:29 127:53]
  InputSwitch in_switch ( // @[Benes.scala 90:27]
    .io_y(in_switch_io_y),
    .io_z(in_switch_io_z),
    .io_in(in_switch_io_in)
  );
  InputSwitch in_switch_1 ( // @[Benes.scala 90:27]
    .io_y(in_switch_1_io_y),
    .io_z(in_switch_1_io_z),
    .io_in(in_switch_1_io_in)
  );
  InputSwitch in_switch_2 ( // @[Benes.scala 90:27]
    .io_y(in_switch_2_io_y),
    .io_z(in_switch_2_io_z),
    .io_in(in_switch_2_io_in)
  );
  InputSwitch in_switch_3 ( // @[Benes.scala 90:27]
    .io_y(in_switch_3_io_y),
    .io_z(in_switch_3_io_z),
    .io_in(in_switch_3_io_in)
  );
  InputSwitch in_switch_4 ( // @[Benes.scala 90:27]
    .io_y(in_switch_4_io_y),
    .io_z(in_switch_4_io_z),
    .io_in(in_switch_4_io_in)
  );
  InputSwitch in_switch_5 ( // @[Benes.scala 90:27]
    .io_y(in_switch_5_io_y),
    .io_z(in_switch_5_io_z),
    .io_in(in_switch_5_io_in)
  );
  InputSwitch in_switch_6 ( // @[Benes.scala 90:27]
    .io_y(in_switch_6_io_y),
    .io_z(in_switch_6_io_z),
    .io_in(in_switch_6_io_in)
  );
  InputSwitch in_switch_7 ( // @[Benes.scala 90:27]
    .io_y(in_switch_7_io_y),
    .io_z(in_switch_7_io_z),
    .io_in(in_switch_7_io_in)
  );
  InputSwitch in_switch_8 ( // @[Benes.scala 90:27]
    .io_y(in_switch_8_io_y),
    .io_z(in_switch_8_io_z),
    .io_in(in_switch_8_io_in)
  );
  InputSwitch in_switch_9 ( // @[Benes.scala 90:27]
    .io_y(in_switch_9_io_y),
    .io_z(in_switch_9_io_z),
    .io_in(in_switch_9_io_in)
  );
  InputSwitch in_switch_10 ( // @[Benes.scala 90:27]
    .io_y(in_switch_10_io_y),
    .io_z(in_switch_10_io_z),
    .io_in(in_switch_10_io_in)
  );
  InputSwitch in_switch_11 ( // @[Benes.scala 90:27]
    .io_y(in_switch_11_io_y),
    .io_z(in_switch_11_io_z),
    .io_in(in_switch_11_io_in)
  );
  InputSwitch in_switch_12 ( // @[Benes.scala 90:27]
    .io_y(in_switch_12_io_y),
    .io_z(in_switch_12_io_z),
    .io_in(in_switch_12_io_in)
  );
  InputSwitch in_switch_13 ( // @[Benes.scala 90:27]
    .io_y(in_switch_13_io_y),
    .io_z(in_switch_13_io_z),
    .io_in(in_switch_13_io_in)
  );
  InputSwitch in_switch_14 ( // @[Benes.scala 90:27]
    .io_y(in_switch_14_io_y),
    .io_z(in_switch_14_io_z),
    .io_in(in_switch_14_io_in)
  );
  InputSwitch in_switch_15 ( // @[Benes.scala 90:27]
    .io_y(in_switch_15_io_y),
    .io_z(in_switch_15_io_z),
    .io_in(in_switch_15_io_in)
  );
  InputSwitch in_switch_16 ( // @[Benes.scala 90:27]
    .io_y(in_switch_16_io_y),
    .io_z(in_switch_16_io_z),
    .io_in(in_switch_16_io_in)
  );
  InputSwitch in_switch_17 ( // @[Benes.scala 90:27]
    .io_y(in_switch_17_io_y),
    .io_z(in_switch_17_io_z),
    .io_in(in_switch_17_io_in)
  );
  InputSwitch in_switch_18 ( // @[Benes.scala 90:27]
    .io_y(in_switch_18_io_y),
    .io_z(in_switch_18_io_z),
    .io_in(in_switch_18_io_in)
  );
  InputSwitch in_switch_19 ( // @[Benes.scala 90:27]
    .io_y(in_switch_19_io_y),
    .io_z(in_switch_19_io_z),
    .io_in(in_switch_19_io_in)
  );
  InputSwitch in_switch_20 ( // @[Benes.scala 90:27]
    .io_y(in_switch_20_io_y),
    .io_z(in_switch_20_io_z),
    .io_in(in_switch_20_io_in)
  );
  InputSwitch in_switch_21 ( // @[Benes.scala 90:27]
    .io_y(in_switch_21_io_y),
    .io_z(in_switch_21_io_z),
    .io_in(in_switch_21_io_in)
  );
  InputSwitch in_switch_22 ( // @[Benes.scala 90:27]
    .io_y(in_switch_22_io_y),
    .io_z(in_switch_22_io_z),
    .io_in(in_switch_22_io_in)
  );
  InputSwitch in_switch_23 ( // @[Benes.scala 90:27]
    .io_y(in_switch_23_io_y),
    .io_z(in_switch_23_io_z),
    .io_in(in_switch_23_io_in)
  );
  InputSwitch in_switch_24 ( // @[Benes.scala 90:27]
    .io_y(in_switch_24_io_y),
    .io_z(in_switch_24_io_z),
    .io_in(in_switch_24_io_in)
  );
  InputSwitch in_switch_25 ( // @[Benes.scala 90:27]
    .io_y(in_switch_25_io_y),
    .io_z(in_switch_25_io_z),
    .io_in(in_switch_25_io_in)
  );
  InputSwitch in_switch_26 ( // @[Benes.scala 90:27]
    .io_y(in_switch_26_io_y),
    .io_z(in_switch_26_io_z),
    .io_in(in_switch_26_io_in)
  );
  InputSwitch in_switch_27 ( // @[Benes.scala 90:27]
    .io_y(in_switch_27_io_y),
    .io_z(in_switch_27_io_z),
    .io_in(in_switch_27_io_in)
  );
  InputSwitch in_switch_28 ( // @[Benes.scala 90:27]
    .io_y(in_switch_28_io_y),
    .io_z(in_switch_28_io_z),
    .io_in(in_switch_28_io_in)
  );
  InputSwitch in_switch_29 ( // @[Benes.scala 90:27]
    .io_y(in_switch_29_io_y),
    .io_z(in_switch_29_io_z),
    .io_in(in_switch_29_io_in)
  );
  InputSwitch in_switch_30 ( // @[Benes.scala 90:27]
    .io_y(in_switch_30_io_y),
    .io_z(in_switch_30_io_z),
    .io_in(in_switch_30_io_in)
  );
  InputSwitch in_switch_31 ( // @[Benes.scala 90:27]
    .io_y(in_switch_31_io_y),
    .io_z(in_switch_31_io_z),
    .io_in(in_switch_31_io_in)
  );
  OutputSwitch out_switch ( // @[Benes.scala 99:28]
    .io_y(out_switch_io_y),
    .io_in0(out_switch_io_in0)
  );
  OutputSwitch out_switch_1 ( // @[Benes.scala 99:28]
    .io_y(out_switch_1_io_y),
    .io_in0(out_switch_1_io_in0)
  );
  OutputSwitch out_switch_2 ( // @[Benes.scala 99:28]
    .io_y(out_switch_2_io_y),
    .io_in0(out_switch_2_io_in0)
  );
  OutputSwitch out_switch_3 ( // @[Benes.scala 99:28]
    .io_y(out_switch_3_io_y),
    .io_in0(out_switch_3_io_in0)
  );
  OutputSwitch out_switch_4 ( // @[Benes.scala 99:28]
    .io_y(out_switch_4_io_y),
    .io_in0(out_switch_4_io_in0)
  );
  OutputSwitch out_switch_5 ( // @[Benes.scala 99:28]
    .io_y(out_switch_5_io_y),
    .io_in0(out_switch_5_io_in0)
  );
  OutputSwitch out_switch_6 ( // @[Benes.scala 99:28]
    .io_y(out_switch_6_io_y),
    .io_in0(out_switch_6_io_in0)
  );
  OutputSwitch out_switch_7 ( // @[Benes.scala 99:28]
    .io_y(out_switch_7_io_y),
    .io_in0(out_switch_7_io_in0)
  );
  OutputSwitch out_switch_8 ( // @[Benes.scala 99:28]
    .io_y(out_switch_8_io_y),
    .io_in0(out_switch_8_io_in0)
  );
  OutputSwitch out_switch_9 ( // @[Benes.scala 99:28]
    .io_y(out_switch_9_io_y),
    .io_in0(out_switch_9_io_in0)
  );
  OutputSwitch out_switch_10 ( // @[Benes.scala 99:28]
    .io_y(out_switch_10_io_y),
    .io_in0(out_switch_10_io_in0)
  );
  OutputSwitch out_switch_11 ( // @[Benes.scala 99:28]
    .io_y(out_switch_11_io_y),
    .io_in0(out_switch_11_io_in0)
  );
  OutputSwitch out_switch_12 ( // @[Benes.scala 99:28]
    .io_y(out_switch_12_io_y),
    .io_in0(out_switch_12_io_in0)
  );
  OutputSwitch out_switch_13 ( // @[Benes.scala 99:28]
    .io_y(out_switch_13_io_y),
    .io_in0(out_switch_13_io_in0)
  );
  OutputSwitch out_switch_14 ( // @[Benes.scala 99:28]
    .io_y(out_switch_14_io_y),
    .io_in0(out_switch_14_io_in0)
  );
  OutputSwitch out_switch_15 ( // @[Benes.scala 99:28]
    .io_y(out_switch_15_io_y),
    .io_in0(out_switch_15_io_in0)
  );
  OutputSwitch out_switch_16 ( // @[Benes.scala 99:28]
    .io_y(out_switch_16_io_y),
    .io_in0(out_switch_16_io_in0)
  );
  OutputSwitch out_switch_17 ( // @[Benes.scala 99:28]
    .io_y(out_switch_17_io_y),
    .io_in0(out_switch_17_io_in0)
  );
  OutputSwitch out_switch_18 ( // @[Benes.scala 99:28]
    .io_y(out_switch_18_io_y),
    .io_in0(out_switch_18_io_in0)
  );
  OutputSwitch out_switch_19 ( // @[Benes.scala 99:28]
    .io_y(out_switch_19_io_y),
    .io_in0(out_switch_19_io_in0)
  );
  OutputSwitch out_switch_20 ( // @[Benes.scala 99:28]
    .io_y(out_switch_20_io_y),
    .io_in0(out_switch_20_io_in0)
  );
  OutputSwitch out_switch_21 ( // @[Benes.scala 99:28]
    .io_y(out_switch_21_io_y),
    .io_in0(out_switch_21_io_in0)
  );
  OutputSwitch out_switch_22 ( // @[Benes.scala 99:28]
    .io_y(out_switch_22_io_y),
    .io_in0(out_switch_22_io_in0)
  );
  OutputSwitch out_switch_23 ( // @[Benes.scala 99:28]
    .io_y(out_switch_23_io_y),
    .io_in0(out_switch_23_io_in0)
  );
  OutputSwitch out_switch_24 ( // @[Benes.scala 99:28]
    .io_y(out_switch_24_io_y),
    .io_in0(out_switch_24_io_in0)
  );
  OutputSwitch out_switch_25 ( // @[Benes.scala 99:28]
    .io_y(out_switch_25_io_y),
    .io_in0(out_switch_25_io_in0)
  );
  OutputSwitch out_switch_26 ( // @[Benes.scala 99:28]
    .io_y(out_switch_26_io_y),
    .io_in0(out_switch_26_io_in0)
  );
  OutputSwitch out_switch_27 ( // @[Benes.scala 99:28]
    .io_y(out_switch_27_io_y),
    .io_in0(out_switch_27_io_in0)
  );
  OutputSwitch out_switch_28 ( // @[Benes.scala 99:28]
    .io_y(out_switch_28_io_y),
    .io_in0(out_switch_28_io_in0)
  );
  OutputSwitch out_switch_29 ( // @[Benes.scala 99:28]
    .io_y(out_switch_29_io_y),
    .io_in0(out_switch_29_io_in0)
  );
  OutputSwitch out_switch_30 ( // @[Benes.scala 99:28]
    .io_y(out_switch_30_io_y),
    .io_in0(out_switch_30_io_in0)
  );
  OutputSwitch out_switch_31 ( // @[Benes.scala 99:28]
    .io_y(out_switch_31_io_y),
    .io_in0(out_switch_31_io_in0)
  );
  Switch imm_switch ( // @[Benes.scala 109:30]
    .io_y(imm_switch_io_y),
    .io_z(imm_switch_io_z),
    .io_in0(imm_switch_io_in0)
  );
  Switch imm_switch_1 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_1_io_y),
    .io_z(imm_switch_1_io_z),
    .io_in0(imm_switch_1_io_in0)
  );
  Switch imm_switch_2 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_2_io_y),
    .io_z(imm_switch_2_io_z),
    .io_in0(imm_switch_2_io_in0)
  );
  Switch imm_switch_3 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_3_io_y),
    .io_z(imm_switch_3_io_z),
    .io_in0(imm_switch_3_io_in0)
  );
  Switch imm_switch_4 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_4_io_y),
    .io_z(imm_switch_4_io_z),
    .io_in0(imm_switch_4_io_in0)
  );
  Switch imm_switch_5 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_5_io_y),
    .io_z(imm_switch_5_io_z),
    .io_in0(imm_switch_5_io_in0)
  );
  Switch imm_switch_6 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_6_io_y),
    .io_z(imm_switch_6_io_z),
    .io_in0(imm_switch_6_io_in0)
  );
  Switch imm_switch_7 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_7_io_y),
    .io_z(imm_switch_7_io_z),
    .io_in0(imm_switch_7_io_in0)
  );
  Switch imm_switch_8 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_8_io_y),
    .io_z(imm_switch_8_io_z),
    .io_in0(imm_switch_8_io_in0)
  );
  Switch imm_switch_9 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_9_io_y),
    .io_z(imm_switch_9_io_z),
    .io_in0(imm_switch_9_io_in0)
  );
  Switch imm_switch_10 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_10_io_y),
    .io_z(imm_switch_10_io_z),
    .io_in0(imm_switch_10_io_in0)
  );
  Switch imm_switch_11 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_11_io_y),
    .io_z(imm_switch_11_io_z),
    .io_in0(imm_switch_11_io_in0)
  );
  Switch imm_switch_12 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_12_io_y),
    .io_z(imm_switch_12_io_z),
    .io_in0(imm_switch_12_io_in0)
  );
  Switch imm_switch_13 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_13_io_y),
    .io_z(imm_switch_13_io_z),
    .io_in0(imm_switch_13_io_in0)
  );
  Switch imm_switch_14 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_14_io_y),
    .io_z(imm_switch_14_io_z),
    .io_in0(imm_switch_14_io_in0)
  );
  Switch imm_switch_15 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_15_io_y),
    .io_z(imm_switch_15_io_z),
    .io_in0(imm_switch_15_io_in0)
  );
  Switch imm_switch_16 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_16_io_y),
    .io_z(imm_switch_16_io_z),
    .io_in0(imm_switch_16_io_in0)
  );
  Switch imm_switch_17 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_17_io_y),
    .io_z(imm_switch_17_io_z),
    .io_in0(imm_switch_17_io_in0)
  );
  Switch imm_switch_18 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_18_io_y),
    .io_z(imm_switch_18_io_z),
    .io_in0(imm_switch_18_io_in0)
  );
  Switch imm_switch_19 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_19_io_y),
    .io_z(imm_switch_19_io_z),
    .io_in0(imm_switch_19_io_in0)
  );
  Switch imm_switch_20 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_20_io_y),
    .io_z(imm_switch_20_io_z),
    .io_in0(imm_switch_20_io_in0)
  );
  Switch imm_switch_21 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_21_io_y),
    .io_z(imm_switch_21_io_z),
    .io_in0(imm_switch_21_io_in0)
  );
  Switch imm_switch_22 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_22_io_y),
    .io_z(imm_switch_22_io_z),
    .io_in0(imm_switch_22_io_in0)
  );
  Switch imm_switch_23 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_23_io_y),
    .io_z(imm_switch_23_io_z),
    .io_in0(imm_switch_23_io_in0)
  );
  Switch imm_switch_24 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_24_io_y),
    .io_z(imm_switch_24_io_z),
    .io_in0(imm_switch_24_io_in0)
  );
  Switch imm_switch_25 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_25_io_y),
    .io_z(imm_switch_25_io_z),
    .io_in0(imm_switch_25_io_in0)
  );
  Switch imm_switch_26 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_26_io_y),
    .io_z(imm_switch_26_io_z),
    .io_in0(imm_switch_26_io_in0)
  );
  Switch imm_switch_27 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_27_io_y),
    .io_z(imm_switch_27_io_z),
    .io_in0(imm_switch_27_io_in0)
  );
  Switch imm_switch_28 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_28_io_y),
    .io_z(imm_switch_28_io_z),
    .io_in0(imm_switch_28_io_in0)
  );
  Switch imm_switch_29 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_29_io_y),
    .io_z(imm_switch_29_io_z),
    .io_in0(imm_switch_29_io_in0)
  );
  Switch imm_switch_30 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_30_io_y),
    .io_z(imm_switch_30_io_z),
    .io_in0(imm_switch_30_io_in0)
  );
  Switch imm_switch_31 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_31_io_y),
    .io_z(imm_switch_31_io_z),
    .io_in0(imm_switch_31_io_in0)
  );
  Switch imm_switch_32 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_32_io_y),
    .io_z(imm_switch_32_io_z),
    .io_in0(imm_switch_32_io_in0)
  );
  Switch imm_switch_33 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_33_io_y),
    .io_z(imm_switch_33_io_z),
    .io_in0(imm_switch_33_io_in0)
  );
  Switch imm_switch_34 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_34_io_y),
    .io_z(imm_switch_34_io_z),
    .io_in0(imm_switch_34_io_in0)
  );
  Switch imm_switch_35 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_35_io_y),
    .io_z(imm_switch_35_io_z),
    .io_in0(imm_switch_35_io_in0)
  );
  Switch imm_switch_36 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_36_io_y),
    .io_z(imm_switch_36_io_z),
    .io_in0(imm_switch_36_io_in0)
  );
  Switch imm_switch_37 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_37_io_y),
    .io_z(imm_switch_37_io_z),
    .io_in0(imm_switch_37_io_in0)
  );
  Switch imm_switch_38 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_38_io_y),
    .io_z(imm_switch_38_io_z),
    .io_in0(imm_switch_38_io_in0)
  );
  Switch imm_switch_39 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_39_io_y),
    .io_z(imm_switch_39_io_z),
    .io_in0(imm_switch_39_io_in0)
  );
  Switch imm_switch_40 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_40_io_y),
    .io_z(imm_switch_40_io_z),
    .io_in0(imm_switch_40_io_in0)
  );
  Switch imm_switch_41 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_41_io_y),
    .io_z(imm_switch_41_io_z),
    .io_in0(imm_switch_41_io_in0)
  );
  Switch imm_switch_42 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_42_io_y),
    .io_z(imm_switch_42_io_z),
    .io_in0(imm_switch_42_io_in0)
  );
  Switch imm_switch_43 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_43_io_y),
    .io_z(imm_switch_43_io_z),
    .io_in0(imm_switch_43_io_in0)
  );
  Switch imm_switch_44 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_44_io_y),
    .io_z(imm_switch_44_io_z),
    .io_in0(imm_switch_44_io_in0)
  );
  Switch imm_switch_45 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_45_io_y),
    .io_z(imm_switch_45_io_z),
    .io_in0(imm_switch_45_io_in0)
  );
  Switch imm_switch_46 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_46_io_y),
    .io_z(imm_switch_46_io_z),
    .io_in0(imm_switch_46_io_in0)
  );
  Switch imm_switch_47 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_47_io_y),
    .io_z(imm_switch_47_io_z),
    .io_in0(imm_switch_47_io_in0)
  );
  Switch imm_switch_48 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_48_io_y),
    .io_z(imm_switch_48_io_z),
    .io_in0(imm_switch_48_io_in0)
  );
  Switch imm_switch_49 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_49_io_y),
    .io_z(imm_switch_49_io_z),
    .io_in0(imm_switch_49_io_in0)
  );
  Switch imm_switch_50 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_50_io_y),
    .io_z(imm_switch_50_io_z),
    .io_in0(imm_switch_50_io_in0)
  );
  Switch imm_switch_51 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_51_io_y),
    .io_z(imm_switch_51_io_z),
    .io_in0(imm_switch_51_io_in0)
  );
  Switch imm_switch_52 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_52_io_y),
    .io_z(imm_switch_52_io_z),
    .io_in0(imm_switch_52_io_in0)
  );
  Switch imm_switch_53 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_53_io_y),
    .io_z(imm_switch_53_io_z),
    .io_in0(imm_switch_53_io_in0)
  );
  Switch imm_switch_54 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_54_io_y),
    .io_z(imm_switch_54_io_z),
    .io_in0(imm_switch_54_io_in0)
  );
  Switch imm_switch_55 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_55_io_y),
    .io_z(imm_switch_55_io_z),
    .io_in0(imm_switch_55_io_in0)
  );
  Switch imm_switch_56 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_56_io_y),
    .io_z(imm_switch_56_io_z),
    .io_in0(imm_switch_56_io_in0)
  );
  Switch imm_switch_57 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_57_io_y),
    .io_z(imm_switch_57_io_z),
    .io_in0(imm_switch_57_io_in0)
  );
  Switch imm_switch_58 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_58_io_y),
    .io_z(imm_switch_58_io_z),
    .io_in0(imm_switch_58_io_in0)
  );
  Switch imm_switch_59 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_59_io_y),
    .io_z(imm_switch_59_io_z),
    .io_in0(imm_switch_59_io_in0)
  );
  Switch imm_switch_60 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_60_io_y),
    .io_z(imm_switch_60_io_z),
    .io_in0(imm_switch_60_io_in0)
  );
  Switch imm_switch_61 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_61_io_y),
    .io_z(imm_switch_61_io_z),
    .io_in0(imm_switch_61_io_in0)
  );
  Switch imm_switch_62 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_62_io_y),
    .io_z(imm_switch_62_io_z),
    .io_in0(imm_switch_62_io_in0)
  );
  Switch imm_switch_63 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_63_io_y),
    .io_z(imm_switch_63_io_z),
    .io_in0(imm_switch_63_io_in0)
  );
  Switch imm_switch_64 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_64_io_y),
    .io_z(imm_switch_64_io_z),
    .io_in0(imm_switch_64_io_in0)
  );
  Switch imm_switch_65 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_65_io_y),
    .io_z(imm_switch_65_io_z),
    .io_in0(imm_switch_65_io_in0)
  );
  Switch imm_switch_66 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_66_io_y),
    .io_z(imm_switch_66_io_z),
    .io_in0(imm_switch_66_io_in0)
  );
  Switch imm_switch_67 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_67_io_y),
    .io_z(imm_switch_67_io_z),
    .io_in0(imm_switch_67_io_in0)
  );
  Switch imm_switch_68 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_68_io_y),
    .io_z(imm_switch_68_io_z),
    .io_in0(imm_switch_68_io_in0)
  );
  Switch imm_switch_69 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_69_io_y),
    .io_z(imm_switch_69_io_z),
    .io_in0(imm_switch_69_io_in0)
  );
  Switch imm_switch_70 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_70_io_y),
    .io_z(imm_switch_70_io_z),
    .io_in0(imm_switch_70_io_in0)
  );
  Switch imm_switch_71 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_71_io_y),
    .io_z(imm_switch_71_io_z),
    .io_in0(imm_switch_71_io_in0)
  );
  Switch imm_switch_72 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_72_io_y),
    .io_z(imm_switch_72_io_z),
    .io_in0(imm_switch_72_io_in0)
  );
  Switch imm_switch_73 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_73_io_y),
    .io_z(imm_switch_73_io_z),
    .io_in0(imm_switch_73_io_in0)
  );
  Switch imm_switch_74 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_74_io_y),
    .io_z(imm_switch_74_io_z),
    .io_in0(imm_switch_74_io_in0)
  );
  Switch imm_switch_75 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_75_io_y),
    .io_z(imm_switch_75_io_z),
    .io_in0(imm_switch_75_io_in0)
  );
  Switch imm_switch_76 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_76_io_y),
    .io_z(imm_switch_76_io_z),
    .io_in0(imm_switch_76_io_in0)
  );
  Switch imm_switch_77 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_77_io_y),
    .io_z(imm_switch_77_io_z),
    .io_in0(imm_switch_77_io_in0)
  );
  Switch imm_switch_78 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_78_io_y),
    .io_z(imm_switch_78_io_z),
    .io_in0(imm_switch_78_io_in0)
  );
  Switch imm_switch_79 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_79_io_y),
    .io_z(imm_switch_79_io_z),
    .io_in0(imm_switch_79_io_in0)
  );
  Switch imm_switch_80 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_80_io_y),
    .io_z(imm_switch_80_io_z),
    .io_in0(imm_switch_80_io_in0)
  );
  Switch imm_switch_81 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_81_io_y),
    .io_z(imm_switch_81_io_z),
    .io_in0(imm_switch_81_io_in0)
  );
  Switch imm_switch_82 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_82_io_y),
    .io_z(imm_switch_82_io_z),
    .io_in0(imm_switch_82_io_in0)
  );
  Switch imm_switch_83 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_83_io_y),
    .io_z(imm_switch_83_io_z),
    .io_in0(imm_switch_83_io_in0)
  );
  Switch imm_switch_84 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_84_io_y),
    .io_z(imm_switch_84_io_z),
    .io_in0(imm_switch_84_io_in0)
  );
  Switch imm_switch_85 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_85_io_y),
    .io_z(imm_switch_85_io_z),
    .io_in0(imm_switch_85_io_in0)
  );
  Switch imm_switch_86 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_86_io_y),
    .io_z(imm_switch_86_io_z),
    .io_in0(imm_switch_86_io_in0)
  );
  Switch imm_switch_87 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_87_io_y),
    .io_z(imm_switch_87_io_z),
    .io_in0(imm_switch_87_io_in0)
  );
  Switch imm_switch_88 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_88_io_y),
    .io_z(imm_switch_88_io_z),
    .io_in0(imm_switch_88_io_in0)
  );
  Switch imm_switch_89 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_89_io_y),
    .io_z(imm_switch_89_io_z),
    .io_in0(imm_switch_89_io_in0)
  );
  Switch imm_switch_90 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_90_io_y),
    .io_z(imm_switch_90_io_z),
    .io_in0(imm_switch_90_io_in0)
  );
  Switch imm_switch_91 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_91_io_y),
    .io_z(imm_switch_91_io_z),
    .io_in0(imm_switch_91_io_in0)
  );
  Switch imm_switch_92 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_92_io_y),
    .io_z(imm_switch_92_io_z),
    .io_in0(imm_switch_92_io_in0)
  );
  Switch imm_switch_93 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_93_io_y),
    .io_z(imm_switch_93_io_z),
    .io_in0(imm_switch_93_io_in0)
  );
  Switch imm_switch_94 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_94_io_y),
    .io_z(imm_switch_94_io_z),
    .io_in0(imm_switch_94_io_in0)
  );
  Switch imm_switch_95 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_95_io_y),
    .io_z(imm_switch_95_io_z),
    .io_in0(imm_switch_95_io_in0)
  );
  Switch imm_switch_96 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_96_io_y),
    .io_z(imm_switch_96_io_z),
    .io_in0(imm_switch_96_io_in0)
  );
  Switch imm_switch_97 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_97_io_y),
    .io_z(imm_switch_97_io_z),
    .io_in0(imm_switch_97_io_in0)
  );
  Switch imm_switch_98 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_98_io_y),
    .io_z(imm_switch_98_io_z),
    .io_in0(imm_switch_98_io_in0)
  );
  Switch imm_switch_99 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_99_io_y),
    .io_z(imm_switch_99_io_z),
    .io_in0(imm_switch_99_io_in0)
  );
  Switch imm_switch_100 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_100_io_y),
    .io_z(imm_switch_100_io_z),
    .io_in0(imm_switch_100_io_in0)
  );
  Switch imm_switch_101 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_101_io_y),
    .io_z(imm_switch_101_io_z),
    .io_in0(imm_switch_101_io_in0)
  );
  Switch imm_switch_102 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_102_io_y),
    .io_z(imm_switch_102_io_z),
    .io_in0(imm_switch_102_io_in0)
  );
  Switch imm_switch_103 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_103_io_y),
    .io_z(imm_switch_103_io_z),
    .io_in0(imm_switch_103_io_in0)
  );
  Switch imm_switch_104 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_104_io_y),
    .io_z(imm_switch_104_io_z),
    .io_in0(imm_switch_104_io_in0)
  );
  Switch imm_switch_105 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_105_io_y),
    .io_z(imm_switch_105_io_z),
    .io_in0(imm_switch_105_io_in0)
  );
  Switch imm_switch_106 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_106_io_y),
    .io_z(imm_switch_106_io_z),
    .io_in0(imm_switch_106_io_in0)
  );
  Switch imm_switch_107 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_107_io_y),
    .io_z(imm_switch_107_io_z),
    .io_in0(imm_switch_107_io_in0)
  );
  Switch imm_switch_108 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_108_io_y),
    .io_z(imm_switch_108_io_z),
    .io_in0(imm_switch_108_io_in0)
  );
  Switch imm_switch_109 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_109_io_y),
    .io_z(imm_switch_109_io_z),
    .io_in0(imm_switch_109_io_in0)
  );
  Switch imm_switch_110 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_110_io_y),
    .io_z(imm_switch_110_io_z),
    .io_in0(imm_switch_110_io_in0)
  );
  Switch imm_switch_111 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_111_io_y),
    .io_z(imm_switch_111_io_z),
    .io_in0(imm_switch_111_io_in0)
  );
  Switch imm_switch_112 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_112_io_y),
    .io_z(imm_switch_112_io_z),
    .io_in0(imm_switch_112_io_in0)
  );
  Switch imm_switch_113 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_113_io_y),
    .io_z(imm_switch_113_io_z),
    .io_in0(imm_switch_113_io_in0)
  );
  Switch imm_switch_114 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_114_io_y),
    .io_z(imm_switch_114_io_z),
    .io_in0(imm_switch_114_io_in0)
  );
  Switch imm_switch_115 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_115_io_y),
    .io_z(imm_switch_115_io_z),
    .io_in0(imm_switch_115_io_in0)
  );
  Switch imm_switch_116 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_116_io_y),
    .io_z(imm_switch_116_io_z),
    .io_in0(imm_switch_116_io_in0)
  );
  Switch imm_switch_117 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_117_io_y),
    .io_z(imm_switch_117_io_z),
    .io_in0(imm_switch_117_io_in0)
  );
  Switch imm_switch_118 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_118_io_y),
    .io_z(imm_switch_118_io_z),
    .io_in0(imm_switch_118_io_in0)
  );
  Switch imm_switch_119 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_119_io_y),
    .io_z(imm_switch_119_io_z),
    .io_in0(imm_switch_119_io_in0)
  );
  Switch imm_switch_120 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_120_io_y),
    .io_z(imm_switch_120_io_z),
    .io_in0(imm_switch_120_io_in0)
  );
  Switch imm_switch_121 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_121_io_y),
    .io_z(imm_switch_121_io_z),
    .io_in0(imm_switch_121_io_in0)
  );
  Switch imm_switch_122 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_122_io_y),
    .io_z(imm_switch_122_io_z),
    .io_in0(imm_switch_122_io_in0)
  );
  Switch imm_switch_123 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_123_io_y),
    .io_z(imm_switch_123_io_z),
    .io_in0(imm_switch_123_io_in0)
  );
  Switch imm_switch_124 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_124_io_y),
    .io_z(imm_switch_124_io_z),
    .io_in0(imm_switch_124_io_in0)
  );
  Switch imm_switch_125 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_125_io_y),
    .io_z(imm_switch_125_io_z),
    .io_in0(imm_switch_125_io_in0)
  );
  Switch imm_switch_126 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_126_io_y),
    .io_z(imm_switch_126_io_z),
    .io_in0(imm_switch_126_io_in0)
  );
  Switch imm_switch_127 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_127_io_y),
    .io_z(imm_switch_127_io_z),
    .io_in0(imm_switch_127_io_in0)
  );
  Switch imm_switch_128 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_128_io_y),
    .io_z(imm_switch_128_io_z),
    .io_in0(imm_switch_128_io_in0)
  );
  Switch imm_switch_129 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_129_io_y),
    .io_z(imm_switch_129_io_z),
    .io_in0(imm_switch_129_io_in0)
  );
  Switch imm_switch_130 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_130_io_y),
    .io_z(imm_switch_130_io_z),
    .io_in0(imm_switch_130_io_in0)
  );
  Switch imm_switch_131 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_131_io_y),
    .io_z(imm_switch_131_io_z),
    .io_in0(imm_switch_131_io_in0)
  );
  Switch imm_switch_132 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_132_io_y),
    .io_z(imm_switch_132_io_z),
    .io_in0(imm_switch_132_io_in0)
  );
  Switch imm_switch_133 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_133_io_y),
    .io_z(imm_switch_133_io_z),
    .io_in0(imm_switch_133_io_in0)
  );
  Switch imm_switch_134 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_134_io_y),
    .io_z(imm_switch_134_io_z),
    .io_in0(imm_switch_134_io_in0)
  );
  Switch imm_switch_135 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_135_io_y),
    .io_z(imm_switch_135_io_z),
    .io_in0(imm_switch_135_io_in0)
  );
  Switch imm_switch_136 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_136_io_y),
    .io_z(imm_switch_136_io_z),
    .io_in0(imm_switch_136_io_in0)
  );
  Switch imm_switch_137 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_137_io_y),
    .io_z(imm_switch_137_io_z),
    .io_in0(imm_switch_137_io_in0)
  );
  Switch imm_switch_138 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_138_io_y),
    .io_z(imm_switch_138_io_z),
    .io_in0(imm_switch_138_io_in0)
  );
  Switch imm_switch_139 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_139_io_y),
    .io_z(imm_switch_139_io_z),
    .io_in0(imm_switch_139_io_in0)
  );
  Switch imm_switch_140 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_140_io_y),
    .io_z(imm_switch_140_io_z),
    .io_in0(imm_switch_140_io_in0)
  );
  Switch imm_switch_141 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_141_io_y),
    .io_z(imm_switch_141_io_z),
    .io_in0(imm_switch_141_io_in0)
  );
  Switch imm_switch_142 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_142_io_y),
    .io_z(imm_switch_142_io_z),
    .io_in0(imm_switch_142_io_in0)
  );
  Switch imm_switch_143 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_143_io_y),
    .io_z(imm_switch_143_io_z),
    .io_in0(imm_switch_143_io_in0)
  );
  Switch imm_switch_144 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_144_io_y),
    .io_z(imm_switch_144_io_z),
    .io_in0(imm_switch_144_io_in0)
  );
  Switch imm_switch_145 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_145_io_y),
    .io_z(imm_switch_145_io_z),
    .io_in0(imm_switch_145_io_in0)
  );
  Switch imm_switch_146 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_146_io_y),
    .io_z(imm_switch_146_io_z),
    .io_in0(imm_switch_146_io_in0)
  );
  Switch imm_switch_147 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_147_io_y),
    .io_z(imm_switch_147_io_z),
    .io_in0(imm_switch_147_io_in0)
  );
  Switch imm_switch_148 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_148_io_y),
    .io_z(imm_switch_148_io_z),
    .io_in0(imm_switch_148_io_in0)
  );
  Switch imm_switch_149 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_149_io_y),
    .io_z(imm_switch_149_io_z),
    .io_in0(imm_switch_149_io_in0)
  );
  Switch imm_switch_150 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_150_io_y),
    .io_z(imm_switch_150_io_z),
    .io_in0(imm_switch_150_io_in0)
  );
  Switch imm_switch_151 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_151_io_y),
    .io_z(imm_switch_151_io_z),
    .io_in0(imm_switch_151_io_in0)
  );
  Switch imm_switch_152 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_152_io_y),
    .io_z(imm_switch_152_io_z),
    .io_in0(imm_switch_152_io_in0)
  );
  Switch imm_switch_153 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_153_io_y),
    .io_z(imm_switch_153_io_z),
    .io_in0(imm_switch_153_io_in0)
  );
  Switch imm_switch_154 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_154_io_y),
    .io_z(imm_switch_154_io_z),
    .io_in0(imm_switch_154_io_in0)
  );
  Switch imm_switch_155 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_155_io_y),
    .io_z(imm_switch_155_io_z),
    .io_in0(imm_switch_155_io_in0)
  );
  Switch imm_switch_156 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_156_io_y),
    .io_z(imm_switch_156_io_z),
    .io_in0(imm_switch_156_io_in0)
  );
  Switch imm_switch_157 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_157_io_y),
    .io_z(imm_switch_157_io_z),
    .io_in0(imm_switch_157_io_in0)
  );
  Switch imm_switch_158 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_158_io_y),
    .io_z(imm_switch_158_io_z),
    .io_in0(imm_switch_158_io_in0)
  );
  Switch imm_switch_159 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_159_io_y),
    .io_z(imm_switch_159_io_z),
    .io_in0(imm_switch_159_io_in0)
  );
  Switch imm_switch_160 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_160_io_y),
    .io_z(imm_switch_160_io_z),
    .io_in0(imm_switch_160_io_in0)
  );
  Switch imm_switch_161 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_161_io_y),
    .io_z(imm_switch_161_io_z),
    .io_in0(imm_switch_161_io_in0)
  );
  Switch imm_switch_162 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_162_io_y),
    .io_z(imm_switch_162_io_z),
    .io_in0(imm_switch_162_io_in0)
  );
  Switch imm_switch_163 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_163_io_y),
    .io_z(imm_switch_163_io_z),
    .io_in0(imm_switch_163_io_in0)
  );
  Switch imm_switch_164 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_164_io_y),
    .io_z(imm_switch_164_io_z),
    .io_in0(imm_switch_164_io_in0)
  );
  Switch imm_switch_165 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_165_io_y),
    .io_z(imm_switch_165_io_z),
    .io_in0(imm_switch_165_io_in0)
  );
  Switch imm_switch_166 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_166_io_y),
    .io_z(imm_switch_166_io_z),
    .io_in0(imm_switch_166_io_in0)
  );
  Switch imm_switch_167 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_167_io_y),
    .io_z(imm_switch_167_io_z),
    .io_in0(imm_switch_167_io_in0)
  );
  Switch imm_switch_168 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_168_io_y),
    .io_z(imm_switch_168_io_z),
    .io_in0(imm_switch_168_io_in0)
  );
  Switch imm_switch_169 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_169_io_y),
    .io_z(imm_switch_169_io_z),
    .io_in0(imm_switch_169_io_in0)
  );
  Switch imm_switch_170 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_170_io_y),
    .io_z(imm_switch_170_io_z),
    .io_in0(imm_switch_170_io_in0)
  );
  Switch imm_switch_171 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_171_io_y),
    .io_z(imm_switch_171_io_z),
    .io_in0(imm_switch_171_io_in0)
  );
  Switch imm_switch_172 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_172_io_y),
    .io_z(imm_switch_172_io_z),
    .io_in0(imm_switch_172_io_in0)
  );
  Switch imm_switch_173 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_173_io_y),
    .io_z(imm_switch_173_io_z),
    .io_in0(imm_switch_173_io_in0)
  );
  Switch imm_switch_174 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_174_io_y),
    .io_z(imm_switch_174_io_z),
    .io_in0(imm_switch_174_io_in0)
  );
  Switch imm_switch_175 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_175_io_y),
    .io_z(imm_switch_175_io_z),
    .io_in0(imm_switch_175_io_in0)
  );
  Switch imm_switch_176 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_176_io_y),
    .io_z(imm_switch_176_io_z),
    .io_in0(imm_switch_176_io_in0)
  );
  Switch imm_switch_177 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_177_io_y),
    .io_z(imm_switch_177_io_z),
    .io_in0(imm_switch_177_io_in0)
  );
  Switch imm_switch_178 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_178_io_y),
    .io_z(imm_switch_178_io_z),
    .io_in0(imm_switch_178_io_in0)
  );
  Switch imm_switch_179 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_179_io_y),
    .io_z(imm_switch_179_io_z),
    .io_in0(imm_switch_179_io_in0)
  );
  Switch imm_switch_180 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_180_io_y),
    .io_z(imm_switch_180_io_z),
    .io_in0(imm_switch_180_io_in0)
  );
  Switch imm_switch_181 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_181_io_y),
    .io_z(imm_switch_181_io_z),
    .io_in0(imm_switch_181_io_in0)
  );
  Switch imm_switch_182 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_182_io_y),
    .io_z(imm_switch_182_io_z),
    .io_in0(imm_switch_182_io_in0)
  );
  Switch imm_switch_183 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_183_io_y),
    .io_z(imm_switch_183_io_z),
    .io_in0(imm_switch_183_io_in0)
  );
  Switch imm_switch_184 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_184_io_y),
    .io_z(imm_switch_184_io_z),
    .io_in0(imm_switch_184_io_in0)
  );
  Switch imm_switch_185 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_185_io_y),
    .io_z(imm_switch_185_io_z),
    .io_in0(imm_switch_185_io_in0)
  );
  Switch imm_switch_186 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_186_io_y),
    .io_z(imm_switch_186_io_z),
    .io_in0(imm_switch_186_io_in0)
  );
  Switch imm_switch_187 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_187_io_y),
    .io_z(imm_switch_187_io_z),
    .io_in0(imm_switch_187_io_in0)
  );
  Switch imm_switch_188 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_188_io_y),
    .io_z(imm_switch_188_io_z),
    .io_in0(imm_switch_188_io_in0)
  );
  Switch imm_switch_189 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_189_io_y),
    .io_z(imm_switch_189_io_z),
    .io_in0(imm_switch_189_io_in0)
  );
  Switch imm_switch_190 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_190_io_y),
    .io_z(imm_switch_190_io_z),
    .io_in0(imm_switch_190_io_in0)
  );
  Switch imm_switch_191 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_191_io_y),
    .io_z(imm_switch_191_io_z),
    .io_in0(imm_switch_191_io_in0)
  );
  Switch imm_switch_192 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_192_io_y),
    .io_z(imm_switch_192_io_z),
    .io_in0(imm_switch_192_io_in0)
  );
  Switch imm_switch_193 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_193_io_y),
    .io_z(imm_switch_193_io_z),
    .io_in0(imm_switch_193_io_in0)
  );
  Switch imm_switch_194 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_194_io_y),
    .io_z(imm_switch_194_io_z),
    .io_in0(imm_switch_194_io_in0)
  );
  Switch imm_switch_195 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_195_io_y),
    .io_z(imm_switch_195_io_z),
    .io_in0(imm_switch_195_io_in0)
  );
  Switch imm_switch_196 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_196_io_y),
    .io_z(imm_switch_196_io_z),
    .io_in0(imm_switch_196_io_in0)
  );
  Switch imm_switch_197 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_197_io_y),
    .io_z(imm_switch_197_io_z),
    .io_in0(imm_switch_197_io_in0)
  );
  Switch imm_switch_198 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_198_io_y),
    .io_z(imm_switch_198_io_z),
    .io_in0(imm_switch_198_io_in0)
  );
  Switch imm_switch_199 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_199_io_y),
    .io_z(imm_switch_199_io_z),
    .io_in0(imm_switch_199_io_in0)
  );
  Switch imm_switch_200 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_200_io_y),
    .io_z(imm_switch_200_io_z),
    .io_in0(imm_switch_200_io_in0)
  );
  Switch imm_switch_201 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_201_io_y),
    .io_z(imm_switch_201_io_z),
    .io_in0(imm_switch_201_io_in0)
  );
  Switch imm_switch_202 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_202_io_y),
    .io_z(imm_switch_202_io_z),
    .io_in0(imm_switch_202_io_in0)
  );
  Switch imm_switch_203 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_203_io_y),
    .io_z(imm_switch_203_io_z),
    .io_in0(imm_switch_203_io_in0)
  );
  Switch imm_switch_204 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_204_io_y),
    .io_z(imm_switch_204_io_z),
    .io_in0(imm_switch_204_io_in0)
  );
  Switch imm_switch_205 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_205_io_y),
    .io_z(imm_switch_205_io_z),
    .io_in0(imm_switch_205_io_in0)
  );
  Switch imm_switch_206 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_206_io_y),
    .io_z(imm_switch_206_io_z),
    .io_in0(imm_switch_206_io_in0)
  );
  Switch imm_switch_207 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_207_io_y),
    .io_z(imm_switch_207_io_z),
    .io_in0(imm_switch_207_io_in0)
  );
  Switch imm_switch_208 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_208_io_y),
    .io_z(imm_switch_208_io_z),
    .io_in0(imm_switch_208_io_in0)
  );
  Switch imm_switch_209 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_209_io_y),
    .io_z(imm_switch_209_io_z),
    .io_in0(imm_switch_209_io_in0)
  );
  Switch imm_switch_210 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_210_io_y),
    .io_z(imm_switch_210_io_z),
    .io_in0(imm_switch_210_io_in0)
  );
  Switch imm_switch_211 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_211_io_y),
    .io_z(imm_switch_211_io_z),
    .io_in0(imm_switch_211_io_in0)
  );
  Switch imm_switch_212 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_212_io_y),
    .io_z(imm_switch_212_io_z),
    .io_in0(imm_switch_212_io_in0)
  );
  Switch imm_switch_213 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_213_io_y),
    .io_z(imm_switch_213_io_z),
    .io_in0(imm_switch_213_io_in0)
  );
  Switch imm_switch_214 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_214_io_y),
    .io_z(imm_switch_214_io_z),
    .io_in0(imm_switch_214_io_in0)
  );
  Switch imm_switch_215 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_215_io_y),
    .io_z(imm_switch_215_io_z),
    .io_in0(imm_switch_215_io_in0)
  );
  Switch imm_switch_216 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_216_io_y),
    .io_z(imm_switch_216_io_z),
    .io_in0(imm_switch_216_io_in0)
  );
  Switch imm_switch_217 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_217_io_y),
    .io_z(imm_switch_217_io_z),
    .io_in0(imm_switch_217_io_in0)
  );
  Switch imm_switch_218 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_218_io_y),
    .io_z(imm_switch_218_io_z),
    .io_in0(imm_switch_218_io_in0)
  );
  Switch imm_switch_219 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_219_io_y),
    .io_z(imm_switch_219_io_z),
    .io_in0(imm_switch_219_io_in0)
  );
  Switch imm_switch_220 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_220_io_y),
    .io_z(imm_switch_220_io_z),
    .io_in0(imm_switch_220_io_in0)
  );
  Switch imm_switch_221 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_221_io_y),
    .io_z(imm_switch_221_io_z),
    .io_in0(imm_switch_221_io_in0)
  );
  Switch imm_switch_222 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_222_io_y),
    .io_z(imm_switch_222_io_z),
    .io_in0(imm_switch_222_io_in0)
  );
  Switch imm_switch_223 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_223_io_y),
    .io_z(imm_switch_223_io_z),
    .io_in0(imm_switch_223_io_in0)
  );
  Switch imm_switch_224 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_224_io_y),
    .io_z(imm_switch_224_io_z),
    .io_in0(imm_switch_224_io_in0)
  );
  Switch imm_switch_225 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_225_io_y),
    .io_z(imm_switch_225_io_z),
    .io_in0(imm_switch_225_io_in0)
  );
  Switch imm_switch_226 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_226_io_y),
    .io_z(imm_switch_226_io_z),
    .io_in0(imm_switch_226_io_in0)
  );
  Switch imm_switch_227 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_227_io_y),
    .io_z(imm_switch_227_io_z),
    .io_in0(imm_switch_227_io_in0)
  );
  Switch imm_switch_228 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_228_io_y),
    .io_z(imm_switch_228_io_z),
    .io_in0(imm_switch_228_io_in0)
  );
  Switch imm_switch_229 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_229_io_y),
    .io_z(imm_switch_229_io_z),
    .io_in0(imm_switch_229_io_in0)
  );
  Switch imm_switch_230 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_230_io_y),
    .io_z(imm_switch_230_io_z),
    .io_in0(imm_switch_230_io_in0)
  );
  Switch imm_switch_231 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_231_io_y),
    .io_z(imm_switch_231_io_z),
    .io_in0(imm_switch_231_io_in0)
  );
  Switch imm_switch_232 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_232_io_y),
    .io_z(imm_switch_232_io_z),
    .io_in0(imm_switch_232_io_in0)
  );
  Switch imm_switch_233 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_233_io_y),
    .io_z(imm_switch_233_io_z),
    .io_in0(imm_switch_233_io_in0)
  );
  Switch imm_switch_234 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_234_io_y),
    .io_z(imm_switch_234_io_z),
    .io_in0(imm_switch_234_io_in0)
  );
  Switch imm_switch_235 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_235_io_y),
    .io_z(imm_switch_235_io_z),
    .io_in0(imm_switch_235_io_in0)
  );
  Switch imm_switch_236 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_236_io_y),
    .io_z(imm_switch_236_io_z),
    .io_in0(imm_switch_236_io_in0)
  );
  Switch imm_switch_237 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_237_io_y),
    .io_z(imm_switch_237_io_z),
    .io_in0(imm_switch_237_io_in0)
  );
  Switch imm_switch_238 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_238_io_y),
    .io_z(imm_switch_238_io_z),
    .io_in0(imm_switch_238_io_in0)
  );
  Switch imm_switch_239 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_239_io_y),
    .io_z(imm_switch_239_io_z),
    .io_in0(imm_switch_239_io_in0)
  );
  Switch imm_switch_240 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_240_io_y),
    .io_z(imm_switch_240_io_z),
    .io_in0(imm_switch_240_io_in0)
  );
  Switch imm_switch_241 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_241_io_y),
    .io_z(imm_switch_241_io_z),
    .io_in0(imm_switch_241_io_in0)
  );
  Switch imm_switch_242 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_242_io_y),
    .io_z(imm_switch_242_io_z),
    .io_in0(imm_switch_242_io_in0)
  );
  Switch imm_switch_243 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_243_io_y),
    .io_z(imm_switch_243_io_z),
    .io_in0(imm_switch_243_io_in0)
  );
  Switch imm_switch_244 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_244_io_y),
    .io_z(imm_switch_244_io_z),
    .io_in0(imm_switch_244_io_in0)
  );
  Switch imm_switch_245 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_245_io_y),
    .io_z(imm_switch_245_io_z),
    .io_in0(imm_switch_245_io_in0)
  );
  Switch imm_switch_246 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_246_io_y),
    .io_z(imm_switch_246_io_z),
    .io_in0(imm_switch_246_io_in0)
  );
  Switch imm_switch_247 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_247_io_y),
    .io_z(imm_switch_247_io_z),
    .io_in0(imm_switch_247_io_in0)
  );
  Switch imm_switch_248 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_248_io_y),
    .io_z(imm_switch_248_io_z),
    .io_in0(imm_switch_248_io_in0)
  );
  Switch imm_switch_249 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_249_io_y),
    .io_z(imm_switch_249_io_z),
    .io_in0(imm_switch_249_io_in0)
  );
  Switch imm_switch_250 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_250_io_y),
    .io_z(imm_switch_250_io_z),
    .io_in0(imm_switch_250_io_in0)
  );
  Switch imm_switch_251 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_251_io_y),
    .io_z(imm_switch_251_io_z),
    .io_in0(imm_switch_251_io_in0)
  );
  Switch imm_switch_252 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_252_io_y),
    .io_z(imm_switch_252_io_z),
    .io_in0(imm_switch_252_io_in0)
  );
  Switch imm_switch_253 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_253_io_y),
    .io_z(imm_switch_253_io_z),
    .io_in0(imm_switch_253_io_in0)
  );
  Switch imm_switch_254 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_254_io_y),
    .io_z(imm_switch_254_io_z),
    .io_in0(imm_switch_254_io_in0)
  );
  Switch imm_switch_255 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_255_io_y),
    .io_z(imm_switch_255_io_z),
    .io_in0(imm_switch_255_io_in0)
  );
  Switch imm_switch_256 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_256_io_y),
    .io_z(imm_switch_256_io_z),
    .io_in0(imm_switch_256_io_in0)
  );
  Switch imm_switch_257 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_257_io_y),
    .io_z(imm_switch_257_io_z),
    .io_in0(imm_switch_257_io_in0)
  );
  Switch imm_switch_258 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_258_io_y),
    .io_z(imm_switch_258_io_z),
    .io_in0(imm_switch_258_io_in0)
  );
  Switch imm_switch_259 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_259_io_y),
    .io_z(imm_switch_259_io_z),
    .io_in0(imm_switch_259_io_in0)
  );
  Switch imm_switch_260 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_260_io_y),
    .io_z(imm_switch_260_io_z),
    .io_in0(imm_switch_260_io_in0)
  );
  Switch imm_switch_261 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_261_io_y),
    .io_z(imm_switch_261_io_z),
    .io_in0(imm_switch_261_io_in0)
  );
  Switch imm_switch_262 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_262_io_y),
    .io_z(imm_switch_262_io_z),
    .io_in0(imm_switch_262_io_in0)
  );
  Switch imm_switch_263 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_263_io_y),
    .io_z(imm_switch_263_io_z),
    .io_in0(imm_switch_263_io_in0)
  );
  Switch imm_switch_264 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_264_io_y),
    .io_z(imm_switch_264_io_z),
    .io_in0(imm_switch_264_io_in0)
  );
  Switch imm_switch_265 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_265_io_y),
    .io_z(imm_switch_265_io_z),
    .io_in0(imm_switch_265_io_in0)
  );
  Switch imm_switch_266 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_266_io_y),
    .io_z(imm_switch_266_io_z),
    .io_in0(imm_switch_266_io_in0)
  );
  Switch imm_switch_267 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_267_io_y),
    .io_z(imm_switch_267_io_z),
    .io_in0(imm_switch_267_io_in0)
  );
  Switch imm_switch_268 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_268_io_y),
    .io_z(imm_switch_268_io_z),
    .io_in0(imm_switch_268_io_in0)
  );
  Switch imm_switch_269 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_269_io_y),
    .io_z(imm_switch_269_io_z),
    .io_in0(imm_switch_269_io_in0)
  );
  Switch imm_switch_270 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_270_io_y),
    .io_z(imm_switch_270_io_z),
    .io_in0(imm_switch_270_io_in0)
  );
  Switch imm_switch_271 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_271_io_y),
    .io_z(imm_switch_271_io_z),
    .io_in0(imm_switch_271_io_in0)
  );
  Switch imm_switch_272 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_272_io_y),
    .io_z(imm_switch_272_io_z),
    .io_in0(imm_switch_272_io_in0)
  );
  Switch imm_switch_273 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_273_io_y),
    .io_z(imm_switch_273_io_z),
    .io_in0(imm_switch_273_io_in0)
  );
  Switch imm_switch_274 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_274_io_y),
    .io_z(imm_switch_274_io_z),
    .io_in0(imm_switch_274_io_in0)
  );
  Switch imm_switch_275 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_275_io_y),
    .io_z(imm_switch_275_io_z),
    .io_in0(imm_switch_275_io_in0)
  );
  Switch imm_switch_276 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_276_io_y),
    .io_z(imm_switch_276_io_z),
    .io_in0(imm_switch_276_io_in0)
  );
  Switch imm_switch_277 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_277_io_y),
    .io_z(imm_switch_277_io_z),
    .io_in0(imm_switch_277_io_in0)
  );
  Switch imm_switch_278 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_278_io_y),
    .io_z(imm_switch_278_io_z),
    .io_in0(imm_switch_278_io_in0)
  );
  Switch imm_switch_279 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_279_io_y),
    .io_z(imm_switch_279_io_z),
    .io_in0(imm_switch_279_io_in0)
  );
  Switch imm_switch_280 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_280_io_y),
    .io_z(imm_switch_280_io_z),
    .io_in0(imm_switch_280_io_in0)
  );
  Switch imm_switch_281 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_281_io_y),
    .io_z(imm_switch_281_io_z),
    .io_in0(imm_switch_281_io_in0)
  );
  Switch imm_switch_282 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_282_io_y),
    .io_z(imm_switch_282_io_z),
    .io_in0(imm_switch_282_io_in0)
  );
  Switch imm_switch_283 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_283_io_y),
    .io_z(imm_switch_283_io_z),
    .io_in0(imm_switch_283_io_in0)
  );
  Switch imm_switch_284 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_284_io_y),
    .io_z(imm_switch_284_io_z),
    .io_in0(imm_switch_284_io_in0)
  );
  Switch imm_switch_285 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_285_io_y),
    .io_z(imm_switch_285_io_z),
    .io_in0(imm_switch_285_io_in0)
  );
  Switch imm_switch_286 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_286_io_y),
    .io_z(imm_switch_286_io_z),
    .io_in0(imm_switch_286_io_in0)
  );
  Switch imm_switch_287 ( // @[Benes.scala 109:30]
    .io_y(imm_switch_287_io_y),
    .io_z(imm_switch_287_io_z),
    .io_in0(imm_switch_287_io_in0)
  );
  assign io_o_dist_bus2_0 = reset ? 16'h0 : w_dist_bus_0; // @[Benes.scala 86:24]
  assign io_o_dist_bus2_1 = reset ? 16'h0 : w_dist_bus_1; // @[Benes.scala 86:24]
  assign io_o_dist_bus2_2 = reset ? 16'h0 : w_dist_bus_2; // @[Benes.scala 86:24]
  assign io_o_dist_bus2_3 = reset ? 16'h0 : w_dist_bus_3; // @[Benes.scala 86:24]
  assign io_o_dist_bus2_4 = reset ? 16'h0 : w_dist_bus_4; // @[Benes.scala 86:24]
  assign io_o_dist_bus2_5 = reset ? 16'h0 : w_dist_bus_5; // @[Benes.scala 86:24]
  assign io_o_dist_bus2_6 = reset ? 16'h0 : w_dist_bus_6; // @[Benes.scala 86:24]
  assign io_o_dist_bus2_7 = reset ? 16'h0 : w_dist_bus_7; // @[Benes.scala 86:24]
  assign io_o_dist_bus2_8 = reset ? 16'h0 : w_dist_bus_8; // @[Benes.scala 86:24]
  assign io_o_dist_bus2_9 = reset ? 16'h0 : w_dist_bus_9; // @[Benes.scala 86:24]
  assign io_o_dist_bus2_10 = reset ? 16'h0 : w_dist_bus_10; // @[Benes.scala 86:24]
  assign io_o_dist_bus2_11 = reset ? 16'h0 : w_dist_bus_11; // @[Benes.scala 86:24]
  assign io_o_dist_bus2_12 = reset ? 16'h0 : w_dist_bus_12; // @[Benes.scala 86:24]
  assign io_o_dist_bus2_13 = reset ? 16'h0 : w_dist_bus_13; // @[Benes.scala 86:24]
  assign io_o_dist_bus2_14 = reset ? 16'h0 : w_dist_bus_14; // @[Benes.scala 86:24]
  assign io_o_dist_bus2_15 = reset ? 16'h0 : w_dist_bus_15; // @[Benes.scala 86:24]
  assign io_o_dist_bus2_16 = reset ? 16'h0 : w_dist_bus_16; // @[Benes.scala 86:24]
  assign io_o_dist_bus2_17 = reset ? 16'h0 : w_dist_bus_17; // @[Benes.scala 86:24]
  assign io_o_dist_bus2_18 = reset ? 16'h0 : w_dist_bus_18; // @[Benes.scala 86:24]
  assign io_o_dist_bus2_19 = reset ? 16'h0 : w_dist_bus_19; // @[Benes.scala 86:24]
  assign io_o_dist_bus2_20 = reset ? 16'h0 : w_dist_bus_20; // @[Benes.scala 86:24]
  assign io_o_dist_bus2_21 = reset ? 16'h0 : w_dist_bus_21; // @[Benes.scala 86:24]
  assign io_o_dist_bus2_22 = reset ? 16'h0 : w_dist_bus_22; // @[Benes.scala 86:24]
  assign io_o_dist_bus2_23 = reset ? 16'h0 : w_dist_bus_23; // @[Benes.scala 86:24]
  assign io_o_dist_bus2_24 = reset ? 16'h0 : w_dist_bus_24; // @[Benes.scala 86:24]
  assign io_o_dist_bus2_25 = reset ? 16'h0 : w_dist_bus_25; // @[Benes.scala 86:24]
  assign io_o_dist_bus2_26 = reset ? 16'h0 : w_dist_bus_26; // @[Benes.scala 86:24]
  assign io_o_dist_bus2_27 = reset ? 16'h0 : w_dist_bus_27; // @[Benes.scala 86:24]
  assign io_o_dist_bus2_28 = reset ? 16'h0 : w_dist_bus_28; // @[Benes.scala 86:24]
  assign io_o_dist_bus2_29 = reset ? 16'h0 : w_dist_bus_29; // @[Benes.scala 86:24]
  assign io_o_dist_bus2_30 = reset ? 16'h0 : w_dist_bus_30; // @[Benes.scala 86:24]
  assign io_o_dist_bus2_31 = reset ? 16'h0 : w_dist_bus_31; // @[Benes.scala 86:24]
  assign in_switch_io_in = r_data_bus_ff_0; // @[Benes.scala 91:21]
  assign in_switch_1_io_in = r_data_bus_ff_1; // @[Benes.scala 91:21]
  assign in_switch_2_io_in = r_data_bus_ff_2; // @[Benes.scala 91:21]
  assign in_switch_3_io_in = r_data_bus_ff_3; // @[Benes.scala 91:21]
  assign in_switch_4_io_in = r_data_bus_ff_4; // @[Benes.scala 91:21]
  assign in_switch_5_io_in = r_data_bus_ff_5; // @[Benes.scala 91:21]
  assign in_switch_6_io_in = r_data_bus_ff_6; // @[Benes.scala 91:21]
  assign in_switch_7_io_in = r_data_bus_ff_7; // @[Benes.scala 91:21]
  assign in_switch_8_io_in = r_data_bus_ff_8; // @[Benes.scala 91:21]
  assign in_switch_9_io_in = r_data_bus_ff_9; // @[Benes.scala 91:21]
  assign in_switch_10_io_in = r_data_bus_ff_10; // @[Benes.scala 91:21]
  assign in_switch_11_io_in = r_data_bus_ff_11; // @[Benes.scala 91:21]
  assign in_switch_12_io_in = r_data_bus_ff_12; // @[Benes.scala 91:21]
  assign in_switch_13_io_in = r_data_bus_ff_13; // @[Benes.scala 91:21]
  assign in_switch_14_io_in = r_data_bus_ff_14; // @[Benes.scala 91:21]
  assign in_switch_15_io_in = r_data_bus_ff_15; // @[Benes.scala 91:21]
  assign in_switch_16_io_in = r_data_bus_ff_16; // @[Benes.scala 91:21]
  assign in_switch_17_io_in = r_data_bus_ff_17; // @[Benes.scala 91:21]
  assign in_switch_18_io_in = r_data_bus_ff_18; // @[Benes.scala 91:21]
  assign in_switch_19_io_in = r_data_bus_ff_19; // @[Benes.scala 91:21]
  assign in_switch_20_io_in = r_data_bus_ff_20; // @[Benes.scala 91:21]
  assign in_switch_21_io_in = r_data_bus_ff_21; // @[Benes.scala 91:21]
  assign in_switch_22_io_in = r_data_bus_ff_22; // @[Benes.scala 91:21]
  assign in_switch_23_io_in = r_data_bus_ff_23; // @[Benes.scala 91:21]
  assign in_switch_24_io_in = r_data_bus_ff_24; // @[Benes.scala 91:21]
  assign in_switch_25_io_in = r_data_bus_ff_25; // @[Benes.scala 91:21]
  assign in_switch_26_io_in = r_data_bus_ff_26; // @[Benes.scala 91:21]
  assign in_switch_27_io_in = r_data_bus_ff_27; // @[Benes.scala 91:21]
  assign in_switch_28_io_in = r_data_bus_ff_28; // @[Benes.scala 91:21]
  assign in_switch_29_io_in = r_data_bus_ff_29; // @[Benes.scala 91:21]
  assign in_switch_30_io_in = r_data_bus_ff_30; // @[Benes.scala 91:21]
  assign in_switch_31_io_in = r_data_bus_ff_31; // @[Benes.scala 91:21]
  assign out_switch_io_in0 = w_internal_18; // @[Benes.scala 100:23]
  assign out_switch_1_io_in0 = w_internal_38; // @[Benes.scala 100:23]
  assign out_switch_2_io_in0 = w_internal_58; // @[Benes.scala 100:23]
  assign out_switch_3_io_in0 = w_internal_78; // @[Benes.scala 100:23]
  assign out_switch_4_io_in0 = w_internal_98; // @[Benes.scala 100:23]
  assign out_switch_5_io_in0 = w_internal_118; // @[Benes.scala 100:23]
  assign out_switch_6_io_in0 = w_internal_138; // @[Benes.scala 100:23]
  assign out_switch_7_io_in0 = w_internal_158; // @[Benes.scala 100:23]
  assign out_switch_8_io_in0 = w_internal_178; // @[Benes.scala 100:23]
  assign out_switch_9_io_in0 = w_internal_198; // @[Benes.scala 100:23]
  assign out_switch_10_io_in0 = w_internal_218; // @[Benes.scala 100:23]
  assign out_switch_11_io_in0 = w_internal_238; // @[Benes.scala 100:23]
  assign out_switch_12_io_in0 = w_internal_258; // @[Benes.scala 100:23]
  assign out_switch_13_io_in0 = w_internal_278; // @[Benes.scala 100:23]
  assign out_switch_14_io_in0 = w_internal_298; // @[Benes.scala 100:23]
  assign out_switch_15_io_in0 = w_internal_318; // @[Benes.scala 100:23]
  assign out_switch_16_io_in0 = w_internal_338; // @[Benes.scala 100:23]
  assign out_switch_17_io_in0 = w_internal_358; // @[Benes.scala 100:23]
  assign out_switch_18_io_in0 = w_internal_378; // @[Benes.scala 100:23]
  assign out_switch_19_io_in0 = w_internal_398; // @[Benes.scala 100:23]
  assign out_switch_20_io_in0 = w_internal_418; // @[Benes.scala 100:23]
  assign out_switch_21_io_in0 = w_internal_438; // @[Benes.scala 100:23]
  assign out_switch_22_io_in0 = w_internal_458; // @[Benes.scala 100:23]
  assign out_switch_23_io_in0 = w_internal_478; // @[Benes.scala 100:23]
  assign out_switch_24_io_in0 = w_internal_498; // @[Benes.scala 100:23]
  assign out_switch_25_io_in0 = w_internal_518; // @[Benes.scala 100:23]
  assign out_switch_26_io_in0 = w_internal_538; // @[Benes.scala 100:23]
  assign out_switch_27_io_in0 = w_internal_558; // @[Benes.scala 100:23]
  assign out_switch_28_io_in0 = w_internal_578; // @[Benes.scala 100:23]
  assign out_switch_29_io_in0 = w_internal_598; // @[Benes.scala 100:23]
  assign out_switch_30_io_in0 = w_internal_618; // @[Benes.scala 100:23]
  assign out_switch_31_io_in0 = w_internal_638; // @[Benes.scala 100:23]
  assign imm_switch_io_in0 = w_internal_0; // @[Benes.scala 110:25]
  assign imm_switch_1_io_in0 = w_internal_2; // @[Benes.scala 110:25]
  assign imm_switch_2_io_in0 = w_internal_4; // @[Benes.scala 110:25]
  assign imm_switch_3_io_in0 = w_internal_6; // @[Benes.scala 110:25]
  assign imm_switch_4_io_in0 = w_internal_8; // @[Benes.scala 110:25]
  assign imm_switch_5_io_in0 = w_internal_10; // @[Benes.scala 110:25]
  assign imm_switch_6_io_in0 = w_internal_12; // @[Benes.scala 110:25]
  assign imm_switch_7_io_in0 = w_internal_14; // @[Benes.scala 110:25]
  assign imm_switch_8_io_in0 = w_internal_16; // @[Benes.scala 110:25]
  assign imm_switch_9_io_in0 = w_internal_20; // @[Benes.scala 110:25]
  assign imm_switch_10_io_in0 = w_internal_22; // @[Benes.scala 110:25]
  assign imm_switch_11_io_in0 = w_internal_24; // @[Benes.scala 110:25]
  assign imm_switch_12_io_in0 = w_internal_26; // @[Benes.scala 110:25]
  assign imm_switch_13_io_in0 = w_internal_28; // @[Benes.scala 110:25]
  assign imm_switch_14_io_in0 = w_internal_30; // @[Benes.scala 110:25]
  assign imm_switch_15_io_in0 = w_internal_32; // @[Benes.scala 110:25]
  assign imm_switch_16_io_in0 = w_internal_34; // @[Benes.scala 110:25]
  assign imm_switch_17_io_in0 = w_internal_36; // @[Benes.scala 110:25]
  assign imm_switch_18_io_in0 = w_internal_40; // @[Benes.scala 110:25]
  assign imm_switch_19_io_in0 = w_internal_42; // @[Benes.scala 110:25]
  assign imm_switch_20_io_in0 = w_internal_44; // @[Benes.scala 110:25]
  assign imm_switch_21_io_in0 = w_internal_46; // @[Benes.scala 110:25]
  assign imm_switch_22_io_in0 = w_internal_48; // @[Benes.scala 110:25]
  assign imm_switch_23_io_in0 = w_internal_50; // @[Benes.scala 110:25]
  assign imm_switch_24_io_in0 = w_internal_52; // @[Benes.scala 110:25]
  assign imm_switch_25_io_in0 = w_internal_54; // @[Benes.scala 110:25]
  assign imm_switch_26_io_in0 = w_internal_56; // @[Benes.scala 110:25]
  assign imm_switch_27_io_in0 = w_internal_60; // @[Benes.scala 110:25]
  assign imm_switch_28_io_in0 = w_internal_62; // @[Benes.scala 110:25]
  assign imm_switch_29_io_in0 = w_internal_64; // @[Benes.scala 110:25]
  assign imm_switch_30_io_in0 = w_internal_66; // @[Benes.scala 110:25]
  assign imm_switch_31_io_in0 = w_internal_68; // @[Benes.scala 110:25]
  assign imm_switch_32_io_in0 = w_internal_70; // @[Benes.scala 110:25]
  assign imm_switch_33_io_in0 = w_internal_72; // @[Benes.scala 110:25]
  assign imm_switch_34_io_in0 = w_internal_74; // @[Benes.scala 110:25]
  assign imm_switch_35_io_in0 = w_internal_76; // @[Benes.scala 110:25]
  assign imm_switch_36_io_in0 = w_internal_80; // @[Benes.scala 110:25]
  assign imm_switch_37_io_in0 = w_internal_82; // @[Benes.scala 110:25]
  assign imm_switch_38_io_in0 = w_internal_84; // @[Benes.scala 110:25]
  assign imm_switch_39_io_in0 = w_internal_86; // @[Benes.scala 110:25]
  assign imm_switch_40_io_in0 = w_internal_88; // @[Benes.scala 110:25]
  assign imm_switch_41_io_in0 = w_internal_90; // @[Benes.scala 110:25]
  assign imm_switch_42_io_in0 = w_internal_92; // @[Benes.scala 110:25]
  assign imm_switch_43_io_in0 = w_internal_94; // @[Benes.scala 110:25]
  assign imm_switch_44_io_in0 = w_internal_96; // @[Benes.scala 110:25]
  assign imm_switch_45_io_in0 = w_internal_100; // @[Benes.scala 110:25]
  assign imm_switch_46_io_in0 = w_internal_102; // @[Benes.scala 110:25]
  assign imm_switch_47_io_in0 = w_internal_104; // @[Benes.scala 110:25]
  assign imm_switch_48_io_in0 = w_internal_106; // @[Benes.scala 110:25]
  assign imm_switch_49_io_in0 = w_internal_108; // @[Benes.scala 110:25]
  assign imm_switch_50_io_in0 = w_internal_110; // @[Benes.scala 110:25]
  assign imm_switch_51_io_in0 = w_internal_112; // @[Benes.scala 110:25]
  assign imm_switch_52_io_in0 = w_internal_114; // @[Benes.scala 110:25]
  assign imm_switch_53_io_in0 = w_internal_116; // @[Benes.scala 110:25]
  assign imm_switch_54_io_in0 = w_internal_120; // @[Benes.scala 110:25]
  assign imm_switch_55_io_in0 = w_internal_122; // @[Benes.scala 110:25]
  assign imm_switch_56_io_in0 = w_internal_124; // @[Benes.scala 110:25]
  assign imm_switch_57_io_in0 = w_internal_126; // @[Benes.scala 110:25]
  assign imm_switch_58_io_in0 = w_internal_128; // @[Benes.scala 110:25]
  assign imm_switch_59_io_in0 = w_internal_130; // @[Benes.scala 110:25]
  assign imm_switch_60_io_in0 = w_internal_132; // @[Benes.scala 110:25]
  assign imm_switch_61_io_in0 = w_internal_134; // @[Benes.scala 110:25]
  assign imm_switch_62_io_in0 = w_internal_136; // @[Benes.scala 110:25]
  assign imm_switch_63_io_in0 = w_internal_140; // @[Benes.scala 110:25]
  assign imm_switch_64_io_in0 = w_internal_142; // @[Benes.scala 110:25]
  assign imm_switch_65_io_in0 = w_internal_144; // @[Benes.scala 110:25]
  assign imm_switch_66_io_in0 = w_internal_146; // @[Benes.scala 110:25]
  assign imm_switch_67_io_in0 = w_internal_148; // @[Benes.scala 110:25]
  assign imm_switch_68_io_in0 = w_internal_150; // @[Benes.scala 110:25]
  assign imm_switch_69_io_in0 = w_internal_152; // @[Benes.scala 110:25]
  assign imm_switch_70_io_in0 = w_internal_154; // @[Benes.scala 110:25]
  assign imm_switch_71_io_in0 = w_internal_156; // @[Benes.scala 110:25]
  assign imm_switch_72_io_in0 = w_internal_160; // @[Benes.scala 110:25]
  assign imm_switch_73_io_in0 = w_internal_162; // @[Benes.scala 110:25]
  assign imm_switch_74_io_in0 = w_internal_164; // @[Benes.scala 110:25]
  assign imm_switch_75_io_in0 = w_internal_166; // @[Benes.scala 110:25]
  assign imm_switch_76_io_in0 = w_internal_168; // @[Benes.scala 110:25]
  assign imm_switch_77_io_in0 = w_internal_170; // @[Benes.scala 110:25]
  assign imm_switch_78_io_in0 = w_internal_172; // @[Benes.scala 110:25]
  assign imm_switch_79_io_in0 = w_internal_174; // @[Benes.scala 110:25]
  assign imm_switch_80_io_in0 = w_internal_176; // @[Benes.scala 110:25]
  assign imm_switch_81_io_in0 = w_internal_180; // @[Benes.scala 110:25]
  assign imm_switch_82_io_in0 = w_internal_182; // @[Benes.scala 110:25]
  assign imm_switch_83_io_in0 = w_internal_184; // @[Benes.scala 110:25]
  assign imm_switch_84_io_in0 = w_internal_186; // @[Benes.scala 110:25]
  assign imm_switch_85_io_in0 = w_internal_188; // @[Benes.scala 110:25]
  assign imm_switch_86_io_in0 = w_internal_190; // @[Benes.scala 110:25]
  assign imm_switch_87_io_in0 = w_internal_192; // @[Benes.scala 110:25]
  assign imm_switch_88_io_in0 = w_internal_194; // @[Benes.scala 110:25]
  assign imm_switch_89_io_in0 = w_internal_196; // @[Benes.scala 110:25]
  assign imm_switch_90_io_in0 = w_internal_200; // @[Benes.scala 110:25]
  assign imm_switch_91_io_in0 = w_internal_202; // @[Benes.scala 110:25]
  assign imm_switch_92_io_in0 = w_internal_204; // @[Benes.scala 110:25]
  assign imm_switch_93_io_in0 = w_internal_206; // @[Benes.scala 110:25]
  assign imm_switch_94_io_in0 = w_internal_208; // @[Benes.scala 110:25]
  assign imm_switch_95_io_in0 = w_internal_210; // @[Benes.scala 110:25]
  assign imm_switch_96_io_in0 = w_internal_212; // @[Benes.scala 110:25]
  assign imm_switch_97_io_in0 = w_internal_214; // @[Benes.scala 110:25]
  assign imm_switch_98_io_in0 = w_internal_216; // @[Benes.scala 110:25]
  assign imm_switch_99_io_in0 = w_internal_220; // @[Benes.scala 110:25]
  assign imm_switch_100_io_in0 = w_internal_222; // @[Benes.scala 110:25]
  assign imm_switch_101_io_in0 = w_internal_224; // @[Benes.scala 110:25]
  assign imm_switch_102_io_in0 = w_internal_226; // @[Benes.scala 110:25]
  assign imm_switch_103_io_in0 = w_internal_228; // @[Benes.scala 110:25]
  assign imm_switch_104_io_in0 = w_internal_230; // @[Benes.scala 110:25]
  assign imm_switch_105_io_in0 = w_internal_232; // @[Benes.scala 110:25]
  assign imm_switch_106_io_in0 = w_internal_234; // @[Benes.scala 110:25]
  assign imm_switch_107_io_in0 = w_internal_236; // @[Benes.scala 110:25]
  assign imm_switch_108_io_in0 = w_internal_240; // @[Benes.scala 110:25]
  assign imm_switch_109_io_in0 = w_internal_242; // @[Benes.scala 110:25]
  assign imm_switch_110_io_in0 = w_internal_244; // @[Benes.scala 110:25]
  assign imm_switch_111_io_in0 = w_internal_246; // @[Benes.scala 110:25]
  assign imm_switch_112_io_in0 = w_internal_248; // @[Benes.scala 110:25]
  assign imm_switch_113_io_in0 = w_internal_250; // @[Benes.scala 110:25]
  assign imm_switch_114_io_in0 = w_internal_252; // @[Benes.scala 110:25]
  assign imm_switch_115_io_in0 = w_internal_254; // @[Benes.scala 110:25]
  assign imm_switch_116_io_in0 = w_internal_256; // @[Benes.scala 110:25]
  assign imm_switch_117_io_in0 = w_internal_260; // @[Benes.scala 110:25]
  assign imm_switch_118_io_in0 = w_internal_262; // @[Benes.scala 110:25]
  assign imm_switch_119_io_in0 = w_internal_264; // @[Benes.scala 110:25]
  assign imm_switch_120_io_in0 = w_internal_266; // @[Benes.scala 110:25]
  assign imm_switch_121_io_in0 = w_internal_268; // @[Benes.scala 110:25]
  assign imm_switch_122_io_in0 = w_internal_270; // @[Benes.scala 110:25]
  assign imm_switch_123_io_in0 = w_internal_272; // @[Benes.scala 110:25]
  assign imm_switch_124_io_in0 = w_internal_274; // @[Benes.scala 110:25]
  assign imm_switch_125_io_in0 = w_internal_276; // @[Benes.scala 110:25]
  assign imm_switch_126_io_in0 = w_internal_280; // @[Benes.scala 110:25]
  assign imm_switch_127_io_in0 = w_internal_282; // @[Benes.scala 110:25]
  assign imm_switch_128_io_in0 = w_internal_284; // @[Benes.scala 110:25]
  assign imm_switch_129_io_in0 = w_internal_286; // @[Benes.scala 110:25]
  assign imm_switch_130_io_in0 = w_internal_288; // @[Benes.scala 110:25]
  assign imm_switch_131_io_in0 = w_internal_290; // @[Benes.scala 110:25]
  assign imm_switch_132_io_in0 = w_internal_292; // @[Benes.scala 110:25]
  assign imm_switch_133_io_in0 = w_internal_294; // @[Benes.scala 110:25]
  assign imm_switch_134_io_in0 = w_internal_296; // @[Benes.scala 110:25]
  assign imm_switch_135_io_in0 = w_internal_300; // @[Benes.scala 110:25]
  assign imm_switch_136_io_in0 = w_internal_302; // @[Benes.scala 110:25]
  assign imm_switch_137_io_in0 = w_internal_304; // @[Benes.scala 110:25]
  assign imm_switch_138_io_in0 = w_internal_306; // @[Benes.scala 110:25]
  assign imm_switch_139_io_in0 = w_internal_308; // @[Benes.scala 110:25]
  assign imm_switch_140_io_in0 = w_internal_310; // @[Benes.scala 110:25]
  assign imm_switch_141_io_in0 = w_internal_312; // @[Benes.scala 110:25]
  assign imm_switch_142_io_in0 = w_internal_314; // @[Benes.scala 110:25]
  assign imm_switch_143_io_in0 = w_internal_316; // @[Benes.scala 110:25]
  assign imm_switch_144_io_in0 = w_internal_320; // @[Benes.scala 110:25]
  assign imm_switch_145_io_in0 = w_internal_322; // @[Benes.scala 110:25]
  assign imm_switch_146_io_in0 = w_internal_324; // @[Benes.scala 110:25]
  assign imm_switch_147_io_in0 = w_internal_326; // @[Benes.scala 110:25]
  assign imm_switch_148_io_in0 = w_internal_328; // @[Benes.scala 110:25]
  assign imm_switch_149_io_in0 = w_internal_330; // @[Benes.scala 110:25]
  assign imm_switch_150_io_in0 = w_internal_332; // @[Benes.scala 110:25]
  assign imm_switch_151_io_in0 = w_internal_334; // @[Benes.scala 110:25]
  assign imm_switch_152_io_in0 = w_internal_336; // @[Benes.scala 110:25]
  assign imm_switch_153_io_in0 = w_internal_340; // @[Benes.scala 110:25]
  assign imm_switch_154_io_in0 = w_internal_342; // @[Benes.scala 110:25]
  assign imm_switch_155_io_in0 = w_internal_344; // @[Benes.scala 110:25]
  assign imm_switch_156_io_in0 = w_internal_346; // @[Benes.scala 110:25]
  assign imm_switch_157_io_in0 = w_internal_348; // @[Benes.scala 110:25]
  assign imm_switch_158_io_in0 = w_internal_350; // @[Benes.scala 110:25]
  assign imm_switch_159_io_in0 = w_internal_352; // @[Benes.scala 110:25]
  assign imm_switch_160_io_in0 = w_internal_354; // @[Benes.scala 110:25]
  assign imm_switch_161_io_in0 = w_internal_356; // @[Benes.scala 110:25]
  assign imm_switch_162_io_in0 = w_internal_360; // @[Benes.scala 110:25]
  assign imm_switch_163_io_in0 = w_internal_362; // @[Benes.scala 110:25]
  assign imm_switch_164_io_in0 = w_internal_364; // @[Benes.scala 110:25]
  assign imm_switch_165_io_in0 = w_internal_366; // @[Benes.scala 110:25]
  assign imm_switch_166_io_in0 = w_internal_368; // @[Benes.scala 110:25]
  assign imm_switch_167_io_in0 = w_internal_370; // @[Benes.scala 110:25]
  assign imm_switch_168_io_in0 = w_internal_372; // @[Benes.scala 110:25]
  assign imm_switch_169_io_in0 = w_internal_374; // @[Benes.scala 110:25]
  assign imm_switch_170_io_in0 = w_internal_376; // @[Benes.scala 110:25]
  assign imm_switch_171_io_in0 = w_internal_380; // @[Benes.scala 110:25]
  assign imm_switch_172_io_in0 = w_internal_382; // @[Benes.scala 110:25]
  assign imm_switch_173_io_in0 = w_internal_384; // @[Benes.scala 110:25]
  assign imm_switch_174_io_in0 = w_internal_386; // @[Benes.scala 110:25]
  assign imm_switch_175_io_in0 = w_internal_388; // @[Benes.scala 110:25]
  assign imm_switch_176_io_in0 = w_internal_390; // @[Benes.scala 110:25]
  assign imm_switch_177_io_in0 = w_internal_392; // @[Benes.scala 110:25]
  assign imm_switch_178_io_in0 = w_internal_394; // @[Benes.scala 110:25]
  assign imm_switch_179_io_in0 = w_internal_396; // @[Benes.scala 110:25]
  assign imm_switch_180_io_in0 = w_internal_400; // @[Benes.scala 110:25]
  assign imm_switch_181_io_in0 = w_internal_402; // @[Benes.scala 110:25]
  assign imm_switch_182_io_in0 = w_internal_404; // @[Benes.scala 110:25]
  assign imm_switch_183_io_in0 = w_internal_406; // @[Benes.scala 110:25]
  assign imm_switch_184_io_in0 = w_internal_408; // @[Benes.scala 110:25]
  assign imm_switch_185_io_in0 = w_internal_410; // @[Benes.scala 110:25]
  assign imm_switch_186_io_in0 = w_internal_412; // @[Benes.scala 110:25]
  assign imm_switch_187_io_in0 = w_internal_414; // @[Benes.scala 110:25]
  assign imm_switch_188_io_in0 = w_internal_416; // @[Benes.scala 110:25]
  assign imm_switch_189_io_in0 = w_internal_420; // @[Benes.scala 110:25]
  assign imm_switch_190_io_in0 = w_internal_422; // @[Benes.scala 110:25]
  assign imm_switch_191_io_in0 = w_internal_424; // @[Benes.scala 110:25]
  assign imm_switch_192_io_in0 = w_internal_426; // @[Benes.scala 110:25]
  assign imm_switch_193_io_in0 = w_internal_428; // @[Benes.scala 110:25]
  assign imm_switch_194_io_in0 = w_internal_430; // @[Benes.scala 110:25]
  assign imm_switch_195_io_in0 = w_internal_432; // @[Benes.scala 110:25]
  assign imm_switch_196_io_in0 = w_internal_434; // @[Benes.scala 110:25]
  assign imm_switch_197_io_in0 = w_internal_436; // @[Benes.scala 110:25]
  assign imm_switch_198_io_in0 = w_internal_440; // @[Benes.scala 110:25]
  assign imm_switch_199_io_in0 = w_internal_442; // @[Benes.scala 110:25]
  assign imm_switch_200_io_in0 = w_internal_444; // @[Benes.scala 110:25]
  assign imm_switch_201_io_in0 = w_internal_446; // @[Benes.scala 110:25]
  assign imm_switch_202_io_in0 = w_internal_448; // @[Benes.scala 110:25]
  assign imm_switch_203_io_in0 = w_internal_450; // @[Benes.scala 110:25]
  assign imm_switch_204_io_in0 = w_internal_452; // @[Benes.scala 110:25]
  assign imm_switch_205_io_in0 = w_internal_454; // @[Benes.scala 110:25]
  assign imm_switch_206_io_in0 = w_internal_456; // @[Benes.scala 110:25]
  assign imm_switch_207_io_in0 = w_internal_460; // @[Benes.scala 110:25]
  assign imm_switch_208_io_in0 = w_internal_462; // @[Benes.scala 110:25]
  assign imm_switch_209_io_in0 = w_internal_464; // @[Benes.scala 110:25]
  assign imm_switch_210_io_in0 = w_internal_466; // @[Benes.scala 110:25]
  assign imm_switch_211_io_in0 = w_internal_468; // @[Benes.scala 110:25]
  assign imm_switch_212_io_in0 = w_internal_470; // @[Benes.scala 110:25]
  assign imm_switch_213_io_in0 = w_internal_472; // @[Benes.scala 110:25]
  assign imm_switch_214_io_in0 = w_internal_474; // @[Benes.scala 110:25]
  assign imm_switch_215_io_in0 = w_internal_476; // @[Benes.scala 110:25]
  assign imm_switch_216_io_in0 = w_internal_480; // @[Benes.scala 110:25]
  assign imm_switch_217_io_in0 = w_internal_482; // @[Benes.scala 110:25]
  assign imm_switch_218_io_in0 = w_internal_484; // @[Benes.scala 110:25]
  assign imm_switch_219_io_in0 = w_internal_486; // @[Benes.scala 110:25]
  assign imm_switch_220_io_in0 = w_internal_488; // @[Benes.scala 110:25]
  assign imm_switch_221_io_in0 = w_internal_490; // @[Benes.scala 110:25]
  assign imm_switch_222_io_in0 = w_internal_492; // @[Benes.scala 110:25]
  assign imm_switch_223_io_in0 = w_internal_494; // @[Benes.scala 110:25]
  assign imm_switch_224_io_in0 = w_internal_496; // @[Benes.scala 110:25]
  assign imm_switch_225_io_in0 = w_internal_500; // @[Benes.scala 110:25]
  assign imm_switch_226_io_in0 = w_internal_502; // @[Benes.scala 110:25]
  assign imm_switch_227_io_in0 = w_internal_504; // @[Benes.scala 110:25]
  assign imm_switch_228_io_in0 = w_internal_506; // @[Benes.scala 110:25]
  assign imm_switch_229_io_in0 = w_internal_508; // @[Benes.scala 110:25]
  assign imm_switch_230_io_in0 = w_internal_510; // @[Benes.scala 110:25]
  assign imm_switch_231_io_in0 = w_internal_512; // @[Benes.scala 110:25]
  assign imm_switch_232_io_in0 = w_internal_514; // @[Benes.scala 110:25]
  assign imm_switch_233_io_in0 = w_internal_516; // @[Benes.scala 110:25]
  assign imm_switch_234_io_in0 = w_internal_520; // @[Benes.scala 110:25]
  assign imm_switch_235_io_in0 = w_internal_522; // @[Benes.scala 110:25]
  assign imm_switch_236_io_in0 = w_internal_524; // @[Benes.scala 110:25]
  assign imm_switch_237_io_in0 = w_internal_526; // @[Benes.scala 110:25]
  assign imm_switch_238_io_in0 = w_internal_528; // @[Benes.scala 110:25]
  assign imm_switch_239_io_in0 = w_internal_530; // @[Benes.scala 110:25]
  assign imm_switch_240_io_in0 = w_internal_532; // @[Benes.scala 110:25]
  assign imm_switch_241_io_in0 = w_internal_534; // @[Benes.scala 110:25]
  assign imm_switch_242_io_in0 = w_internal_536; // @[Benes.scala 110:25]
  assign imm_switch_243_io_in0 = w_internal_540; // @[Benes.scala 110:25]
  assign imm_switch_244_io_in0 = w_internal_542; // @[Benes.scala 110:25]
  assign imm_switch_245_io_in0 = w_internal_544; // @[Benes.scala 110:25]
  assign imm_switch_246_io_in0 = w_internal_546; // @[Benes.scala 110:25]
  assign imm_switch_247_io_in0 = w_internal_548; // @[Benes.scala 110:25]
  assign imm_switch_248_io_in0 = w_internal_550; // @[Benes.scala 110:25]
  assign imm_switch_249_io_in0 = w_internal_552; // @[Benes.scala 110:25]
  assign imm_switch_250_io_in0 = w_internal_554; // @[Benes.scala 110:25]
  assign imm_switch_251_io_in0 = w_internal_556; // @[Benes.scala 110:25]
  assign imm_switch_252_io_in0 = w_internal_560; // @[Benes.scala 110:25]
  assign imm_switch_253_io_in0 = w_internal_562; // @[Benes.scala 110:25]
  assign imm_switch_254_io_in0 = w_internal_564; // @[Benes.scala 110:25]
  assign imm_switch_255_io_in0 = w_internal_566; // @[Benes.scala 110:25]
  assign imm_switch_256_io_in0 = w_internal_568; // @[Benes.scala 110:25]
  assign imm_switch_257_io_in0 = w_internal_570; // @[Benes.scala 110:25]
  assign imm_switch_258_io_in0 = w_internal_572; // @[Benes.scala 110:25]
  assign imm_switch_259_io_in0 = w_internal_574; // @[Benes.scala 110:25]
  assign imm_switch_260_io_in0 = w_internal_576; // @[Benes.scala 110:25]
  assign imm_switch_261_io_in0 = w_internal_580; // @[Benes.scala 110:25]
  assign imm_switch_262_io_in0 = w_internal_582; // @[Benes.scala 110:25]
  assign imm_switch_263_io_in0 = w_internal_584; // @[Benes.scala 110:25]
  assign imm_switch_264_io_in0 = w_internal_586; // @[Benes.scala 110:25]
  assign imm_switch_265_io_in0 = w_internal_588; // @[Benes.scala 110:25]
  assign imm_switch_266_io_in0 = w_internal_590; // @[Benes.scala 110:25]
  assign imm_switch_267_io_in0 = w_internal_592; // @[Benes.scala 110:25]
  assign imm_switch_268_io_in0 = w_internal_594; // @[Benes.scala 110:25]
  assign imm_switch_269_io_in0 = w_internal_596; // @[Benes.scala 110:25]
  assign imm_switch_270_io_in0 = w_internal_600; // @[Benes.scala 110:25]
  assign imm_switch_271_io_in0 = w_internal_602; // @[Benes.scala 110:25]
  assign imm_switch_272_io_in0 = w_internal_604; // @[Benes.scala 110:25]
  assign imm_switch_273_io_in0 = w_internal_606; // @[Benes.scala 110:25]
  assign imm_switch_274_io_in0 = w_internal_608; // @[Benes.scala 110:25]
  assign imm_switch_275_io_in0 = w_internal_610; // @[Benes.scala 110:25]
  assign imm_switch_276_io_in0 = w_internal_612; // @[Benes.scala 110:25]
  assign imm_switch_277_io_in0 = w_internal_614; // @[Benes.scala 110:25]
  assign imm_switch_278_io_in0 = w_internal_616; // @[Benes.scala 110:25]
  assign imm_switch_279_io_in0 = w_internal_620; // @[Benes.scala 110:25]
  assign imm_switch_280_io_in0 = w_internal_622; // @[Benes.scala 110:25]
  assign imm_switch_281_io_in0 = w_internal_624; // @[Benes.scala 110:25]
  assign imm_switch_282_io_in0 = w_internal_626; // @[Benes.scala 110:25]
  assign imm_switch_283_io_in0 = w_internal_628; // @[Benes.scala 110:25]
  assign imm_switch_284_io_in0 = w_internal_630; // @[Benes.scala 110:25]
  assign imm_switch_285_io_in0 = w_internal_632; // @[Benes.scala 110:25]
  assign imm_switch_286_io_in0 = w_internal_634; // @[Benes.scala 110:25]
  assign imm_switch_287_io_in0 = w_internal_636; // @[Benes.scala 110:25]
  always @(posedge clock) begin
    if (reset) begin // @[Benes.scala 77:32]
      r_data_bus_ff_0 <= 16'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_data_bus_ff_0 <= 16'h0;
    end else begin
      r_data_bus_ff_0 <= 16'h1;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_data_bus_ff_1 <= 16'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_data_bus_ff_1 <= 16'h0;
    end else begin
      r_data_bus_ff_1 <= 16'h2;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_data_bus_ff_2 <= 16'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_data_bus_ff_2 <= 16'h0;
    end else begin
      r_data_bus_ff_2 <= 16'h3;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_data_bus_ff_3 <= 16'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_data_bus_ff_3 <= 16'h0;
    end else begin
      r_data_bus_ff_3 <= 16'h4;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_data_bus_ff_4 <= 16'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_data_bus_ff_4 <= 16'h0;
    end else begin
      r_data_bus_ff_4 <= 16'h5;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_data_bus_ff_5 <= 16'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_data_bus_ff_5 <= 16'h0;
    end else begin
      r_data_bus_ff_5 <= 16'h6;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_data_bus_ff_6 <= 16'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_data_bus_ff_6 <= 16'h0;
    end else begin
      r_data_bus_ff_6 <= 16'h7;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_data_bus_ff_7 <= 16'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_data_bus_ff_7 <= 16'h0;
    end else begin
      r_data_bus_ff_7 <= 16'h8;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_data_bus_ff_8 <= 16'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_data_bus_ff_8 <= 16'h0;
    end else begin
      r_data_bus_ff_8 <= 16'h9;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_data_bus_ff_9 <= 16'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_data_bus_ff_9 <= 16'h0;
    end else begin
      r_data_bus_ff_9 <= 16'ha;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_data_bus_ff_10 <= 16'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_data_bus_ff_10 <= 16'h0;
    end else begin
      r_data_bus_ff_10 <= 16'h1;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_data_bus_ff_11 <= 16'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_data_bus_ff_11 <= 16'h0;
    end else begin
      r_data_bus_ff_11 <= 16'h2;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_data_bus_ff_12 <= 16'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_data_bus_ff_12 <= 16'h0;
    end else begin
      r_data_bus_ff_12 <= 16'h3;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_data_bus_ff_13 <= 16'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_data_bus_ff_13 <= 16'h0;
    end else begin
      r_data_bus_ff_13 <= 16'h4;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_data_bus_ff_14 <= 16'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_data_bus_ff_14 <= 16'h0;
    end else begin
      r_data_bus_ff_14 <= 16'h5;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_data_bus_ff_15 <= 16'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_data_bus_ff_15 <= 16'h0;
    end else begin
      r_data_bus_ff_15 <= 16'h6;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_data_bus_ff_16 <= 16'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_data_bus_ff_16 <= 16'h0;
    end else begin
      r_data_bus_ff_16 <= 16'h7;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_data_bus_ff_17 <= 16'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_data_bus_ff_17 <= 16'h0;
    end else begin
      r_data_bus_ff_17 <= 16'h8;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_data_bus_ff_18 <= 16'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_data_bus_ff_18 <= 16'h0;
    end else begin
      r_data_bus_ff_18 <= 16'h9;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_data_bus_ff_19 <= 16'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_data_bus_ff_19 <= 16'h0;
    end else begin
      r_data_bus_ff_19 <= 16'ha;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_data_bus_ff_20 <= 16'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_data_bus_ff_20 <= 16'h0;
    end else begin
      r_data_bus_ff_20 <= 16'h1;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_data_bus_ff_21 <= 16'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_data_bus_ff_21 <= 16'h0;
    end else begin
      r_data_bus_ff_21 <= 16'h2;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_data_bus_ff_22 <= 16'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_data_bus_ff_22 <= 16'h0;
    end else begin
      r_data_bus_ff_22 <= 16'h3;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_data_bus_ff_23 <= 16'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_data_bus_ff_23 <= 16'h0;
    end else begin
      r_data_bus_ff_23 <= 16'h4;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_data_bus_ff_24 <= 16'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_data_bus_ff_24 <= 16'h0;
    end else begin
      r_data_bus_ff_24 <= 16'h5;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_data_bus_ff_25 <= 16'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_data_bus_ff_25 <= 16'h0;
    end else begin
      r_data_bus_ff_25 <= 16'h6;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_data_bus_ff_26 <= 16'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_data_bus_ff_26 <= 16'h0;
    end else begin
      r_data_bus_ff_26 <= 16'h7;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_data_bus_ff_27 <= 16'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_data_bus_ff_27 <= 16'h0;
    end else begin
      r_data_bus_ff_27 <= 16'h8;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_data_bus_ff_28 <= 16'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_data_bus_ff_28 <= 16'h0;
    end else begin
      r_data_bus_ff_28 <= 16'h9;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_data_bus_ff_29 <= 16'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_data_bus_ff_29 <= 16'h0;
    end else begin
      r_data_bus_ff_29 <= 16'ha;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_data_bus_ff_30 <= 16'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_data_bus_ff_30 <= 16'h0;
    end else begin
      r_data_bus_ff_30 <= 16'h1f;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_data_bus_ff_31 <= 16'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_data_bus_ff_31 <= 16'h0;
    end else begin
      r_data_bus_ff_31 <= 16'h20;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_data_bus_ff_0 = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  r_data_bus_ff_1 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  r_data_bus_ff_2 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  r_data_bus_ff_3 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  r_data_bus_ff_4 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  r_data_bus_ff_5 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  r_data_bus_ff_6 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  r_data_bus_ff_7 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  r_data_bus_ff_8 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  r_data_bus_ff_9 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  r_data_bus_ff_10 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  r_data_bus_ff_11 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  r_data_bus_ff_12 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  r_data_bus_ff_13 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  r_data_bus_ff_14 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  r_data_bus_ff_15 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  r_data_bus_ff_16 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  r_data_bus_ff_17 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  r_data_bus_ff_18 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  r_data_bus_ff_19 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  r_data_bus_ff_20 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  r_data_bus_ff_21 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  r_data_bus_ff_22 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  r_data_bus_ff_23 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  r_data_bus_ff_24 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  r_data_bus_ff_25 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  r_data_bus_ff_26 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  r_data_bus_ff_27 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  r_data_bus_ff_28 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  r_data_bus_ff_29 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  r_data_bus_ff_30 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  r_data_bus_ff_31 = _RAND_31[15:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module buffer_multiplication(
  input  [15:0] io_buffer2_0,
  input  [15:0] io_buffer2_1,
  input  [15:0] io_buffer2_2,
  input  [15:0] io_buffer2_3,
  input  [15:0] io_buffer2_4,
  input  [15:0] io_buffer2_5,
  input  [15:0] io_buffer2_6,
  input  [15:0] io_buffer2_7,
  input  [15:0] io_buffer2_8,
  input  [15:0] io_buffer2_9,
  input  [15:0] io_buffer2_10,
  input  [15:0] io_buffer2_11,
  input  [15:0] io_buffer2_12,
  input  [15:0] io_buffer2_13,
  input  [15:0] io_buffer2_14,
  input  [15:0] io_buffer2_15,
  input  [15:0] io_buffer2_16,
  input  [15:0] io_buffer2_17,
  input  [15:0] io_buffer2_18,
  input  [15:0] io_buffer2_19,
  input  [15:0] io_buffer2_20,
  input  [15:0] io_buffer2_21,
  input  [15:0] io_buffer2_22,
  input  [15:0] io_buffer2_23,
  input  [15:0] io_buffer2_24,
  input  [15:0] io_buffer2_25,
  input  [15:0] io_buffer2_26,
  input  [15:0] io_buffer2_27,
  input  [15:0] io_buffer2_28,
  input  [15:0] io_buffer2_29,
  input  [15:0] io_buffer2_30,
  input  [15:0] io_buffer2_31,
  output [15:0] io_out_0,
  output [15:0] io_out_1,
  output [15:0] io_out_2,
  output [15:0] io_out_3,
  output [15:0] io_out_4,
  output [15:0] io_out_5,
  output [15:0] io_out_6,
  output [15:0] io_out_7,
  output [15:0] io_out_8,
  output [15:0] io_out_9,
  output [15:0] io_out_10,
  output [15:0] io_out_11,
  output [15:0] io_out_12,
  output [15:0] io_out_13,
  output [15:0] io_out_14,
  output [15:0] io_out_15,
  output [15:0] io_out_16,
  output [15:0] io_out_17,
  output [15:0] io_out_18,
  output [15:0] io_out_19,
  output [15:0] io_out_20,
  output [15:0] io_out_21,
  output [15:0] io_out_22,
  output [15:0] io_out_23,
  output [15:0] io_out_24,
  output [15:0] io_out_25,
  output [15:0] io_out_26,
  output [15:0] io_out_27,
  output [15:0] io_out_28,
  output [15:0] io_out_29,
  output [15:0] io_out_30,
  output [15:0] io_out_31
);
  wire [31:0] elementMul = 16'h1 * io_buffer2_0; // @[buffer_multiplication.scala 17:42]
  wire [31:0] result_elementMul = 16'h2 * io_buffer2_1; // @[buffer_multiplication.scala 17:42]
  wire [31:0] result_result_elementMul = 16'h3 * io_buffer2_2; // @[buffer_multiplication.scala 17:42]
  wire [31:0] result_result_result_elementMul = 16'h4 * io_buffer2_3; // @[buffer_multiplication.scala 17:42]
  wire [31:0] result_result_result_result_elementMul = 16'h5 * io_buffer2_4; // @[buffer_multiplication.scala 17:42]
  wire [31:0] result_result_result_result_result_elementMul = 16'h6 * io_buffer2_5; // @[buffer_multiplication.scala 17:42]
  wire [31:0] result_result_result_result_result_result_elementMul = 16'h7 * io_buffer2_6; // @[buffer_multiplication.scala 17:42]
  wire [31:0] result_result_result_result_result_result_result_elementMul = 16'h8 * io_buffer2_7; // @[buffer_multiplication.scala 17:42]
  wire [31:0] result_result_result_result_result_result_result_result_elementMul = 16'h9 * io_buffer2_8; // @[buffer_multiplication.scala 17:42]
  wire [31:0] result_result_result_result_result_result_result_result_result_elementMul = 16'ha * io_buffer2_9; // @[buffer_multiplication.scala 17:42]
  wire [31:0] result_result_result_result_result_result_result_result_result_result_elementMul = 16'h1 * io_buffer2_10; // @[buffer_multiplication.scala 17:42]
  wire [31:0] result_result_result_result_result_result_result_result_result_result_result_elementMul = 16'h2 *
    io_buffer2_11; // @[buffer_multiplication.scala 17:42]
  wire [31:0] result_result_result_result_result_result_result_result_result_result_result_result_elementMul = 16'h3 *
    io_buffer2_12; // @[buffer_multiplication.scala 17:42]
  wire [31:0] result_result_result_result_result_result_result_result_result_result_result_result_result_elementMul = 16'h4
     * io_buffer2_13; // @[buffer_multiplication.scala 17:42]
  wire [31:0]
    result_result_result_result_result_result_result_result_result_result_result_result_result_result_elementMul = 16'h5
     * io_buffer2_14; // @[buffer_multiplication.scala 17:42]
  wire [31:0]
    result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_elementMul
     = 16'h6 * io_buffer2_15; // @[buffer_multiplication.scala 17:42]
  wire [31:0]
    result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_elementMul
     = 16'h7 * io_buffer2_16; // @[buffer_multiplication.scala 17:42]
  wire [31:0]
    result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_elementMul
     = 16'h8 * io_buffer2_17; // @[buffer_multiplication.scala 17:42]
  wire [31:0]
    result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_elementMul
     = 16'h9 * io_buffer2_18; // @[buffer_multiplication.scala 17:42]
  wire [31:0]
    result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_elementMul
     = 16'ha * io_buffer2_19; // @[buffer_multiplication.scala 17:42]
  wire [31:0]
    result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_elementMul
     = 16'h1 * io_buffer2_20; // @[buffer_multiplication.scala 17:42]
  wire [31:0]
    result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_elementMul
     = 16'h2 * io_buffer2_21; // @[buffer_multiplication.scala 17:42]
  wire [31:0]
    result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_elementMul
     = 16'h3 * io_buffer2_22; // @[buffer_multiplication.scala 17:42]
  wire [31:0]
    result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_elementMul
     = 16'h4 * io_buffer2_23; // @[buffer_multiplication.scala 17:42]
  wire [31:0]
    result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_elementMul
     = 16'h5 * io_buffer2_24; // @[buffer_multiplication.scala 17:42]
  wire [31:0]
    result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_elementMul
     = 16'h6 * io_buffer2_25; // @[buffer_multiplication.scala 17:42]
  wire [31:0]
    result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_elementMul
     = 16'h7 * io_buffer2_26; // @[buffer_multiplication.scala 17:42]
  wire [31:0]
    result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_elementMul
     = 16'h8 * io_buffer2_27; // @[buffer_multiplication.scala 17:42]
  wire [31:0]
    result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_elementMul
     = 16'h9 * io_buffer2_28; // @[buffer_multiplication.scala 17:42]
  wire [31:0]
    result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_elementMul
     = 16'ha * io_buffer2_29; // @[buffer_multiplication.scala 17:42]
  wire [31:0]
    result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_elementMul
     = 16'h1f * io_buffer2_30; // @[buffer_multiplication.scala 17:42]
  wire [31:0]
    result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_elementMul
     = 16'h20 * io_buffer2_31; // @[buffer_multiplication.scala 17:42]
  assign io_out_0 = elementMul[15:0]; // @[buffer_multiplication.scala 15:20 19:27]
  assign io_out_1 = result_elementMul[15:0]; // @[buffer_multiplication.scala 15:20 19:27]
  assign io_out_2 = result_result_elementMul[15:0]; // @[buffer_multiplication.scala 15:20 19:27]
  assign io_out_3 = result_result_result_elementMul[15:0]; // @[buffer_multiplication.scala 15:20 19:27]
  assign io_out_4 = result_result_result_result_elementMul[15:0]; // @[buffer_multiplication.scala 15:20 19:27]
  assign io_out_5 = result_result_result_result_result_elementMul[15:0]; // @[buffer_multiplication.scala 15:20 19:27]
  assign io_out_6 = result_result_result_result_result_result_elementMul[15:0]; // @[buffer_multiplication.scala 15:20 19:27]
  assign io_out_7 = result_result_result_result_result_result_result_elementMul[15:0]; // @[buffer_multiplication.scala 15:20 19:27]
  assign io_out_8 = result_result_result_result_result_result_result_result_elementMul[15:0]; // @[buffer_multiplication.scala 15:20 19:27]
  assign io_out_9 = result_result_result_result_result_result_result_result_result_elementMul[15:0]; // @[buffer_multiplication.scala 15:20 19:27]
  assign io_out_10 = result_result_result_result_result_result_result_result_result_result_elementMul[15:0]; // @[buffer_multiplication.scala 15:20 19:27]
  assign io_out_11 = result_result_result_result_result_result_result_result_result_result_result_elementMul[15:0]; // @[buffer_multiplication.scala 15:20 19:27]
  assign io_out_12 = result_result_result_result_result_result_result_result_result_result_result_result_elementMul[15:0
    ]; // @[buffer_multiplication.scala 15:20 19:27]
  assign io_out_13 =
    result_result_result_result_result_result_result_result_result_result_result_result_result_elementMul[15:0]; // @[buffer_multiplication.scala 15:20 19:27]
  assign io_out_14 =
    result_result_result_result_result_result_result_result_result_result_result_result_result_result_elementMul[15:0]; // @[buffer_multiplication.scala 15:20 19:27]
  assign io_out_15 =
    result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_elementMul[
    15:0]; // @[buffer_multiplication.scala 15:20 19:27]
  assign io_out_16 =
    result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_elementMul
    [15:0]; // @[buffer_multiplication.scala 15:20 19:27]
  assign io_out_17 =
    result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_elementMul
    [15:0]; // @[buffer_multiplication.scala 15:20 19:27]
  assign io_out_18 =
    result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_elementMul
    [15:0]; // @[buffer_multiplication.scala 15:20 19:27]
  assign io_out_19 =
    result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_elementMul
    [15:0]; // @[buffer_multiplication.scala 15:20 19:27]
  assign io_out_20 =
    result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_elementMul
    [15:0]; // @[buffer_multiplication.scala 15:20 19:27]
  assign io_out_21 =
    result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_elementMul
    [15:0]; // @[buffer_multiplication.scala 15:20 19:27]
  assign io_out_22 =
    result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_elementMul
    [15:0]; // @[buffer_multiplication.scala 15:20 19:27]
  assign io_out_23 =
    result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_elementMul
    [15:0]; // @[buffer_multiplication.scala 15:20 19:27]
  assign io_out_24 =
    result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_elementMul
    [15:0]; // @[buffer_multiplication.scala 15:20 19:27]
  assign io_out_25 =
    result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_elementMul
    [15:0]; // @[buffer_multiplication.scala 15:20 19:27]
  assign io_out_26 =
    result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_elementMul
    [15:0]; // @[buffer_multiplication.scala 15:20 19:27]
  assign io_out_27 =
    result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_elementMul
    [15:0]; // @[buffer_multiplication.scala 15:20 19:27]
  assign io_out_28 =
    result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_elementMul
    [15:0]; // @[buffer_multiplication.scala 15:20 19:27]
  assign io_out_29 =
    result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_elementMul
    [15:0]; // @[buffer_multiplication.scala 15:20 19:27]
  assign io_out_30 =
    result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_elementMul
    [15:0]; // @[buffer_multiplication.scala 15:20 19:27]
  assign io_out_31 =
    result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_result_elementMul
    [15:0]; // @[buffer_multiplication.scala 15:20 19:27]
endmodule
module ReductionMux(
  input  [31:0] io_i_data_0,
  input  [31:0] io_i_data_1,
  output [31:0] io_o_data_0,
  output [31:0] io_o_data_1
);
  assign io_o_data_0 = io_i_data_0; // @[ReductionMux.scala 31:39 33:18 35:18]
  assign io_o_data_1 = io_i_data_1; // @[ReductionMux.scala 37:22]
endmodule
module SimpleAdder(
  input  [31:0] io_A,
  input  [31:0] io_B,
  output [31:0] io_O
);
  assign io_O = io_A + io_B; // @[SimpleAdder.scala 14:18]
endmodule
module EdgeAdderSwitch(
  input         clock,
  input         reset,
  input         io_i_valid,
  input  [63:0] io_i_data_bus_0,
  input  [63:0] io_i_data_bus_1,
  input  [2:0]  io_i_add_en,
  input  [4:0]  io_i_cmd,
  output [63:0] io_o_vn,
  output [1:0]  io_o_vn_valid,
  output [31:0] io_o_adder
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] reductionMux_io_i_data_0; // @[EdgeAdderSwitch.scala 19:28]
  wire [31:0] reductionMux_io_i_data_1; // @[EdgeAdderSwitch.scala 19:28]
  wire [31:0] reductionMux_io_o_data_0; // @[EdgeAdderSwitch.scala 19:28]
  wire [31:0] reductionMux_io_o_data_1; // @[EdgeAdderSwitch.scala 19:28]
  wire [31:0] adder32_io_A; // @[EdgeAdderSwitch.scala 23:23]
  wire [31:0] adder32_io_B; // @[EdgeAdderSwitch.scala 23:23]
  wire [31:0] adder32_io_O; // @[EdgeAdderSwitch.scala 23:23]
  reg  r_valid; // @[EdgeAdderSwitch.scala 27:24]
  reg [31:0] r_adder; // @[EdgeAdderSwitch.scala 28:24]
  reg [63:0] r_vn; // @[EdgeAdderSwitch.scala 29:21]
  reg [1:0] r_vn_valid; // @[EdgeAdderSwitch.scala 30:27]
  reg [2:0] r_add_en; // @[EdgeAdderSwitch.scala 31:25]
  wire [95:0] _r_vn_T = {io_i_data_bus_0,32'h0}; // @[Cat.scala 33:92]
  wire [95:0] _r_vn_T_1 = {32'h0,io_i_data_bus_1}; // @[Cat.scala 33:92]
  wire [63:0] _r_vn_T_2 = {reductionMux_io_o_data_0,reductionMux_io_o_data_1}; // @[Cat.scala 33:92]
  wire [1:0] _GEN_0 = 5'h0 == io_i_cmd ? 2'h0 : r_vn_valid; // @[EdgeAdderSwitch.scala 38:23 54:20 30:27]
  wire [63:0] _GEN_1 = 5'h5 == io_i_cmd ? _r_vn_T_2 : r_vn; // @[EdgeAdderSwitch.scala 38:23 50:14 29:21]
  wire [1:0] _GEN_2 = 5'h5 == io_i_cmd ? 2'h3 : _GEN_0; // @[EdgeAdderSwitch.scala 38:23 51:20]
  wire [31:0] _GEN_3 = 5'h4 == io_i_cmd ? reductionMux_io_o_data_0 : r_adder; // @[EdgeAdderSwitch.scala 38:23 45:17 28:24]
  wire [95:0] _GEN_4 = 5'h4 == io_i_cmd ? _r_vn_T_1 : {{32'd0}, _GEN_1}; // @[EdgeAdderSwitch.scala 38:23 46:14]
  wire [1:0] _GEN_5 = 5'h4 == io_i_cmd ? 2'h2 : _GEN_2; // @[EdgeAdderSwitch.scala 38:23 47:20]
  wire [95:0] _GEN_7 = 5'h3 == io_i_cmd ? _r_vn_T : _GEN_4; // @[EdgeAdderSwitch.scala 38:23 41:14]
  wire [95:0] _GEN_10 = r_valid ? _GEN_7 : {{32'd0}, r_vn}; // @[EdgeAdderSwitch.scala 29:21 37:25]
  wire [95:0] _GEN_13 = reset ? 96'h0 : _GEN_10; // @[EdgeAdderSwitch.scala 33:14 35:10]
  wire [31:0] _GEN_15 = r_add_en == 3'h0 ? r_adder : adder32_io_O; // @[EdgeAdderSwitch.scala 64:22 65:18 67:18]
  wire [95:0] _GEN_19 = reset ? 96'h0 : _GEN_13; // @[EdgeAdderSwitch.scala 29:{21,21}]
  ReductionMux reductionMux ( // @[EdgeAdderSwitch.scala 19:28]
    .io_i_data_0(reductionMux_io_i_data_0),
    .io_i_data_1(reductionMux_io_i_data_1),
    .io_o_data_0(reductionMux_io_o_data_0),
    .io_o_data_1(reductionMux_io_o_data_1)
  );
  SimpleAdder adder32 ( // @[EdgeAdderSwitch.scala 23:23]
    .io_A(adder32_io_A),
    .io_B(adder32_io_B),
    .io_O(adder32_io_O)
  );
  assign io_o_vn = reset ? 64'h0 : r_vn; // @[EdgeAdderSwitch.scala 59:14 61:13 69:13]
  assign io_o_vn_valid = reset ? 2'h0 : r_vn_valid; // @[EdgeAdderSwitch.scala 59:14 62:19 70:19]
  assign io_o_adder = reset ? 32'h0 : _GEN_15; // @[EdgeAdderSwitch.scala 59:14 60:16]
  assign reductionMux_io_i_data_0 = io_i_data_bus_0[31:0]; // @[EdgeAdderSwitch.scala 20:26]
  assign reductionMux_io_i_data_1 = io_i_data_bus_1[31:0]; // @[EdgeAdderSwitch.scala 20:26]
  assign adder32_io_A = reductionMux_io_o_data_1; // @[EdgeAdderSwitch.scala 24:16]
  assign adder32_io_B = reductionMux_io_o_data_0; // @[EdgeAdderSwitch.scala 25:16]
  always @(posedge clock) begin
    if (reset) begin // @[EdgeAdderSwitch.scala 27:24]
      r_valid <= 1'h0; // @[EdgeAdderSwitch.scala 27:24]
    end else begin
      r_valid <= io_i_valid; // @[EdgeAdderSwitch.scala 27:24]
    end
    if (reset) begin // @[EdgeAdderSwitch.scala 28:24]
      r_adder <= 32'h0; // @[EdgeAdderSwitch.scala 28:24]
    end else if (reset) begin // @[EdgeAdderSwitch.scala 33:14]
      r_adder <= 32'h0; // @[EdgeAdderSwitch.scala 34:13]
    end else if (r_valid) begin // @[EdgeAdderSwitch.scala 37:25]
      if (5'h3 == io_i_cmd) begin // @[EdgeAdderSwitch.scala 38:23]
        r_adder <= reductionMux_io_o_data_1; // @[EdgeAdderSwitch.scala 40:17]
      end else begin
        r_adder <= _GEN_3;
      end
    end
    r_vn <= _GEN_19[63:0]; // @[EdgeAdderSwitch.scala 29:{21,21}]
    if (reset) begin // @[EdgeAdderSwitch.scala 30:27]
      r_vn_valid <= 2'h0; // @[EdgeAdderSwitch.scala 30:27]
    end else if (reset) begin // @[EdgeAdderSwitch.scala 33:14]
      r_vn_valid <= 2'h0; // @[EdgeAdderSwitch.scala 36:16]
    end else if (r_valid) begin // @[EdgeAdderSwitch.scala 37:25]
      if (5'h3 == io_i_cmd) begin // @[EdgeAdderSwitch.scala 38:23]
        r_vn_valid <= 2'h1; // @[EdgeAdderSwitch.scala 42:20]
      end else begin
        r_vn_valid <= _GEN_5;
      end
    end
    if (reset) begin // @[EdgeAdderSwitch.scala 31:25]
      r_add_en <= 3'h0; // @[EdgeAdderSwitch.scala 31:25]
    end else begin
      r_add_en <= io_i_add_en; // @[EdgeAdderSwitch.scala 31:25]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  r_adder = _RAND_1[31:0];
  _RAND_2 = {2{`RANDOM}};
  r_vn = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  r_vn_valid = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  r_add_en = _RAND_4[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AdderSwitch(
  input         clock,
  input         reset,
  input         io_i_valid,
  input  [31:0] io_i_data_bus_0,
  input  [31:0] io_i_data_bus_1,
  input  [2:0]  io_i_add_en,
  input  [2:0]  io_i_cmd,
  output [1:0]  io_o_vn_valid,
  output [63:0] io_o_vn,
  output [31:0] io_o_adder_0,
  output [31:0] io_o_adder_1
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] reductionMux_io_i_data_0; // @[AdderSwitch.scala 21:28]
  wire [31:0] reductionMux_io_i_data_1; // @[AdderSwitch.scala 21:28]
  wire [31:0] reductionMux_io_o_data_0; // @[AdderSwitch.scala 21:28]
  wire [31:0] reductionMux_io_o_data_1; // @[AdderSwitch.scala 21:28]
  wire [31:0] adder32_io_A; // @[AdderSwitch.scala 25:23]
  wire [31:0] adder32_io_B; // @[AdderSwitch.scala 25:23]
  wire [31:0] adder32_io_O; // @[AdderSwitch.scala 25:23]
  reg [63:0] r_adder; // @[AdderSwitch.scala 29:24]
  reg [63:0] r_vn; // @[AdderSwitch.scala 30:21]
  reg [1:0] r_vn_valid; // @[AdderSwitch.scala 31:27]
  reg [2:0] r_add_en; // @[AdderSwitch.scala 32:25]
  wire [63:0] _r_adder_T = {reductionMux_io_o_data_0,reductionMux_io_o_data_1}; // @[Cat.scala 33:92]
  wire [62:0] _r_adder_T_1 = {31'h0,reductionMux_io_o_data_1}; // @[Cat.scala 33:92]
  wire [62:0] _r_adder_T_2 = {reductionMux_io_o_data_0,31'h0}; // @[Cat.scala 33:92]
  wire [1:0] _GEN_0 = 3'h0 == io_i_cmd ? 2'h0 : r_vn_valid; // @[AdderSwitch.scala 39:23 59:20 31:27]
  wire [63:0] _GEN_1 = 3'h5 == io_i_cmd ? _r_adder_T : r_vn; // @[AdderSwitch.scala 39:23 55:14 30:21]
  wire [1:0] _GEN_2 = 3'h5 == io_i_cmd ? 2'h3 : _GEN_0; // @[AdderSwitch.scala 39:23 56:20]
  wire [63:0] _GEN_3 = 3'h4 == io_i_cmd ? {{1'd0}, _r_adder_T_2} : r_adder; // @[AdderSwitch.scala 39:23 50:17 29:24]
  wire [63:0] _GEN_4 = 3'h4 == io_i_cmd ? {{32'd0}, io_i_data_bus_1} : _GEN_1; // @[AdderSwitch.scala 39:23 51:14]
  wire [1:0] _GEN_5 = 3'h4 == io_i_cmd ? 2'h2 : _GEN_2; // @[AdderSwitch.scala 39:23 52:20]
  wire [63:0] _GEN_6 = 3'h3 == io_i_cmd ? {{1'd0}, _r_adder_T_1} : _GEN_3; // @[AdderSwitch.scala 39:23 45:17]
  wire [63:0] _GEN_7 = 3'h3 == io_i_cmd ? {{32'd0}, io_i_data_bus_0} : _GEN_4; // @[AdderSwitch.scala 39:23 46:14]
  wire [1:0] _GEN_8 = 3'h3 == io_i_cmd ? 2'h1 : _GEN_5; // @[AdderSwitch.scala 39:23 47:20]
  wire [31:0] _WIRE_2_0 = adder32_io_O; // @[AdderSwitch.scala 72:{28,28}]
  wire [31:0] _GEN_18 = r_add_en == 3'h0 ? r_adder[31:0] : _WIRE_2_0; // @[AdderSwitch.scala 69:22 70:18 72:18]
  wire [31:0] _GEN_19 = r_add_en == 3'h0 ? r_adder[63:32] : _WIRE_2_0; // @[AdderSwitch.scala 69:22 70:18 72:18]
  ReductionMux reductionMux ( // @[AdderSwitch.scala 21:28]
    .io_i_data_0(reductionMux_io_i_data_0),
    .io_i_data_1(reductionMux_io_i_data_1),
    .io_o_data_0(reductionMux_io_o_data_0),
    .io_o_data_1(reductionMux_io_o_data_1)
  );
  SimpleAdder adder32 ( // @[AdderSwitch.scala 25:23]
    .io_A(adder32_io_A),
    .io_B(adder32_io_B),
    .io_O(adder32_io_O)
  );
  assign io_o_vn_valid = reset ? 2'h0 : r_vn_valid; // @[AdderSwitch.scala 64:14 67:19 75:19]
  assign io_o_vn = reset ? 64'h0 : r_vn; // @[AdderSwitch.scala 64:14 66:13 74:13]
  assign io_o_adder_0 = reset ? 32'h0 : _GEN_18; // @[AdderSwitch.scala 64:14 65:16]
  assign io_o_adder_1 = reset ? 32'h0 : _GEN_19; // @[AdderSwitch.scala 64:14 65:16]
  assign reductionMux_io_i_data_0 = io_i_data_bus_0; // @[AdderSwitch.scala 22:26]
  assign reductionMux_io_i_data_1 = io_i_data_bus_1; // @[AdderSwitch.scala 22:26]
  assign adder32_io_A = reductionMux_io_o_data_1; // @[AdderSwitch.scala 26:16]
  assign adder32_io_B = reductionMux_io_o_data_0; // @[AdderSwitch.scala 27:16]
  always @(posedge clock) begin
    if (reset) begin // @[AdderSwitch.scala 29:24]
      r_adder <= 64'h0; // @[AdderSwitch.scala 29:24]
    end else if (reset) begin // @[AdderSwitch.scala 34:14]
      r_adder <= 64'h0; // @[AdderSwitch.scala 35:13]
    end else if (io_i_valid) begin // @[AdderSwitch.scala 38:28]
      if (3'h1 == io_i_cmd) begin // @[AdderSwitch.scala 39:23]
        r_adder <= _r_adder_T; // @[AdderSwitch.scala 41:17]
      end else begin
        r_adder <= _GEN_6;
      end
    end
    if (reset) begin // @[AdderSwitch.scala 30:21]
      r_vn <= 64'h0; // @[AdderSwitch.scala 30:21]
    end else if (reset) begin // @[AdderSwitch.scala 34:14]
      r_vn <= 64'h0; // @[AdderSwitch.scala 36:10]
    end else if (io_i_valid) begin // @[AdderSwitch.scala 38:28]
      if (!(3'h1 == io_i_cmd)) begin // @[AdderSwitch.scala 39:23]
        r_vn <= _GEN_7;
      end
    end
    if (reset) begin // @[AdderSwitch.scala 31:27]
      r_vn_valid <= 2'h0; // @[AdderSwitch.scala 31:27]
    end else if (reset) begin // @[AdderSwitch.scala 34:14]
      r_vn_valid <= 2'h0; // @[AdderSwitch.scala 37:16]
    end else if (io_i_valid) begin // @[AdderSwitch.scala 38:28]
      if (3'h1 == io_i_cmd) begin // @[AdderSwitch.scala 39:23]
        r_vn_valid <= 2'h0; // @[AdderSwitch.scala 42:20]
      end else begin
        r_vn_valid <= _GEN_8;
      end
    end
    if (reset) begin // @[AdderSwitch.scala 32:25]
      r_add_en <= 3'h0; // @[AdderSwitch.scala 32:25]
    end else begin
      r_add_en <= io_i_add_en; // @[AdderSwitch.scala 32:25]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  r_adder = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  r_vn = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  r_vn_valid = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  r_add_en = _RAND_3[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ReductionMux_3(
  input  [31:0] io_i_data_0,
  input  [31:0] io_i_data_1,
  input  [31:0] io_i_data_2,
  input  [31:0] io_i_data_3,
  input  [1:0]  io_i_sel,
  output [31:0] io_o_data_0,
  output [31:0] io_o_data_1
);
  wire  w_sel_in_left = io_i_sel[0]; // @[ReductionMux.scala 28:32]
  wire  w_sel_in_right = io_i_sel[1]; // @[ReductionMux.scala 29:33]
  assign io_o_data_0 = w_sel_in_left ? io_i_data_1 : io_i_data_0; // @[ReductionMux.scala 33:{18,18}]
  assign io_o_data_1 = w_sel_in_right ? io_i_data_3 : io_i_data_2; // @[ReductionMux.scala 37:{22,22}]
endmodule
module EdgeAdderSwitch_2(
  input         clock,
  input         reset,
  input         io_i_valid,
  input  [63:0] io_i_data_bus_0,
  input  [63:0] io_i_data_bus_1,
  input  [63:0] io_i_data_bus_2,
  input  [63:0] io_i_data_bus_3,
  input  [2:0]  io_i_add_en,
  input  [4:0]  io_i_cmd,
  input  [1:0]  io_i_sel,
  output [63:0] io_o_vn,
  output [1:0]  io_o_vn_valid,
  output [31:0] io_o_adder
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] reductionMux_io_i_data_0; // @[EdgeAdderSwitch.scala 19:28]
  wire [31:0] reductionMux_io_i_data_1; // @[EdgeAdderSwitch.scala 19:28]
  wire [31:0] reductionMux_io_i_data_2; // @[EdgeAdderSwitch.scala 19:28]
  wire [31:0] reductionMux_io_i_data_3; // @[EdgeAdderSwitch.scala 19:28]
  wire [1:0] reductionMux_io_i_sel; // @[EdgeAdderSwitch.scala 19:28]
  wire [31:0] reductionMux_io_o_data_0; // @[EdgeAdderSwitch.scala 19:28]
  wire [31:0] reductionMux_io_o_data_1; // @[EdgeAdderSwitch.scala 19:28]
  wire [31:0] adder32_io_A; // @[EdgeAdderSwitch.scala 23:23]
  wire [31:0] adder32_io_B; // @[EdgeAdderSwitch.scala 23:23]
  wire [31:0] adder32_io_O; // @[EdgeAdderSwitch.scala 23:23]
  reg  r_valid; // @[EdgeAdderSwitch.scala 27:24]
  reg [31:0] r_adder; // @[EdgeAdderSwitch.scala 28:24]
  reg [63:0] r_vn; // @[EdgeAdderSwitch.scala 29:21]
  reg [1:0] r_vn_valid; // @[EdgeAdderSwitch.scala 30:27]
  reg [2:0] r_add_en; // @[EdgeAdderSwitch.scala 31:25]
  wire [95:0] _r_vn_T = {io_i_data_bus_0,32'h0}; // @[Cat.scala 33:92]
  wire [95:0] _r_vn_T_1 = {32'h0,io_i_data_bus_3}; // @[Cat.scala 33:92]
  wire [63:0] _r_vn_T_2 = {reductionMux_io_o_data_0,reductionMux_io_o_data_1}; // @[Cat.scala 33:92]
  wire [1:0] _GEN_0 = 5'h0 == io_i_cmd ? 2'h0 : r_vn_valid; // @[EdgeAdderSwitch.scala 38:23 54:20 30:27]
  wire [63:0] _GEN_1 = 5'h5 == io_i_cmd ? _r_vn_T_2 : r_vn; // @[EdgeAdderSwitch.scala 38:23 50:14 29:21]
  wire [1:0] _GEN_2 = 5'h5 == io_i_cmd ? 2'h3 : _GEN_0; // @[EdgeAdderSwitch.scala 38:23 51:20]
  wire [31:0] _GEN_3 = 5'h4 == io_i_cmd ? reductionMux_io_o_data_0 : r_adder; // @[EdgeAdderSwitch.scala 38:23 45:17 28:24]
  wire [95:0] _GEN_4 = 5'h4 == io_i_cmd ? _r_vn_T_1 : {{32'd0}, _GEN_1}; // @[EdgeAdderSwitch.scala 38:23 46:14]
  wire [1:0] _GEN_5 = 5'h4 == io_i_cmd ? 2'h2 : _GEN_2; // @[EdgeAdderSwitch.scala 38:23 47:20]
  wire [95:0] _GEN_7 = 5'h3 == io_i_cmd ? _r_vn_T : _GEN_4; // @[EdgeAdderSwitch.scala 38:23 41:14]
  wire [95:0] _GEN_10 = r_valid ? _GEN_7 : {{32'd0}, r_vn}; // @[EdgeAdderSwitch.scala 29:21 37:25]
  wire [95:0] _GEN_13 = reset ? 96'h0 : _GEN_10; // @[EdgeAdderSwitch.scala 33:14 35:10]
  wire [31:0] _GEN_15 = r_add_en == 3'h0 ? r_adder : adder32_io_O; // @[EdgeAdderSwitch.scala 64:22 65:18 67:18]
  wire [95:0] _GEN_19 = reset ? 96'h0 : _GEN_13; // @[EdgeAdderSwitch.scala 29:{21,21}]
  ReductionMux_3 reductionMux ( // @[EdgeAdderSwitch.scala 19:28]
    .io_i_data_0(reductionMux_io_i_data_0),
    .io_i_data_1(reductionMux_io_i_data_1),
    .io_i_data_2(reductionMux_io_i_data_2),
    .io_i_data_3(reductionMux_io_i_data_3),
    .io_i_sel(reductionMux_io_i_sel),
    .io_o_data_0(reductionMux_io_o_data_0),
    .io_o_data_1(reductionMux_io_o_data_1)
  );
  SimpleAdder adder32 ( // @[EdgeAdderSwitch.scala 23:23]
    .io_A(adder32_io_A),
    .io_B(adder32_io_B),
    .io_O(adder32_io_O)
  );
  assign io_o_vn = reset ? 64'h0 : r_vn; // @[EdgeAdderSwitch.scala 59:14 61:13 69:13]
  assign io_o_vn_valid = reset ? 2'h0 : r_vn_valid; // @[EdgeAdderSwitch.scala 59:14 62:19 70:19]
  assign io_o_adder = reset ? 32'h0 : _GEN_15; // @[EdgeAdderSwitch.scala 59:14 60:16]
  assign reductionMux_io_i_data_0 = io_i_data_bus_0[31:0]; // @[EdgeAdderSwitch.scala 20:26]
  assign reductionMux_io_i_data_1 = io_i_data_bus_1[31:0]; // @[EdgeAdderSwitch.scala 20:26]
  assign reductionMux_io_i_data_2 = io_i_data_bus_2[31:0]; // @[EdgeAdderSwitch.scala 20:26]
  assign reductionMux_io_i_data_3 = io_i_data_bus_3[31:0]; // @[EdgeAdderSwitch.scala 20:26]
  assign reductionMux_io_i_sel = io_i_sel; // @[EdgeAdderSwitch.scala 21:25]
  assign adder32_io_A = reductionMux_io_o_data_1; // @[EdgeAdderSwitch.scala 24:16]
  assign adder32_io_B = reductionMux_io_o_data_0; // @[EdgeAdderSwitch.scala 25:16]
  always @(posedge clock) begin
    if (reset) begin // @[EdgeAdderSwitch.scala 27:24]
      r_valid <= 1'h0; // @[EdgeAdderSwitch.scala 27:24]
    end else begin
      r_valid <= io_i_valid; // @[EdgeAdderSwitch.scala 27:24]
    end
    if (reset) begin // @[EdgeAdderSwitch.scala 28:24]
      r_adder <= 32'h0; // @[EdgeAdderSwitch.scala 28:24]
    end else if (reset) begin // @[EdgeAdderSwitch.scala 33:14]
      r_adder <= 32'h0; // @[EdgeAdderSwitch.scala 34:13]
    end else if (r_valid) begin // @[EdgeAdderSwitch.scala 37:25]
      if (5'h3 == io_i_cmd) begin // @[EdgeAdderSwitch.scala 38:23]
        r_adder <= reductionMux_io_o_data_1; // @[EdgeAdderSwitch.scala 40:17]
      end else begin
        r_adder <= _GEN_3;
      end
    end
    r_vn <= _GEN_19[63:0]; // @[EdgeAdderSwitch.scala 29:{21,21}]
    if (reset) begin // @[EdgeAdderSwitch.scala 30:27]
      r_vn_valid <= 2'h0; // @[EdgeAdderSwitch.scala 30:27]
    end else if (reset) begin // @[EdgeAdderSwitch.scala 33:14]
      r_vn_valid <= 2'h0; // @[EdgeAdderSwitch.scala 36:16]
    end else if (r_valid) begin // @[EdgeAdderSwitch.scala 37:25]
      if (5'h3 == io_i_cmd) begin // @[EdgeAdderSwitch.scala 38:23]
        r_vn_valid <= 2'h1; // @[EdgeAdderSwitch.scala 42:20]
      end else begin
        r_vn_valid <= _GEN_5;
      end
    end
    if (reset) begin // @[EdgeAdderSwitch.scala 31:25]
      r_add_en <= 3'h0; // @[EdgeAdderSwitch.scala 31:25]
    end else begin
      r_add_en <= io_i_add_en; // @[EdgeAdderSwitch.scala 31:25]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  r_adder = _RAND_1[31:0];
  _RAND_2 = {2{`RANDOM}};
  r_vn = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  r_vn_valid = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  r_add_en = _RAND_4[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ReductionMux_7(
  input  [31:0] io_i_data_0,
  input  [31:0] io_i_data_1,
  input  [31:0] io_i_data_2,
  input  [31:0] io_i_data_3,
  input  [31:0] io_i_data_4,
  input  [31:0] io_i_data_5,
  input  [3:0]  io_i_sel,
  output [31:0] io_o_data_0,
  output [31:0] io_o_data_1
);
  wire [1:0] w_sel_in_left = io_i_sel[1:0]; // @[ReductionMux.scala 28:32]
  wire [1:0] w_sel_in_right = io_i_sel[3:2]; // @[ReductionMux.scala 29:33]
  wire [31:0] _GEN_1 = 2'h1 == w_sel_in_left ? io_i_data_1 : io_i_data_0; // @[ReductionMux.scala 33:{18,18}]
  wire [31:0] _GEN_2 = 2'h2 == w_sel_in_left ? io_i_data_2 : _GEN_1; // @[ReductionMux.scala 33:{18,18}]
  wire [31:0] _GEN_5 = 2'h1 == w_sel_in_right ? io_i_data_4 : io_i_data_3; // @[ReductionMux.scala 37:{22,22}]
  wire [31:0] _GEN_6 = 2'h2 == w_sel_in_right ? io_i_data_5 : _GEN_5; // @[ReductionMux.scala 37:{22,22}]
  assign io_o_data_0 = w_sel_in_left < 2'h2 ? _GEN_2 : 32'h0; // @[ReductionMux.scala 31:39 33:18 35:18]
  assign io_o_data_1 = w_sel_in_right < 2'h3 ? _GEN_6 : 32'h0; // @[ReductionMux.scala 37:22]
endmodule
module EdgeAdderSwitch_3(
  input         clock,
  input         reset,
  input         io_i_valid,
  input  [63:0] io_i_data_bus_0,
  input  [63:0] io_i_data_bus_1,
  input  [63:0] io_i_data_bus_2,
  input  [63:0] io_i_data_bus_3,
  input  [63:0] io_i_data_bus_4,
  input  [63:0] io_i_data_bus_5,
  input  [2:0]  io_i_add_en,
  input  [4:0]  io_i_cmd,
  input  [3:0]  io_i_sel,
  output [63:0] io_o_vn,
  output [1:0]  io_o_vn_valid,
  output [31:0] io_o_adder
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] reductionMux_io_i_data_0; // @[EdgeAdderSwitch.scala 19:28]
  wire [31:0] reductionMux_io_i_data_1; // @[EdgeAdderSwitch.scala 19:28]
  wire [31:0] reductionMux_io_i_data_2; // @[EdgeAdderSwitch.scala 19:28]
  wire [31:0] reductionMux_io_i_data_3; // @[EdgeAdderSwitch.scala 19:28]
  wire [31:0] reductionMux_io_i_data_4; // @[EdgeAdderSwitch.scala 19:28]
  wire [31:0] reductionMux_io_i_data_5; // @[EdgeAdderSwitch.scala 19:28]
  wire [3:0] reductionMux_io_i_sel; // @[EdgeAdderSwitch.scala 19:28]
  wire [31:0] reductionMux_io_o_data_0; // @[EdgeAdderSwitch.scala 19:28]
  wire [31:0] reductionMux_io_o_data_1; // @[EdgeAdderSwitch.scala 19:28]
  wire [31:0] adder32_io_A; // @[EdgeAdderSwitch.scala 23:23]
  wire [31:0] adder32_io_B; // @[EdgeAdderSwitch.scala 23:23]
  wire [31:0] adder32_io_O; // @[EdgeAdderSwitch.scala 23:23]
  reg  r_valid; // @[EdgeAdderSwitch.scala 27:24]
  reg [31:0] r_adder; // @[EdgeAdderSwitch.scala 28:24]
  reg [63:0] r_vn; // @[EdgeAdderSwitch.scala 29:21]
  reg [1:0] r_vn_valid; // @[EdgeAdderSwitch.scala 30:27]
  reg [2:0] r_add_en; // @[EdgeAdderSwitch.scala 31:25]
  wire [95:0] _r_vn_T = {io_i_data_bus_0,32'h0}; // @[Cat.scala 33:92]
  wire [95:0] _r_vn_T_1 = {32'h0,io_i_data_bus_5}; // @[Cat.scala 33:92]
  wire [63:0] _r_vn_T_2 = {reductionMux_io_o_data_0,reductionMux_io_o_data_1}; // @[Cat.scala 33:92]
  wire [1:0] _GEN_0 = 5'h0 == io_i_cmd ? 2'h0 : r_vn_valid; // @[EdgeAdderSwitch.scala 38:23 54:20 30:27]
  wire [63:0] _GEN_1 = 5'h5 == io_i_cmd ? _r_vn_T_2 : r_vn; // @[EdgeAdderSwitch.scala 38:23 50:14 29:21]
  wire [1:0] _GEN_2 = 5'h5 == io_i_cmd ? 2'h3 : _GEN_0; // @[EdgeAdderSwitch.scala 38:23 51:20]
  wire [31:0] _GEN_3 = 5'h4 == io_i_cmd ? reductionMux_io_o_data_0 : r_adder; // @[EdgeAdderSwitch.scala 38:23 45:17 28:24]
  wire [95:0] _GEN_4 = 5'h4 == io_i_cmd ? _r_vn_T_1 : {{32'd0}, _GEN_1}; // @[EdgeAdderSwitch.scala 38:23 46:14]
  wire [1:0] _GEN_5 = 5'h4 == io_i_cmd ? 2'h2 : _GEN_2; // @[EdgeAdderSwitch.scala 38:23 47:20]
  wire [95:0] _GEN_7 = 5'h3 == io_i_cmd ? _r_vn_T : _GEN_4; // @[EdgeAdderSwitch.scala 38:23 41:14]
  wire [95:0] _GEN_10 = r_valid ? _GEN_7 : {{32'd0}, r_vn}; // @[EdgeAdderSwitch.scala 29:21 37:25]
  wire [95:0] _GEN_13 = reset ? 96'h0 : _GEN_10; // @[EdgeAdderSwitch.scala 33:14 35:10]
  wire [31:0] _GEN_15 = r_add_en == 3'h0 ? r_adder : adder32_io_O; // @[EdgeAdderSwitch.scala 64:22 65:18 67:18]
  wire [95:0] _GEN_19 = reset ? 96'h0 : _GEN_13; // @[EdgeAdderSwitch.scala 29:{21,21}]
  ReductionMux_7 reductionMux ( // @[EdgeAdderSwitch.scala 19:28]
    .io_i_data_0(reductionMux_io_i_data_0),
    .io_i_data_1(reductionMux_io_i_data_1),
    .io_i_data_2(reductionMux_io_i_data_2),
    .io_i_data_3(reductionMux_io_i_data_3),
    .io_i_data_4(reductionMux_io_i_data_4),
    .io_i_data_5(reductionMux_io_i_data_5),
    .io_i_sel(reductionMux_io_i_sel),
    .io_o_data_0(reductionMux_io_o_data_0),
    .io_o_data_1(reductionMux_io_o_data_1)
  );
  SimpleAdder adder32 ( // @[EdgeAdderSwitch.scala 23:23]
    .io_A(adder32_io_A),
    .io_B(adder32_io_B),
    .io_O(adder32_io_O)
  );
  assign io_o_vn = reset ? 64'h0 : r_vn; // @[EdgeAdderSwitch.scala 59:14 61:13 69:13]
  assign io_o_vn_valid = reset ? 2'h0 : r_vn_valid; // @[EdgeAdderSwitch.scala 59:14 62:19 70:19]
  assign io_o_adder = reset ? 32'h0 : _GEN_15; // @[EdgeAdderSwitch.scala 59:14 60:16]
  assign reductionMux_io_i_data_0 = io_i_data_bus_0[31:0]; // @[EdgeAdderSwitch.scala 20:26]
  assign reductionMux_io_i_data_1 = io_i_data_bus_1[31:0]; // @[EdgeAdderSwitch.scala 20:26]
  assign reductionMux_io_i_data_2 = io_i_data_bus_2[31:0]; // @[EdgeAdderSwitch.scala 20:26]
  assign reductionMux_io_i_data_3 = io_i_data_bus_3[31:0]; // @[EdgeAdderSwitch.scala 20:26]
  assign reductionMux_io_i_data_4 = io_i_data_bus_4[31:0]; // @[EdgeAdderSwitch.scala 20:26]
  assign reductionMux_io_i_data_5 = io_i_data_bus_5[31:0]; // @[EdgeAdderSwitch.scala 20:26]
  assign reductionMux_io_i_sel = io_i_sel; // @[EdgeAdderSwitch.scala 21:25]
  assign adder32_io_A = reductionMux_io_o_data_1; // @[EdgeAdderSwitch.scala 24:16]
  assign adder32_io_B = reductionMux_io_o_data_0; // @[EdgeAdderSwitch.scala 25:16]
  always @(posedge clock) begin
    if (reset) begin // @[EdgeAdderSwitch.scala 27:24]
      r_valid <= 1'h0; // @[EdgeAdderSwitch.scala 27:24]
    end else begin
      r_valid <= io_i_valid; // @[EdgeAdderSwitch.scala 27:24]
    end
    if (reset) begin // @[EdgeAdderSwitch.scala 28:24]
      r_adder <= 32'h0; // @[EdgeAdderSwitch.scala 28:24]
    end else if (reset) begin // @[EdgeAdderSwitch.scala 33:14]
      r_adder <= 32'h0; // @[EdgeAdderSwitch.scala 34:13]
    end else if (r_valid) begin // @[EdgeAdderSwitch.scala 37:25]
      if (5'h3 == io_i_cmd) begin // @[EdgeAdderSwitch.scala 38:23]
        r_adder <= reductionMux_io_o_data_1; // @[EdgeAdderSwitch.scala 40:17]
      end else begin
        r_adder <= _GEN_3;
      end
    end
    r_vn <= _GEN_19[63:0]; // @[EdgeAdderSwitch.scala 29:{21,21}]
    if (reset) begin // @[EdgeAdderSwitch.scala 30:27]
      r_vn_valid <= 2'h0; // @[EdgeAdderSwitch.scala 30:27]
    end else if (reset) begin // @[EdgeAdderSwitch.scala 33:14]
      r_vn_valid <= 2'h0; // @[EdgeAdderSwitch.scala 36:16]
    end else if (r_valid) begin // @[EdgeAdderSwitch.scala 37:25]
      if (5'h3 == io_i_cmd) begin // @[EdgeAdderSwitch.scala 38:23]
        r_vn_valid <= 2'h1; // @[EdgeAdderSwitch.scala 42:20]
      end else begin
        r_vn_valid <= _GEN_5;
      end
    end
    if (reset) begin // @[EdgeAdderSwitch.scala 31:25]
      r_add_en <= 3'h0; // @[EdgeAdderSwitch.scala 31:25]
    end else begin
      r_add_en <= io_i_add_en; // @[EdgeAdderSwitch.scala 31:25]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  r_adder = _RAND_1[31:0];
  _RAND_2 = {2{`RANDOM}};
  r_vn = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  r_vn_valid = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  r_add_en = _RAND_4[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AdderSwitch_7(
  input         clock,
  input         reset,
  input         io_i_valid,
  input  [31:0] io_i_data_bus_0,
  input  [31:0] io_i_data_bus_1,
  input  [31:0] io_i_data_bus_2,
  input  [31:0] io_i_data_bus_3,
  input  [2:0]  io_i_add_en,
  input  [2:0]  io_i_cmd,
  input  [1:0]  io_i_sel,
  output [1:0]  io_o_vn_valid,
  output [63:0] io_o_vn,
  output [31:0] io_o_adder_0,
  output [31:0] io_o_adder_1
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] reductionMux_io_i_data_0; // @[AdderSwitch.scala 21:28]
  wire [31:0] reductionMux_io_i_data_1; // @[AdderSwitch.scala 21:28]
  wire [31:0] reductionMux_io_i_data_2; // @[AdderSwitch.scala 21:28]
  wire [31:0] reductionMux_io_i_data_3; // @[AdderSwitch.scala 21:28]
  wire [1:0] reductionMux_io_i_sel; // @[AdderSwitch.scala 21:28]
  wire [31:0] reductionMux_io_o_data_0; // @[AdderSwitch.scala 21:28]
  wire [31:0] reductionMux_io_o_data_1; // @[AdderSwitch.scala 21:28]
  wire [31:0] adder32_io_A; // @[AdderSwitch.scala 25:23]
  wire [31:0] adder32_io_B; // @[AdderSwitch.scala 25:23]
  wire [31:0] adder32_io_O; // @[AdderSwitch.scala 25:23]
  reg [63:0] r_adder; // @[AdderSwitch.scala 29:24]
  reg [63:0] r_vn; // @[AdderSwitch.scala 30:21]
  reg [1:0] r_vn_valid; // @[AdderSwitch.scala 31:27]
  reg [2:0] r_add_en; // @[AdderSwitch.scala 32:25]
  wire [63:0] _r_adder_T = {reductionMux_io_o_data_0,reductionMux_io_o_data_1}; // @[Cat.scala 33:92]
  wire [62:0] _r_adder_T_1 = {31'h0,reductionMux_io_o_data_1}; // @[Cat.scala 33:92]
  wire [62:0] _r_adder_T_2 = {reductionMux_io_o_data_0,31'h0}; // @[Cat.scala 33:92]
  wire [1:0] _GEN_0 = 3'h0 == io_i_cmd ? 2'h0 : r_vn_valid; // @[AdderSwitch.scala 39:23 59:20 31:27]
  wire [63:0] _GEN_1 = 3'h5 == io_i_cmd ? _r_adder_T : r_vn; // @[AdderSwitch.scala 39:23 55:14 30:21]
  wire [1:0] _GEN_2 = 3'h5 == io_i_cmd ? 2'h3 : _GEN_0; // @[AdderSwitch.scala 39:23 56:20]
  wire [63:0] _GEN_3 = 3'h4 == io_i_cmd ? {{1'd0}, _r_adder_T_2} : r_adder; // @[AdderSwitch.scala 39:23 50:17 29:24]
  wire [63:0] _GEN_4 = 3'h4 == io_i_cmd ? {{32'd0}, io_i_data_bus_1} : _GEN_1; // @[AdderSwitch.scala 39:23 51:14]
  wire [1:0] _GEN_5 = 3'h4 == io_i_cmd ? 2'h2 : _GEN_2; // @[AdderSwitch.scala 39:23 52:20]
  wire [63:0] _GEN_6 = 3'h3 == io_i_cmd ? {{1'd0}, _r_adder_T_1} : _GEN_3; // @[AdderSwitch.scala 39:23 45:17]
  wire [63:0] _GEN_7 = 3'h3 == io_i_cmd ? {{32'd0}, io_i_data_bus_0} : _GEN_4; // @[AdderSwitch.scala 39:23 46:14]
  wire [1:0] _GEN_8 = 3'h3 == io_i_cmd ? 2'h1 : _GEN_5; // @[AdderSwitch.scala 39:23 47:20]
  wire [31:0] _WIRE_2_0 = adder32_io_O; // @[AdderSwitch.scala 72:{28,28}]
  wire [31:0] _GEN_18 = r_add_en == 3'h0 ? r_adder[31:0] : _WIRE_2_0; // @[AdderSwitch.scala 69:22 70:18 72:18]
  wire [31:0] _GEN_19 = r_add_en == 3'h0 ? r_adder[63:32] : _WIRE_2_0; // @[AdderSwitch.scala 69:22 70:18 72:18]
  ReductionMux_3 reductionMux ( // @[AdderSwitch.scala 21:28]
    .io_i_data_0(reductionMux_io_i_data_0),
    .io_i_data_1(reductionMux_io_i_data_1),
    .io_i_data_2(reductionMux_io_i_data_2),
    .io_i_data_3(reductionMux_io_i_data_3),
    .io_i_sel(reductionMux_io_i_sel),
    .io_o_data_0(reductionMux_io_o_data_0),
    .io_o_data_1(reductionMux_io_o_data_1)
  );
  SimpleAdder adder32 ( // @[AdderSwitch.scala 25:23]
    .io_A(adder32_io_A),
    .io_B(adder32_io_B),
    .io_O(adder32_io_O)
  );
  assign io_o_vn_valid = reset ? 2'h0 : r_vn_valid; // @[AdderSwitch.scala 64:14 67:19 75:19]
  assign io_o_vn = reset ? 64'h0 : r_vn; // @[AdderSwitch.scala 64:14 66:13 74:13]
  assign io_o_adder_0 = reset ? 32'h0 : _GEN_18; // @[AdderSwitch.scala 64:14 65:16]
  assign io_o_adder_1 = reset ? 32'h0 : _GEN_19; // @[AdderSwitch.scala 64:14 65:16]
  assign reductionMux_io_i_data_0 = io_i_data_bus_0; // @[AdderSwitch.scala 22:26]
  assign reductionMux_io_i_data_1 = io_i_data_bus_1; // @[AdderSwitch.scala 22:26]
  assign reductionMux_io_i_data_2 = io_i_data_bus_2; // @[AdderSwitch.scala 22:26]
  assign reductionMux_io_i_data_3 = io_i_data_bus_3; // @[AdderSwitch.scala 22:26]
  assign reductionMux_io_i_sel = io_i_sel; // @[AdderSwitch.scala 23:25]
  assign adder32_io_A = reductionMux_io_o_data_1; // @[AdderSwitch.scala 26:16]
  assign adder32_io_B = reductionMux_io_o_data_0; // @[AdderSwitch.scala 27:16]
  always @(posedge clock) begin
    if (reset) begin // @[AdderSwitch.scala 29:24]
      r_adder <= 64'h0; // @[AdderSwitch.scala 29:24]
    end else if (reset) begin // @[AdderSwitch.scala 34:14]
      r_adder <= 64'h0; // @[AdderSwitch.scala 35:13]
    end else if (io_i_valid) begin // @[AdderSwitch.scala 38:28]
      if (3'h1 == io_i_cmd) begin // @[AdderSwitch.scala 39:23]
        r_adder <= _r_adder_T; // @[AdderSwitch.scala 41:17]
      end else begin
        r_adder <= _GEN_6;
      end
    end
    if (reset) begin // @[AdderSwitch.scala 30:21]
      r_vn <= 64'h0; // @[AdderSwitch.scala 30:21]
    end else if (reset) begin // @[AdderSwitch.scala 34:14]
      r_vn <= 64'h0; // @[AdderSwitch.scala 36:10]
    end else if (io_i_valid) begin // @[AdderSwitch.scala 38:28]
      if (!(3'h1 == io_i_cmd)) begin // @[AdderSwitch.scala 39:23]
        r_vn <= _GEN_7;
      end
    end
    if (reset) begin // @[AdderSwitch.scala 31:27]
      r_vn_valid <= 2'h0; // @[AdderSwitch.scala 31:27]
    end else if (reset) begin // @[AdderSwitch.scala 34:14]
      r_vn_valid <= 2'h0; // @[AdderSwitch.scala 37:16]
    end else if (io_i_valid) begin // @[AdderSwitch.scala 38:28]
      if (3'h1 == io_i_cmd) begin // @[AdderSwitch.scala 39:23]
        r_vn_valid <= 2'h0; // @[AdderSwitch.scala 42:20]
      end else begin
        r_vn_valid <= _GEN_8;
      end
    end
    if (reset) begin // @[AdderSwitch.scala 32:25]
      r_add_en <= 3'h0; // @[AdderSwitch.scala 32:25]
    end else begin
      r_add_en <= io_i_add_en; // @[AdderSwitch.scala 32:25]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  r_adder = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  r_vn = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  r_vn_valid = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  r_add_en = _RAND_3[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ReductionMux_15(
  input  [31:0] io_i_data_0,
  input  [31:0] io_i_data_1,
  input  [31:0] io_i_data_2,
  input  [31:0] io_i_data_3,
  input  [31:0] io_i_data_4,
  input  [31:0] io_i_data_5,
  input  [31:0] io_i_data_6,
  input  [31:0] io_i_data_7,
  input  [3:0]  io_i_sel,
  output [31:0] io_o_data_0,
  output [31:0] io_o_data_1
);
  wire [1:0] w_sel_in_left = io_i_sel[1:0]; // @[ReductionMux.scala 28:32]
  wire [1:0] w_sel_in_right = io_i_sel[3:2]; // @[ReductionMux.scala 29:33]
  wire [31:0] _GEN_1 = 2'h1 == w_sel_in_left ? io_i_data_1 : io_i_data_0; // @[ReductionMux.scala 33:{18,18}]
  wire [31:0] _GEN_2 = 2'h2 == w_sel_in_left ? io_i_data_2 : _GEN_1; // @[ReductionMux.scala 33:{18,18}]
  wire [31:0] _GEN_3 = 2'h3 == w_sel_in_left ? io_i_data_3 : _GEN_2; // @[ReductionMux.scala 33:{18,18}]
  wire [31:0] _GEN_6 = 2'h1 == w_sel_in_right ? io_i_data_5 : io_i_data_4; // @[ReductionMux.scala 37:{22,22}]
  wire [31:0] _GEN_7 = 2'h2 == w_sel_in_right ? io_i_data_6 : _GEN_6; // @[ReductionMux.scala 37:{22,22}]
  assign io_o_data_0 = w_sel_in_left < 2'h2 ? _GEN_3 : 32'h0; // @[ReductionMux.scala 31:39 33:18 35:18]
  assign io_o_data_1 = 2'h3 == w_sel_in_right ? io_i_data_7 : _GEN_7; // @[ReductionMux.scala 37:{22,22}]
endmodule
module EdgeAdderSwitch_4(
  input         clock,
  input         reset,
  input         io_i_valid,
  input  [63:0] io_i_data_bus_0,
  input  [63:0] io_i_data_bus_1,
  input  [63:0] io_i_data_bus_2,
  input  [63:0] io_i_data_bus_3,
  input  [63:0] io_i_data_bus_4,
  input  [63:0] io_i_data_bus_5,
  input  [63:0] io_i_data_bus_6,
  input  [63:0] io_i_data_bus_7,
  input  [2:0]  io_i_add_en,
  input  [4:0]  io_i_cmd,
  input  [3:0]  io_i_sel,
  output [63:0] io_o_vn,
  output [1:0]  io_o_vn_valid,
  output [31:0] io_o_adder
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] reductionMux_io_i_data_0; // @[EdgeAdderSwitch.scala 19:28]
  wire [31:0] reductionMux_io_i_data_1; // @[EdgeAdderSwitch.scala 19:28]
  wire [31:0] reductionMux_io_i_data_2; // @[EdgeAdderSwitch.scala 19:28]
  wire [31:0] reductionMux_io_i_data_3; // @[EdgeAdderSwitch.scala 19:28]
  wire [31:0] reductionMux_io_i_data_4; // @[EdgeAdderSwitch.scala 19:28]
  wire [31:0] reductionMux_io_i_data_5; // @[EdgeAdderSwitch.scala 19:28]
  wire [31:0] reductionMux_io_i_data_6; // @[EdgeAdderSwitch.scala 19:28]
  wire [31:0] reductionMux_io_i_data_7; // @[EdgeAdderSwitch.scala 19:28]
  wire [3:0] reductionMux_io_i_sel; // @[EdgeAdderSwitch.scala 19:28]
  wire [31:0] reductionMux_io_o_data_0; // @[EdgeAdderSwitch.scala 19:28]
  wire [31:0] reductionMux_io_o_data_1; // @[EdgeAdderSwitch.scala 19:28]
  wire [31:0] adder32_io_A; // @[EdgeAdderSwitch.scala 23:23]
  wire [31:0] adder32_io_B; // @[EdgeAdderSwitch.scala 23:23]
  wire [31:0] adder32_io_O; // @[EdgeAdderSwitch.scala 23:23]
  reg  r_valid; // @[EdgeAdderSwitch.scala 27:24]
  reg [31:0] r_adder; // @[EdgeAdderSwitch.scala 28:24]
  reg [63:0] r_vn; // @[EdgeAdderSwitch.scala 29:21]
  reg [1:0] r_vn_valid; // @[EdgeAdderSwitch.scala 30:27]
  reg [2:0] r_add_en; // @[EdgeAdderSwitch.scala 31:25]
  wire [95:0] _r_vn_T = {io_i_data_bus_0,32'h0}; // @[Cat.scala 33:92]
  wire [95:0] _r_vn_T_1 = {32'h0,io_i_data_bus_7}; // @[Cat.scala 33:92]
  wire [63:0] _r_vn_T_2 = {reductionMux_io_o_data_0,reductionMux_io_o_data_1}; // @[Cat.scala 33:92]
  wire [1:0] _GEN_0 = 5'h0 == io_i_cmd ? 2'h0 : r_vn_valid; // @[EdgeAdderSwitch.scala 38:23 54:20 30:27]
  wire [63:0] _GEN_1 = 5'h5 == io_i_cmd ? _r_vn_T_2 : r_vn; // @[EdgeAdderSwitch.scala 38:23 50:14 29:21]
  wire [1:0] _GEN_2 = 5'h5 == io_i_cmd ? 2'h3 : _GEN_0; // @[EdgeAdderSwitch.scala 38:23 51:20]
  wire [31:0] _GEN_3 = 5'h4 == io_i_cmd ? reductionMux_io_o_data_0 : r_adder; // @[EdgeAdderSwitch.scala 38:23 45:17 28:24]
  wire [95:0] _GEN_4 = 5'h4 == io_i_cmd ? _r_vn_T_1 : {{32'd0}, _GEN_1}; // @[EdgeAdderSwitch.scala 38:23 46:14]
  wire [1:0] _GEN_5 = 5'h4 == io_i_cmd ? 2'h2 : _GEN_2; // @[EdgeAdderSwitch.scala 38:23 47:20]
  wire [95:0] _GEN_7 = 5'h3 == io_i_cmd ? _r_vn_T : _GEN_4; // @[EdgeAdderSwitch.scala 38:23 41:14]
  wire [95:0] _GEN_10 = r_valid ? _GEN_7 : {{32'd0}, r_vn}; // @[EdgeAdderSwitch.scala 29:21 37:25]
  wire [95:0] _GEN_13 = reset ? 96'h0 : _GEN_10; // @[EdgeAdderSwitch.scala 33:14 35:10]
  wire [31:0] _GEN_15 = r_add_en == 3'h0 ? r_adder : adder32_io_O; // @[EdgeAdderSwitch.scala 64:22 65:18 67:18]
  wire [95:0] _GEN_19 = reset ? 96'h0 : _GEN_13; // @[EdgeAdderSwitch.scala 29:{21,21}]
  ReductionMux_15 reductionMux ( // @[EdgeAdderSwitch.scala 19:28]
    .io_i_data_0(reductionMux_io_i_data_0),
    .io_i_data_1(reductionMux_io_i_data_1),
    .io_i_data_2(reductionMux_io_i_data_2),
    .io_i_data_3(reductionMux_io_i_data_3),
    .io_i_data_4(reductionMux_io_i_data_4),
    .io_i_data_5(reductionMux_io_i_data_5),
    .io_i_data_6(reductionMux_io_i_data_6),
    .io_i_data_7(reductionMux_io_i_data_7),
    .io_i_sel(reductionMux_io_i_sel),
    .io_o_data_0(reductionMux_io_o_data_0),
    .io_o_data_1(reductionMux_io_o_data_1)
  );
  SimpleAdder adder32 ( // @[EdgeAdderSwitch.scala 23:23]
    .io_A(adder32_io_A),
    .io_B(adder32_io_B),
    .io_O(adder32_io_O)
  );
  assign io_o_vn = reset ? 64'h0 : r_vn; // @[EdgeAdderSwitch.scala 59:14 61:13 69:13]
  assign io_o_vn_valid = reset ? 2'h0 : r_vn_valid; // @[EdgeAdderSwitch.scala 59:14 62:19 70:19]
  assign io_o_adder = reset ? 32'h0 : _GEN_15; // @[EdgeAdderSwitch.scala 59:14 60:16]
  assign reductionMux_io_i_data_0 = io_i_data_bus_0[31:0]; // @[EdgeAdderSwitch.scala 20:26]
  assign reductionMux_io_i_data_1 = io_i_data_bus_1[31:0]; // @[EdgeAdderSwitch.scala 20:26]
  assign reductionMux_io_i_data_2 = io_i_data_bus_2[31:0]; // @[EdgeAdderSwitch.scala 20:26]
  assign reductionMux_io_i_data_3 = io_i_data_bus_3[31:0]; // @[EdgeAdderSwitch.scala 20:26]
  assign reductionMux_io_i_data_4 = io_i_data_bus_4[31:0]; // @[EdgeAdderSwitch.scala 20:26]
  assign reductionMux_io_i_data_5 = io_i_data_bus_5[31:0]; // @[EdgeAdderSwitch.scala 20:26]
  assign reductionMux_io_i_data_6 = io_i_data_bus_6[31:0]; // @[EdgeAdderSwitch.scala 20:26]
  assign reductionMux_io_i_data_7 = io_i_data_bus_7[31:0]; // @[EdgeAdderSwitch.scala 20:26]
  assign reductionMux_io_i_sel = io_i_sel; // @[EdgeAdderSwitch.scala 21:25]
  assign adder32_io_A = reductionMux_io_o_data_1; // @[EdgeAdderSwitch.scala 24:16]
  assign adder32_io_B = reductionMux_io_o_data_0; // @[EdgeAdderSwitch.scala 25:16]
  always @(posedge clock) begin
    if (reset) begin // @[EdgeAdderSwitch.scala 27:24]
      r_valid <= 1'h0; // @[EdgeAdderSwitch.scala 27:24]
    end else begin
      r_valid <= io_i_valid; // @[EdgeAdderSwitch.scala 27:24]
    end
    if (reset) begin // @[EdgeAdderSwitch.scala 28:24]
      r_adder <= 32'h0; // @[EdgeAdderSwitch.scala 28:24]
    end else if (reset) begin // @[EdgeAdderSwitch.scala 33:14]
      r_adder <= 32'h0; // @[EdgeAdderSwitch.scala 34:13]
    end else if (r_valid) begin // @[EdgeAdderSwitch.scala 37:25]
      if (5'h3 == io_i_cmd) begin // @[EdgeAdderSwitch.scala 38:23]
        r_adder <= reductionMux_io_o_data_1; // @[EdgeAdderSwitch.scala 40:17]
      end else begin
        r_adder <= _GEN_3;
      end
    end
    r_vn <= _GEN_19[63:0]; // @[EdgeAdderSwitch.scala 29:{21,21}]
    if (reset) begin // @[EdgeAdderSwitch.scala 30:27]
      r_vn_valid <= 2'h0; // @[EdgeAdderSwitch.scala 30:27]
    end else if (reset) begin // @[EdgeAdderSwitch.scala 33:14]
      r_vn_valid <= 2'h0; // @[EdgeAdderSwitch.scala 36:16]
    end else if (r_valid) begin // @[EdgeAdderSwitch.scala 37:25]
      if (5'h3 == io_i_cmd) begin // @[EdgeAdderSwitch.scala 38:23]
        r_vn_valid <= 2'h1; // @[EdgeAdderSwitch.scala 42:20]
      end else begin
        r_vn_valid <= _GEN_5;
      end
    end
    if (reset) begin // @[EdgeAdderSwitch.scala 31:25]
      r_add_en <= 3'h0; // @[EdgeAdderSwitch.scala 31:25]
    end else begin
      r_add_en <= io_i_add_en; // @[EdgeAdderSwitch.scala 31:25]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  r_adder = _RAND_1[31:0];
  _RAND_2 = {2{`RANDOM}};
  r_vn = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  r_vn_valid = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  r_add_en = _RAND_4[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FanNetworkcom(
  input         clock,
  input         reset,
  input         io_i_valid,
  input  [31:0] io_i_data_bus_0,
  input  [31:0] io_i_data_bus_1,
  input  [31:0] io_i_data_bus_2,
  input  [31:0] io_i_data_bus_3,
  input  [31:0] io_i_data_bus_4,
  input  [31:0] io_i_data_bus_5,
  input  [31:0] io_i_data_bus_6,
  input  [31:0] io_i_data_bus_7,
  input  [31:0] io_i_data_bus_8,
  input  [31:0] io_i_data_bus_9,
  input  [31:0] io_i_data_bus_10,
  input  [31:0] io_i_data_bus_11,
  input  [31:0] io_i_data_bus_12,
  input  [31:0] io_i_data_bus_13,
  input  [31:0] io_i_data_bus_14,
  input  [31:0] io_i_data_bus_15,
  input  [31:0] io_i_data_bus_16,
  input  [31:0] io_i_data_bus_17,
  input  [31:0] io_i_data_bus_18,
  input  [31:0] io_i_data_bus_19,
  input  [31:0] io_i_data_bus_20,
  input  [31:0] io_i_data_bus_21,
  input  [31:0] io_i_data_bus_22,
  input  [31:0] io_i_data_bus_23,
  input  [31:0] io_i_data_bus_24,
  input  [31:0] io_i_data_bus_25,
  input  [31:0] io_i_data_bus_26,
  input  [31:0] io_i_data_bus_27,
  input  [31:0] io_i_data_bus_28,
  input  [31:0] io_i_data_bus_29,
  input  [31:0] io_i_data_bus_30,
  input  [31:0] io_i_data_bus_31,
  input         io_i_add_en_bus_0,
  input         io_i_add_en_bus_1,
  input         io_i_add_en_bus_2,
  input         io_i_add_en_bus_3,
  input         io_i_add_en_bus_4,
  input         io_i_add_en_bus_5,
  input         io_i_add_en_bus_6,
  input         io_i_add_en_bus_7,
  input         io_i_add_en_bus_8,
  input         io_i_add_en_bus_9,
  input         io_i_add_en_bus_10,
  input         io_i_add_en_bus_11,
  input         io_i_add_en_bus_12,
  input         io_i_add_en_bus_13,
  input         io_i_add_en_bus_14,
  input         io_i_add_en_bus_15,
  input         io_i_add_en_bus_16,
  input         io_i_add_en_bus_17,
  input         io_i_add_en_bus_18,
  input         io_i_add_en_bus_19,
  input         io_i_add_en_bus_20,
  input         io_i_add_en_bus_21,
  input         io_i_add_en_bus_22,
  input         io_i_add_en_bus_23,
  input         io_i_add_en_bus_24,
  input         io_i_add_en_bus_25,
  input         io_i_add_en_bus_26,
  input         io_i_add_en_bus_27,
  input         io_i_add_en_bus_28,
  input         io_i_add_en_bus_29,
  input         io_i_add_en_bus_30,
  input  [2:0]  io_i_cmd_bus_0,
  input  [2:0]  io_i_cmd_bus_1,
  input  [2:0]  io_i_cmd_bus_2,
  input  [2:0]  io_i_cmd_bus_3,
  input  [2:0]  io_i_cmd_bus_4,
  input  [2:0]  io_i_cmd_bus_5,
  input  [2:0]  io_i_cmd_bus_6,
  input  [2:0]  io_i_cmd_bus_7,
  input  [2:0]  io_i_cmd_bus_8,
  input  [2:0]  io_i_cmd_bus_9,
  input  [2:0]  io_i_cmd_bus_10,
  input  [2:0]  io_i_cmd_bus_11,
  input  [2:0]  io_i_cmd_bus_12,
  input  [2:0]  io_i_cmd_bus_13,
  input  [2:0]  io_i_cmd_bus_14,
  input  [2:0]  io_i_cmd_bus_15,
  input  [2:0]  io_i_cmd_bus_16,
  input  [2:0]  io_i_cmd_bus_17,
  input  [2:0]  io_i_cmd_bus_18,
  input  [2:0]  io_i_cmd_bus_19,
  input  [2:0]  io_i_cmd_bus_20,
  input  [2:0]  io_i_cmd_bus_21,
  input  [2:0]  io_i_cmd_bus_22,
  input  [2:0]  io_i_cmd_bus_23,
  input  [2:0]  io_i_cmd_bus_24,
  input  [2:0]  io_i_cmd_bus_25,
  input  [2:0]  io_i_cmd_bus_26,
  input  [2:0]  io_i_cmd_bus_27,
  input  [2:0]  io_i_cmd_bus_28,
  input  [2:0]  io_i_cmd_bus_29,
  input  [2:0]  io_i_cmd_bus_30,
  input  [1:0]  io_i_sel_bus_0,
  input  [1:0]  io_i_sel_bus_1,
  input  [1:0]  io_i_sel_bus_2,
  input  [1:0]  io_i_sel_bus_3,
  input  [1:0]  io_i_sel_bus_4,
  input  [1:0]  io_i_sel_bus_5,
  input  [1:0]  io_i_sel_bus_6,
  input  [1:0]  io_i_sel_bus_7,
  input  [1:0]  io_i_sel_bus_8,
  input  [1:0]  io_i_sel_bus_9,
  input  [1:0]  io_i_sel_bus_10,
  input  [1:0]  io_i_sel_bus_11,
  input  [1:0]  io_i_sel_bus_12,
  input  [1:0]  io_i_sel_bus_13,
  input  [1:0]  io_i_sel_bus_14,
  input  [1:0]  io_i_sel_bus_15,
  input  [1:0]  io_i_sel_bus_16,
  input  [1:0]  io_i_sel_bus_17,
  input  [1:0]  io_i_sel_bus_18,
  input  [1:0]  io_i_sel_bus_19,
  output        io_o_valid_0,
  output        io_o_valid_1,
  output        io_o_valid_2,
  output        io_o_valid_3,
  output        io_o_valid_4,
  output        io_o_valid_5,
  output        io_o_valid_6,
  output        io_o_valid_7,
  output        io_o_valid_8,
  output        io_o_valid_9,
  output        io_o_valid_10,
  output        io_o_valid_11,
  output        io_o_valid_12,
  output        io_o_valid_13,
  output        io_o_valid_14,
  output        io_o_valid_15,
  output        io_o_valid_16,
  output        io_o_valid_17,
  output        io_o_valid_18,
  output        io_o_valid_19,
  output        io_o_valid_20,
  output        io_o_valid_21,
  output        io_o_valid_22,
  output        io_o_valid_23,
  output        io_o_valid_24,
  output        io_o_valid_25,
  output        io_o_valid_26,
  output        io_o_valid_27,
  output        io_o_valid_28,
  output        io_o_valid_29,
  output        io_o_valid_30,
  output        io_o_valid_31,
  output [31:0] io_o_data_bus_0,
  output [31:0] io_o_data_bus_1,
  output [31:0] io_o_data_bus_2,
  output [31:0] io_o_data_bus_3,
  output [31:0] io_o_data_bus_4,
  output [31:0] io_o_data_bus_5,
  output [31:0] io_o_data_bus_6,
  output [31:0] io_o_data_bus_7,
  output [31:0] io_o_data_bus_8,
  output [31:0] io_o_data_bus_9,
  output [31:0] io_o_data_bus_10,
  output [31:0] io_o_data_bus_11,
  output [31:0] io_o_data_bus_12,
  output [31:0] io_o_data_bus_13,
  output [31:0] io_o_data_bus_14,
  output [31:0] io_o_data_bus_15,
  output [31:0] io_o_data_bus_16,
  output [31:0] io_o_data_bus_17,
  output [31:0] io_o_data_bus_18,
  output [31:0] io_o_data_bus_19,
  output [31:0] io_o_data_bus_20,
  output [31:0] io_o_data_bus_21,
  output [31:0] io_o_data_bus_22,
  output [31:0] io_o_data_bus_23,
  output [31:0] io_o_data_bus_24,
  output [31:0] io_o_data_bus_25,
  output [31:0] io_o_data_bus_26,
  output [31:0] io_o_data_bus_27,
  output [31:0] io_o_data_bus_28,
  output [31:0] io_o_data_bus_29,
  output [31:0] io_o_data_bus_30,
  output [31:0] io_o_data_bus_31,
  output [31:0] io_o_adder_0,
  output [31:0] io_o_adder_1,
  output [31:0] io_o_adder_2,
  output [31:0] io_o_adder_3,
  output [31:0] io_o_adder_4,
  output [31:0] io_o_adder_5,
  output [31:0] io_o_adder_6,
  output [31:0] io_o_adder_7,
  output [31:0] io_o_adder_8,
  output [31:0] io_o_adder_9,
  output [31:0] io_o_adder_10,
  output [31:0] io_o_adder_11,
  output [31:0] io_o_adder_12,
  output [31:0] io_o_adder_13,
  output [31:0] io_o_adder_14,
  output [31:0] io_o_adder_15,
  output [31:0] io_o_adder_16,
  output [31:0] io_o_adder_17,
  output [31:0] io_o_adder_18,
  output [31:0] io_o_adder_19,
  output [31:0] io_o_adder_20,
  output [31:0] io_o_adder_21,
  output [31:0] io_o_adder_22,
  output [31:0] io_o_adder_23,
  output [31:0] io_o_adder_24,
  output [31:0] io_o_adder_25,
  output [31:0] io_o_adder_26,
  output [31:0] io_o_adder_27,
  output [31:0] io_o_adder_28,
  output [31:0] io_o_adder_29,
  output [31:0] io_o_adder_30
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
`endif // RANDOMIZE_REG_INIT
  wire  my_adder_0_clock; // @[FanNetwork.scala 984:28]
  wire  my_adder_0_reset; // @[FanNetwork.scala 984:28]
  wire  my_adder_0_io_i_valid; // @[FanNetwork.scala 984:28]
  wire [63:0] my_adder_0_io_i_data_bus_0; // @[FanNetwork.scala 984:28]
  wire [63:0] my_adder_0_io_i_data_bus_1; // @[FanNetwork.scala 984:28]
  wire [2:0] my_adder_0_io_i_add_en; // @[FanNetwork.scala 984:28]
  wire [4:0] my_adder_0_io_i_cmd; // @[FanNetwork.scala 984:28]
  wire [63:0] my_adder_0_io_o_vn; // @[FanNetwork.scala 984:28]
  wire [1:0] my_adder_0_io_o_vn_valid; // @[FanNetwork.scala 984:28]
  wire [31:0] my_adder_0_io_o_adder; // @[FanNetwork.scala 984:28]
  wire  my_adder_1_clock; // @[FanNetwork.scala 997:28]
  wire  my_adder_1_reset; // @[FanNetwork.scala 997:28]
  wire  my_adder_1_io_i_valid; // @[FanNetwork.scala 997:28]
  wire [63:0] my_adder_1_io_i_data_bus_0; // @[FanNetwork.scala 997:28]
  wire [63:0] my_adder_1_io_i_data_bus_1; // @[FanNetwork.scala 997:28]
  wire [2:0] my_adder_1_io_i_add_en; // @[FanNetwork.scala 997:28]
  wire [4:0] my_adder_1_io_i_cmd; // @[FanNetwork.scala 997:28]
  wire [63:0] my_adder_1_io_o_vn; // @[FanNetwork.scala 997:28]
  wire [1:0] my_adder_1_io_o_vn_valid; // @[FanNetwork.scala 997:28]
  wire [31:0] my_adder_1_io_o_adder; // @[FanNetwork.scala 997:28]
  wire  my_adder_2_clock; // @[FanNetwork.scala 1010:28]
  wire  my_adder_2_reset; // @[FanNetwork.scala 1010:28]
  wire  my_adder_2_io_i_valid; // @[FanNetwork.scala 1010:28]
  wire [31:0] my_adder_2_io_i_data_bus_0; // @[FanNetwork.scala 1010:28]
  wire [31:0] my_adder_2_io_i_data_bus_1; // @[FanNetwork.scala 1010:28]
  wire [2:0] my_adder_2_io_i_add_en; // @[FanNetwork.scala 1010:28]
  wire [2:0] my_adder_2_io_i_cmd; // @[FanNetwork.scala 1010:28]
  wire [1:0] my_adder_2_io_o_vn_valid; // @[FanNetwork.scala 1010:28]
  wire [63:0] my_adder_2_io_o_vn; // @[FanNetwork.scala 1010:28]
  wire [31:0] my_adder_2_io_o_adder_0; // @[FanNetwork.scala 1010:28]
  wire [31:0] my_adder_2_io_o_adder_1; // @[FanNetwork.scala 1010:28]
  wire  my_adder_3_clock; // @[FanNetwork.scala 1028:28]
  wire  my_adder_3_reset; // @[FanNetwork.scala 1028:28]
  wire  my_adder_3_io_i_valid; // @[FanNetwork.scala 1028:28]
  wire [63:0] my_adder_3_io_i_data_bus_0; // @[FanNetwork.scala 1028:28]
  wire [63:0] my_adder_3_io_i_data_bus_1; // @[FanNetwork.scala 1028:28]
  wire [63:0] my_adder_3_io_i_data_bus_2; // @[FanNetwork.scala 1028:28]
  wire [63:0] my_adder_3_io_i_data_bus_3; // @[FanNetwork.scala 1028:28]
  wire [2:0] my_adder_3_io_i_add_en; // @[FanNetwork.scala 1028:28]
  wire [4:0] my_adder_3_io_i_cmd; // @[FanNetwork.scala 1028:28]
  wire [1:0] my_adder_3_io_i_sel; // @[FanNetwork.scala 1028:28]
  wire [63:0] my_adder_3_io_o_vn; // @[FanNetwork.scala 1028:28]
  wire [1:0] my_adder_3_io_o_vn_valid; // @[FanNetwork.scala 1028:28]
  wire [31:0] my_adder_3_io_o_adder; // @[FanNetwork.scala 1028:28]
  wire  my_adder_4_clock; // @[FanNetwork.scala 1043:28]
  wire  my_adder_4_reset; // @[FanNetwork.scala 1043:28]
  wire  my_adder_4_io_i_valid; // @[FanNetwork.scala 1043:28]
  wire [31:0] my_adder_4_io_i_data_bus_0; // @[FanNetwork.scala 1043:28]
  wire [31:0] my_adder_4_io_i_data_bus_1; // @[FanNetwork.scala 1043:28]
  wire [2:0] my_adder_4_io_i_add_en; // @[FanNetwork.scala 1043:28]
  wire [2:0] my_adder_4_io_i_cmd; // @[FanNetwork.scala 1043:28]
  wire [1:0] my_adder_4_io_o_vn_valid; // @[FanNetwork.scala 1043:28]
  wire [63:0] my_adder_4_io_o_vn; // @[FanNetwork.scala 1043:28]
  wire [31:0] my_adder_4_io_o_adder_0; // @[FanNetwork.scala 1043:28]
  wire [31:0] my_adder_4_io_o_adder_1; // @[FanNetwork.scala 1043:28]
  wire  my_adder_5_clock; // @[FanNetwork.scala 1060:28]
  wire  my_adder_5_reset; // @[FanNetwork.scala 1060:28]
  wire  my_adder_5_io_i_valid; // @[FanNetwork.scala 1060:28]
  wire [31:0] my_adder_5_io_i_data_bus_0; // @[FanNetwork.scala 1060:28]
  wire [31:0] my_adder_5_io_i_data_bus_1; // @[FanNetwork.scala 1060:28]
  wire [2:0] my_adder_5_io_i_add_en; // @[FanNetwork.scala 1060:28]
  wire [2:0] my_adder_5_io_i_cmd; // @[FanNetwork.scala 1060:28]
  wire [1:0] my_adder_5_io_o_vn_valid; // @[FanNetwork.scala 1060:28]
  wire [63:0] my_adder_5_io_o_vn; // @[FanNetwork.scala 1060:28]
  wire [31:0] my_adder_5_io_o_adder_0; // @[FanNetwork.scala 1060:28]
  wire [31:0] my_adder_5_io_o_adder_1; // @[FanNetwork.scala 1060:28]
  wire  my_adder_6_clock; // @[FanNetwork.scala 1076:28]
  wire  my_adder_6_reset; // @[FanNetwork.scala 1076:28]
  wire  my_adder_6_io_i_valid; // @[FanNetwork.scala 1076:28]
  wire [31:0] my_adder_6_io_i_data_bus_0; // @[FanNetwork.scala 1076:28]
  wire [31:0] my_adder_6_io_i_data_bus_1; // @[FanNetwork.scala 1076:28]
  wire [2:0] my_adder_6_io_i_add_en; // @[FanNetwork.scala 1076:28]
  wire [2:0] my_adder_6_io_i_cmd; // @[FanNetwork.scala 1076:28]
  wire [1:0] my_adder_6_io_o_vn_valid; // @[FanNetwork.scala 1076:28]
  wire [63:0] my_adder_6_io_o_vn; // @[FanNetwork.scala 1076:28]
  wire [31:0] my_adder_6_io_o_adder_0; // @[FanNetwork.scala 1076:28]
  wire [31:0] my_adder_6_io_o_adder_1; // @[FanNetwork.scala 1076:28]
  wire  my_adder_7_clock; // @[FanNetwork.scala 1092:28]
  wire  my_adder_7_reset; // @[FanNetwork.scala 1092:28]
  wire  my_adder_7_io_i_valid; // @[FanNetwork.scala 1092:28]
  wire [63:0] my_adder_7_io_i_data_bus_0; // @[FanNetwork.scala 1092:28]
  wire [63:0] my_adder_7_io_i_data_bus_1; // @[FanNetwork.scala 1092:28]
  wire [63:0] my_adder_7_io_i_data_bus_2; // @[FanNetwork.scala 1092:28]
  wire [63:0] my_adder_7_io_i_data_bus_3; // @[FanNetwork.scala 1092:28]
  wire [63:0] my_adder_7_io_i_data_bus_4; // @[FanNetwork.scala 1092:28]
  wire [63:0] my_adder_7_io_i_data_bus_5; // @[FanNetwork.scala 1092:28]
  wire [2:0] my_adder_7_io_i_add_en; // @[FanNetwork.scala 1092:28]
  wire [4:0] my_adder_7_io_i_cmd; // @[FanNetwork.scala 1092:28]
  wire [3:0] my_adder_7_io_i_sel; // @[FanNetwork.scala 1092:28]
  wire [63:0] my_adder_7_io_o_vn; // @[FanNetwork.scala 1092:28]
  wire [1:0] my_adder_7_io_o_vn_valid; // @[FanNetwork.scala 1092:28]
  wire [31:0] my_adder_7_io_o_adder; // @[FanNetwork.scala 1092:28]
  wire  my_adder_8_clock; // @[FanNetwork.scala 1109:28]
  wire  my_adder_8_reset; // @[FanNetwork.scala 1109:28]
  wire  my_adder_8_io_i_valid; // @[FanNetwork.scala 1109:28]
  wire [31:0] my_adder_8_io_i_data_bus_0; // @[FanNetwork.scala 1109:28]
  wire [31:0] my_adder_8_io_i_data_bus_1; // @[FanNetwork.scala 1109:28]
  wire [2:0] my_adder_8_io_i_add_en; // @[FanNetwork.scala 1109:28]
  wire [2:0] my_adder_8_io_i_cmd; // @[FanNetwork.scala 1109:28]
  wire [1:0] my_adder_8_io_o_vn_valid; // @[FanNetwork.scala 1109:28]
  wire [63:0] my_adder_8_io_o_vn; // @[FanNetwork.scala 1109:28]
  wire [31:0] my_adder_8_io_o_adder_0; // @[FanNetwork.scala 1109:28]
  wire [31:0] my_adder_8_io_o_adder_1; // @[FanNetwork.scala 1109:28]
  wire  my_adder_9_clock; // @[FanNetwork.scala 1125:28]
  wire  my_adder_9_reset; // @[FanNetwork.scala 1125:28]
  wire  my_adder_9_io_i_valid; // @[FanNetwork.scala 1125:28]
  wire [31:0] my_adder_9_io_i_data_bus_0; // @[FanNetwork.scala 1125:28]
  wire [31:0] my_adder_9_io_i_data_bus_1; // @[FanNetwork.scala 1125:28]
  wire [2:0] my_adder_9_io_i_add_en; // @[FanNetwork.scala 1125:28]
  wire [2:0] my_adder_9_io_i_cmd; // @[FanNetwork.scala 1125:28]
  wire [1:0] my_adder_9_io_o_vn_valid; // @[FanNetwork.scala 1125:28]
  wire [63:0] my_adder_9_io_o_vn; // @[FanNetwork.scala 1125:28]
  wire [31:0] my_adder_9_io_o_adder_0; // @[FanNetwork.scala 1125:28]
  wire [31:0] my_adder_9_io_o_adder_1; // @[FanNetwork.scala 1125:28]
  wire  my_adder_10_clock; // @[FanNetwork.scala 1141:29]
  wire  my_adder_10_reset; // @[FanNetwork.scala 1141:29]
  wire  my_adder_10_io_i_valid; // @[FanNetwork.scala 1141:29]
  wire [31:0] my_adder_10_io_i_data_bus_0; // @[FanNetwork.scala 1141:29]
  wire [31:0] my_adder_10_io_i_data_bus_1; // @[FanNetwork.scala 1141:29]
  wire [2:0] my_adder_10_io_i_add_en; // @[FanNetwork.scala 1141:29]
  wire [2:0] my_adder_10_io_i_cmd; // @[FanNetwork.scala 1141:29]
  wire [1:0] my_adder_10_io_o_vn_valid; // @[FanNetwork.scala 1141:29]
  wire [63:0] my_adder_10_io_o_vn; // @[FanNetwork.scala 1141:29]
  wire [31:0] my_adder_10_io_o_adder_0; // @[FanNetwork.scala 1141:29]
  wire [31:0] my_adder_10_io_o_adder_1; // @[FanNetwork.scala 1141:29]
  wire  my_adder_11_clock; // @[FanNetwork.scala 1158:29]
  wire  my_adder_11_reset; // @[FanNetwork.scala 1158:29]
  wire  my_adder_11_io_i_valid; // @[FanNetwork.scala 1158:29]
  wire [31:0] my_adder_11_io_i_data_bus_0; // @[FanNetwork.scala 1158:29]
  wire [31:0] my_adder_11_io_i_data_bus_1; // @[FanNetwork.scala 1158:29]
  wire [31:0] my_adder_11_io_i_data_bus_2; // @[FanNetwork.scala 1158:29]
  wire [31:0] my_adder_11_io_i_data_bus_3; // @[FanNetwork.scala 1158:29]
  wire [2:0] my_adder_11_io_i_add_en; // @[FanNetwork.scala 1158:29]
  wire [2:0] my_adder_11_io_i_cmd; // @[FanNetwork.scala 1158:29]
  wire [1:0] my_adder_11_io_i_sel; // @[FanNetwork.scala 1158:29]
  wire [1:0] my_adder_11_io_o_vn_valid; // @[FanNetwork.scala 1158:29]
  wire [63:0] my_adder_11_io_o_vn; // @[FanNetwork.scala 1158:29]
  wire [31:0] my_adder_11_io_o_adder_0; // @[FanNetwork.scala 1158:29]
  wire [31:0] my_adder_11_io_o_adder_1; // @[FanNetwork.scala 1158:29]
  wire  my_adder_12_clock; // @[FanNetwork.scala 1177:29]
  wire  my_adder_12_reset; // @[FanNetwork.scala 1177:29]
  wire  my_adder_12_io_i_valid; // @[FanNetwork.scala 1177:29]
  wire [31:0] my_adder_12_io_i_data_bus_0; // @[FanNetwork.scala 1177:29]
  wire [31:0] my_adder_12_io_i_data_bus_1; // @[FanNetwork.scala 1177:29]
  wire [2:0] my_adder_12_io_i_add_en; // @[FanNetwork.scala 1177:29]
  wire [2:0] my_adder_12_io_i_cmd; // @[FanNetwork.scala 1177:29]
  wire [1:0] my_adder_12_io_o_vn_valid; // @[FanNetwork.scala 1177:29]
  wire [63:0] my_adder_12_io_o_vn; // @[FanNetwork.scala 1177:29]
  wire [31:0] my_adder_12_io_o_adder_0; // @[FanNetwork.scala 1177:29]
  wire [31:0] my_adder_12_io_o_adder_1; // @[FanNetwork.scala 1177:29]
  wire  my_adder_13_clock; // @[FanNetwork.scala 1194:29]
  wire  my_adder_13_reset; // @[FanNetwork.scala 1194:29]
  wire  my_adder_13_io_i_valid; // @[FanNetwork.scala 1194:29]
  wire [31:0] my_adder_13_io_i_data_bus_0; // @[FanNetwork.scala 1194:29]
  wire [31:0] my_adder_13_io_i_data_bus_1; // @[FanNetwork.scala 1194:29]
  wire [2:0] my_adder_13_io_i_add_en; // @[FanNetwork.scala 1194:29]
  wire [2:0] my_adder_13_io_i_cmd; // @[FanNetwork.scala 1194:29]
  wire [1:0] my_adder_13_io_o_vn_valid; // @[FanNetwork.scala 1194:29]
  wire [63:0] my_adder_13_io_o_vn; // @[FanNetwork.scala 1194:29]
  wire [31:0] my_adder_13_io_o_adder_0; // @[FanNetwork.scala 1194:29]
  wire [31:0] my_adder_13_io_o_adder_1; // @[FanNetwork.scala 1194:29]
  wire  my_adder_14_clock; // @[FanNetwork.scala 1211:29]
  wire  my_adder_14_reset; // @[FanNetwork.scala 1211:29]
  wire  my_adder_14_io_i_valid; // @[FanNetwork.scala 1211:29]
  wire [31:0] my_adder_14_io_i_data_bus_0; // @[FanNetwork.scala 1211:29]
  wire [31:0] my_adder_14_io_i_data_bus_1; // @[FanNetwork.scala 1211:29]
  wire [2:0] my_adder_14_io_i_add_en; // @[FanNetwork.scala 1211:29]
  wire [2:0] my_adder_14_io_i_cmd; // @[FanNetwork.scala 1211:29]
  wire [1:0] my_adder_14_io_o_vn_valid; // @[FanNetwork.scala 1211:29]
  wire [63:0] my_adder_14_io_o_vn; // @[FanNetwork.scala 1211:29]
  wire [31:0] my_adder_14_io_o_adder_0; // @[FanNetwork.scala 1211:29]
  wire [31:0] my_adder_14_io_o_adder_1; // @[FanNetwork.scala 1211:29]
  wire  my_adder_15_clock; // @[FanNetwork.scala 1228:29]
  wire  my_adder_15_reset; // @[FanNetwork.scala 1228:29]
  wire  my_adder_15_io_i_valid; // @[FanNetwork.scala 1228:29]
  wire [63:0] my_adder_15_io_i_data_bus_0; // @[FanNetwork.scala 1228:29]
  wire [63:0] my_adder_15_io_i_data_bus_1; // @[FanNetwork.scala 1228:29]
  wire [63:0] my_adder_15_io_i_data_bus_2; // @[FanNetwork.scala 1228:29]
  wire [63:0] my_adder_15_io_i_data_bus_3; // @[FanNetwork.scala 1228:29]
  wire [63:0] my_adder_15_io_i_data_bus_4; // @[FanNetwork.scala 1228:29]
  wire [63:0] my_adder_15_io_i_data_bus_5; // @[FanNetwork.scala 1228:29]
  wire [63:0] my_adder_15_io_i_data_bus_6; // @[FanNetwork.scala 1228:29]
  wire [63:0] my_adder_15_io_i_data_bus_7; // @[FanNetwork.scala 1228:29]
  wire [2:0] my_adder_15_io_i_add_en; // @[FanNetwork.scala 1228:29]
  wire [4:0] my_adder_15_io_i_cmd; // @[FanNetwork.scala 1228:29]
  wire [3:0] my_adder_15_io_i_sel; // @[FanNetwork.scala 1228:29]
  wire [63:0] my_adder_15_io_o_vn; // @[FanNetwork.scala 1228:29]
  wire [1:0] my_adder_15_io_o_vn_valid; // @[FanNetwork.scala 1228:29]
  wire [31:0] my_adder_15_io_o_adder; // @[FanNetwork.scala 1228:29]
  wire  my_adder_16_clock; // @[FanNetwork.scala 1245:29]
  wire  my_adder_16_reset; // @[FanNetwork.scala 1245:29]
  wire  my_adder_16_io_i_valid; // @[FanNetwork.scala 1245:29]
  wire [31:0] my_adder_16_io_i_data_bus_0; // @[FanNetwork.scala 1245:29]
  wire [31:0] my_adder_16_io_i_data_bus_1; // @[FanNetwork.scala 1245:29]
  wire [2:0] my_adder_16_io_i_add_en; // @[FanNetwork.scala 1245:29]
  wire [2:0] my_adder_16_io_i_cmd; // @[FanNetwork.scala 1245:29]
  wire [1:0] my_adder_16_io_o_vn_valid; // @[FanNetwork.scala 1245:29]
  wire [63:0] my_adder_16_io_o_vn; // @[FanNetwork.scala 1245:29]
  wire [31:0] my_adder_16_io_o_adder_0; // @[FanNetwork.scala 1245:29]
  wire [31:0] my_adder_16_io_o_adder_1; // @[FanNetwork.scala 1245:29]
  wire  my_adder_17_clock; // @[FanNetwork.scala 1262:29]
  wire  my_adder_17_reset; // @[FanNetwork.scala 1262:29]
  wire  my_adder_17_io_i_valid; // @[FanNetwork.scala 1262:29]
  wire [31:0] my_adder_17_io_i_data_bus_0; // @[FanNetwork.scala 1262:29]
  wire [31:0] my_adder_17_io_i_data_bus_1; // @[FanNetwork.scala 1262:29]
  wire [2:0] my_adder_17_io_i_add_en; // @[FanNetwork.scala 1262:29]
  wire [2:0] my_adder_17_io_i_cmd; // @[FanNetwork.scala 1262:29]
  wire [1:0] my_adder_17_io_o_vn_valid; // @[FanNetwork.scala 1262:29]
  wire [63:0] my_adder_17_io_o_vn; // @[FanNetwork.scala 1262:29]
  wire [31:0] my_adder_17_io_o_adder_0; // @[FanNetwork.scala 1262:29]
  wire [31:0] my_adder_17_io_o_adder_1; // @[FanNetwork.scala 1262:29]
  wire  my_adder_18_clock; // @[FanNetwork.scala 1279:29]
  wire  my_adder_18_reset; // @[FanNetwork.scala 1279:29]
  wire  my_adder_18_io_i_valid; // @[FanNetwork.scala 1279:29]
  wire [31:0] my_adder_18_io_i_data_bus_0; // @[FanNetwork.scala 1279:29]
  wire [31:0] my_adder_18_io_i_data_bus_1; // @[FanNetwork.scala 1279:29]
  wire [2:0] my_adder_18_io_i_add_en; // @[FanNetwork.scala 1279:29]
  wire [2:0] my_adder_18_io_i_cmd; // @[FanNetwork.scala 1279:29]
  wire [1:0] my_adder_18_io_o_vn_valid; // @[FanNetwork.scala 1279:29]
  wire [63:0] my_adder_18_io_o_vn; // @[FanNetwork.scala 1279:29]
  wire [31:0] my_adder_18_io_o_adder_0; // @[FanNetwork.scala 1279:29]
  wire [31:0] my_adder_18_io_o_adder_1; // @[FanNetwork.scala 1279:29]
  wire  my_adder_19_clock; // @[FanNetwork.scala 1296:29]
  wire  my_adder_19_reset; // @[FanNetwork.scala 1296:29]
  wire  my_adder_19_io_i_valid; // @[FanNetwork.scala 1296:29]
  wire [31:0] my_adder_19_io_i_data_bus_0; // @[FanNetwork.scala 1296:29]
  wire [31:0] my_adder_19_io_i_data_bus_1; // @[FanNetwork.scala 1296:29]
  wire [31:0] my_adder_19_io_i_data_bus_2; // @[FanNetwork.scala 1296:29]
  wire [31:0] my_adder_19_io_i_data_bus_3; // @[FanNetwork.scala 1296:29]
  wire [2:0] my_adder_19_io_i_add_en; // @[FanNetwork.scala 1296:29]
  wire [2:0] my_adder_19_io_i_cmd; // @[FanNetwork.scala 1296:29]
  wire [1:0] my_adder_19_io_i_sel; // @[FanNetwork.scala 1296:29]
  wire [1:0] my_adder_19_io_o_vn_valid; // @[FanNetwork.scala 1296:29]
  wire [63:0] my_adder_19_io_o_vn; // @[FanNetwork.scala 1296:29]
  wire [31:0] my_adder_19_io_o_adder_0; // @[FanNetwork.scala 1296:29]
  wire [31:0] my_adder_19_io_o_adder_1; // @[FanNetwork.scala 1296:29]
  wire  my_adder_20_clock; // @[FanNetwork.scala 1314:29]
  wire  my_adder_20_reset; // @[FanNetwork.scala 1314:29]
  wire  my_adder_20_io_i_valid; // @[FanNetwork.scala 1314:29]
  wire [31:0] my_adder_20_io_i_data_bus_0; // @[FanNetwork.scala 1314:29]
  wire [31:0] my_adder_20_io_i_data_bus_1; // @[FanNetwork.scala 1314:29]
  wire [2:0] my_adder_20_io_i_add_en; // @[FanNetwork.scala 1314:29]
  wire [2:0] my_adder_20_io_i_cmd; // @[FanNetwork.scala 1314:29]
  wire [1:0] my_adder_20_io_o_vn_valid; // @[FanNetwork.scala 1314:29]
  wire [63:0] my_adder_20_io_o_vn; // @[FanNetwork.scala 1314:29]
  wire [31:0] my_adder_20_io_o_adder_0; // @[FanNetwork.scala 1314:29]
  wire [31:0] my_adder_20_io_o_adder_1; // @[FanNetwork.scala 1314:29]
  wire  my_adder_21_clock; // @[FanNetwork.scala 1333:29]
  wire  my_adder_21_reset; // @[FanNetwork.scala 1333:29]
  wire  my_adder_21_io_i_valid; // @[FanNetwork.scala 1333:29]
  wire [31:0] my_adder_21_io_i_data_bus_0; // @[FanNetwork.scala 1333:29]
  wire [31:0] my_adder_21_io_i_data_bus_1; // @[FanNetwork.scala 1333:29]
  wire [2:0] my_adder_21_io_i_add_en; // @[FanNetwork.scala 1333:29]
  wire [2:0] my_adder_21_io_i_cmd; // @[FanNetwork.scala 1333:29]
  wire [1:0] my_adder_21_io_o_vn_valid; // @[FanNetwork.scala 1333:29]
  wire [63:0] my_adder_21_io_o_vn; // @[FanNetwork.scala 1333:29]
  wire [31:0] my_adder_21_io_o_adder_0; // @[FanNetwork.scala 1333:29]
  wire [31:0] my_adder_21_io_o_adder_1; // @[FanNetwork.scala 1333:29]
  wire  my_adder_22_clock; // @[FanNetwork.scala 1351:29]
  wire  my_adder_22_reset; // @[FanNetwork.scala 1351:29]
  wire  my_adder_22_io_i_valid; // @[FanNetwork.scala 1351:29]
  wire [31:0] my_adder_22_io_i_data_bus_0; // @[FanNetwork.scala 1351:29]
  wire [31:0] my_adder_22_io_i_data_bus_1; // @[FanNetwork.scala 1351:29]
  wire [2:0] my_adder_22_io_i_add_en; // @[FanNetwork.scala 1351:29]
  wire [2:0] my_adder_22_io_i_cmd; // @[FanNetwork.scala 1351:29]
  wire [1:0] my_adder_22_io_o_vn_valid; // @[FanNetwork.scala 1351:29]
  wire [63:0] my_adder_22_io_o_vn; // @[FanNetwork.scala 1351:29]
  wire [31:0] my_adder_22_io_o_adder_0; // @[FanNetwork.scala 1351:29]
  wire [31:0] my_adder_22_io_o_adder_1; // @[FanNetwork.scala 1351:29]
  wire  my_adder_23_clock; // @[FanNetwork.scala 1368:29]
  wire  my_adder_23_reset; // @[FanNetwork.scala 1368:29]
  wire  my_adder_23_io_i_valid; // @[FanNetwork.scala 1368:29]
  wire [63:0] my_adder_23_io_i_data_bus_0; // @[FanNetwork.scala 1368:29]
  wire [63:0] my_adder_23_io_i_data_bus_1; // @[FanNetwork.scala 1368:29]
  wire [63:0] my_adder_23_io_i_data_bus_2; // @[FanNetwork.scala 1368:29]
  wire [63:0] my_adder_23_io_i_data_bus_3; // @[FanNetwork.scala 1368:29]
  wire [63:0] my_adder_23_io_i_data_bus_4; // @[FanNetwork.scala 1368:29]
  wire [63:0] my_adder_23_io_i_data_bus_5; // @[FanNetwork.scala 1368:29]
  wire [2:0] my_adder_23_io_i_add_en; // @[FanNetwork.scala 1368:29]
  wire [4:0] my_adder_23_io_i_cmd; // @[FanNetwork.scala 1368:29]
  wire [3:0] my_adder_23_io_i_sel; // @[FanNetwork.scala 1368:29]
  wire [63:0] my_adder_23_io_o_vn; // @[FanNetwork.scala 1368:29]
  wire [1:0] my_adder_23_io_o_vn_valid; // @[FanNetwork.scala 1368:29]
  wire [31:0] my_adder_23_io_o_adder; // @[FanNetwork.scala 1368:29]
  wire  my_adder_24_clock; // @[FanNetwork.scala 1383:29]
  wire  my_adder_24_reset; // @[FanNetwork.scala 1383:29]
  wire  my_adder_24_io_i_valid; // @[FanNetwork.scala 1383:29]
  wire [31:0] my_adder_24_io_i_data_bus_0; // @[FanNetwork.scala 1383:29]
  wire [31:0] my_adder_24_io_i_data_bus_1; // @[FanNetwork.scala 1383:29]
  wire [2:0] my_adder_24_io_i_add_en; // @[FanNetwork.scala 1383:29]
  wire [2:0] my_adder_24_io_i_cmd; // @[FanNetwork.scala 1383:29]
  wire [1:0] my_adder_24_io_o_vn_valid; // @[FanNetwork.scala 1383:29]
  wire [63:0] my_adder_24_io_o_vn; // @[FanNetwork.scala 1383:29]
  wire [31:0] my_adder_24_io_o_adder_0; // @[FanNetwork.scala 1383:29]
  wire [31:0] my_adder_24_io_o_adder_1; // @[FanNetwork.scala 1383:29]
  wire  my_adder_25_clock; // @[FanNetwork.scala 1401:29]
  wire  my_adder_25_reset; // @[FanNetwork.scala 1401:29]
  wire  my_adder_25_io_i_valid; // @[FanNetwork.scala 1401:29]
  wire [31:0] my_adder_25_io_i_data_bus_0; // @[FanNetwork.scala 1401:29]
  wire [31:0] my_adder_25_io_i_data_bus_1; // @[FanNetwork.scala 1401:29]
  wire [2:0] my_adder_25_io_i_add_en; // @[FanNetwork.scala 1401:29]
  wire [2:0] my_adder_25_io_i_cmd; // @[FanNetwork.scala 1401:29]
  wire [1:0] my_adder_25_io_o_vn_valid; // @[FanNetwork.scala 1401:29]
  wire [63:0] my_adder_25_io_o_vn; // @[FanNetwork.scala 1401:29]
  wire [31:0] my_adder_25_io_o_adder_0; // @[FanNetwork.scala 1401:29]
  wire [31:0] my_adder_25_io_o_adder_1; // @[FanNetwork.scala 1401:29]
  wire  my_adder_26_clock; // @[FanNetwork.scala 1420:29]
  wire  my_adder_26_reset; // @[FanNetwork.scala 1420:29]
  wire  my_adder_26_io_i_valid; // @[FanNetwork.scala 1420:29]
  wire [31:0] my_adder_26_io_i_data_bus_0; // @[FanNetwork.scala 1420:29]
  wire [31:0] my_adder_26_io_i_data_bus_1; // @[FanNetwork.scala 1420:29]
  wire [2:0] my_adder_26_io_i_add_en; // @[FanNetwork.scala 1420:29]
  wire [2:0] my_adder_26_io_i_cmd; // @[FanNetwork.scala 1420:29]
  wire [1:0] my_adder_26_io_o_vn_valid; // @[FanNetwork.scala 1420:29]
  wire [63:0] my_adder_26_io_o_vn; // @[FanNetwork.scala 1420:29]
  wire [31:0] my_adder_26_io_o_adder_0; // @[FanNetwork.scala 1420:29]
  wire [31:0] my_adder_26_io_o_adder_1; // @[FanNetwork.scala 1420:29]
  wire  my_adder_27_clock; // @[FanNetwork.scala 1437:29]
  wire  my_adder_27_reset; // @[FanNetwork.scala 1437:29]
  wire  my_adder_27_io_i_valid; // @[FanNetwork.scala 1437:29]
  wire [63:0] my_adder_27_io_i_data_bus_0; // @[FanNetwork.scala 1437:29]
  wire [63:0] my_adder_27_io_i_data_bus_1; // @[FanNetwork.scala 1437:29]
  wire [63:0] my_adder_27_io_i_data_bus_2; // @[FanNetwork.scala 1437:29]
  wire [63:0] my_adder_27_io_i_data_bus_3; // @[FanNetwork.scala 1437:29]
  wire [2:0] my_adder_27_io_i_add_en; // @[FanNetwork.scala 1437:29]
  wire [4:0] my_adder_27_io_i_cmd; // @[FanNetwork.scala 1437:29]
  wire [1:0] my_adder_27_io_i_sel; // @[FanNetwork.scala 1437:29]
  wire [63:0] my_adder_27_io_o_vn; // @[FanNetwork.scala 1437:29]
  wire [1:0] my_adder_27_io_o_vn_valid; // @[FanNetwork.scala 1437:29]
  wire [31:0] my_adder_27_io_o_adder; // @[FanNetwork.scala 1437:29]
  wire  my_adder_28_clock; // @[FanNetwork.scala 1456:29]
  wire  my_adder_28_reset; // @[FanNetwork.scala 1456:29]
  wire  my_adder_28_io_i_valid; // @[FanNetwork.scala 1456:29]
  wire [31:0] my_adder_28_io_i_data_bus_0; // @[FanNetwork.scala 1456:29]
  wire [31:0] my_adder_28_io_i_data_bus_1; // @[FanNetwork.scala 1456:29]
  wire [2:0] my_adder_28_io_i_add_en; // @[FanNetwork.scala 1456:29]
  wire [2:0] my_adder_28_io_i_cmd; // @[FanNetwork.scala 1456:29]
  wire [1:0] my_adder_28_io_o_vn_valid; // @[FanNetwork.scala 1456:29]
  wire [63:0] my_adder_28_io_o_vn; // @[FanNetwork.scala 1456:29]
  wire [31:0] my_adder_28_io_o_adder_0; // @[FanNetwork.scala 1456:29]
  wire [31:0] my_adder_28_io_o_adder_1; // @[FanNetwork.scala 1456:29]
  wire  my_adder_29_clock; // @[FanNetwork.scala 1474:29]
  wire  my_adder_29_reset; // @[FanNetwork.scala 1474:29]
  wire  my_adder_29_io_i_valid; // @[FanNetwork.scala 1474:29]
  wire [63:0] my_adder_29_io_i_data_bus_0; // @[FanNetwork.scala 1474:29]
  wire [63:0] my_adder_29_io_i_data_bus_1; // @[FanNetwork.scala 1474:29]
  wire [2:0] my_adder_29_io_i_add_en; // @[FanNetwork.scala 1474:29]
  wire [4:0] my_adder_29_io_i_cmd; // @[FanNetwork.scala 1474:29]
  wire [63:0] my_adder_29_io_o_vn; // @[FanNetwork.scala 1474:29]
  wire [1:0] my_adder_29_io_o_vn_valid; // @[FanNetwork.scala 1474:29]
  wire [31:0] my_adder_29_io_o_adder; // @[FanNetwork.scala 1474:29]
  wire  my_adder_30_clock; // @[FanNetwork.scala 1491:29]
  wire  my_adder_30_reset; // @[FanNetwork.scala 1491:29]
  wire  my_adder_30_io_i_valid; // @[FanNetwork.scala 1491:29]
  wire [63:0] my_adder_30_io_i_data_bus_0; // @[FanNetwork.scala 1491:29]
  wire [63:0] my_adder_30_io_i_data_bus_1; // @[FanNetwork.scala 1491:29]
  wire [2:0] my_adder_30_io_i_add_en; // @[FanNetwork.scala 1491:29]
  wire [4:0] my_adder_30_io_i_cmd; // @[FanNetwork.scala 1491:29]
  wire [63:0] my_adder_30_io_o_vn; // @[FanNetwork.scala 1491:29]
  wire [1:0] my_adder_30_io_o_vn_valid; // @[FanNetwork.scala 1491:29]
  wire [31:0] my_adder_30_io_o_adder; // @[FanNetwork.scala 1491:29]
  reg [31:0] r_fan_ff_lvl_0_to_4_0; // @[FanNetwork.scala 27:38]
  reg [31:0] r_fan_ff_lvl_0_to_4_1; // @[FanNetwork.scala 27:38]
  reg [31:0] r_fan_ff_lvl_0_to_3_0; // @[FanNetwork.scala 28:38]
  reg [31:0] r_fan_ff_lvl_0_to_3_1; // @[FanNetwork.scala 28:38]
  reg [31:0] r_fan_ff_lvl_0_to_3_2; // @[FanNetwork.scala 28:38]
  reg [31:0] r_fan_ff_lvl_0_to_3_3; // @[FanNetwork.scala 28:38]
  reg [31:0] r_fan_ff_lvl_0_to_3_4; // @[FanNetwork.scala 28:38]
  reg [31:0] r_fan_ff_lvl_0_to_3_5; // @[FanNetwork.scala 28:38]
  reg [31:0] r_fan_ff_lvl_0_to_2_0; // @[FanNetwork.scala 29:38]
  reg [31:0] r_fan_ff_lvl_0_to_2_1; // @[FanNetwork.scala 29:38]
  reg [31:0] r_fan_ff_lvl_0_to_2_2; // @[FanNetwork.scala 29:38]
  reg [31:0] r_fan_ff_lvl_0_to_2_3; // @[FanNetwork.scala 29:38]
  reg [31:0] r_fan_ff_lvl_0_to_2_4; // @[FanNetwork.scala 29:38]
  reg [31:0] r_fan_ff_lvl_0_to_2_5; // @[FanNetwork.scala 29:38]
  reg [31:0] r_fan_ff_lvl_0_to_2_6; // @[FanNetwork.scala 29:38]
  reg [31:0] r_fan_ff_lvl_0_to_2_7; // @[FanNetwork.scala 29:38]
  reg [31:0] r_fan_ff_lvl_0_to_2_8; // @[FanNetwork.scala 29:38]
  reg [31:0] r_fan_ff_lvl_0_to_2_9; // @[FanNetwork.scala 29:38]
  reg [31:0] r_fan_ff_lvl_0_to_2_10; // @[FanNetwork.scala 29:38]
  reg [31:0] r_fan_ff_lvl_0_to_2_11; // @[FanNetwork.scala 29:38]
  reg [31:0] r_fan_ff_lvl_0_to_2_12; // @[FanNetwork.scala 29:38]
  reg [31:0] r_fan_ff_lvl_0_to_2_13; // @[FanNetwork.scala 29:38]
  reg [31:0] r_fan_ff_lvl_1_to_4_0; // @[FanNetwork.scala 30:38]
  reg [31:0] r_fan_ff_lvl_1_to_4_1; // @[FanNetwork.scala 30:38]
  reg [31:0] r_fan_ff_lvl_1_to_3_0; // @[FanNetwork.scala 31:38]
  reg [31:0] r_fan_ff_lvl_1_to_3_1; // @[FanNetwork.scala 31:38]
  reg [31:0] r_fan_ff_lvl_1_to_3_2; // @[FanNetwork.scala 31:38]
  reg [31:0] r_fan_ff_lvl_1_to_3_3; // @[FanNetwork.scala 31:38]
  reg [31:0] r_fan_ff_lvl_1_to_3_4; // @[FanNetwork.scala 31:38]
  reg [31:0] r_fan_ff_lvl_1_to_3_5; // @[FanNetwork.scala 31:38]
  reg [31:0] r_fan_ff_lvl_2_to_4_0; // @[FanNetwork.scala 32:38]
  reg [31:0] r_fan_ff_lvl_2_to_4_1; // @[FanNetwork.scala 32:38]
  reg [31:0] r_lvl_output_ff_0; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_1; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_2; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_3; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_4; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_5; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_6; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_7; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_8; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_9; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_10; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_11; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_12; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_13; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_14; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_15; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_16; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_17; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_18; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_19; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_20; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_21; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_22; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_23; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_24; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_25; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_26; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_27; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_28; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_29; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_30; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_31; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_32; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_33; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_34; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_35; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_36; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_37; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_38; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_39; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_40; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_41; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_42; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_43; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_44; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_45; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_46; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_47; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_48; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_49; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_50; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_51; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_52; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_53; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_54; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_55; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_56; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_57; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_58; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_59; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_60; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_61; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_62; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_63; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_64; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_65; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_66; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_67; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_68; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_69; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_70; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_71; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_72; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_73; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_74; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_75; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_76; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_77; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_78; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_79; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_80; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_81; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_82; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_83; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_84; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_85; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_86; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_87; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_88; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_89; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_90; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_91; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_92; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_93; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_94; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_95; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_96; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_97; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_98; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_99; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_100; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_101; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_102; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_103; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_104; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_105; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_106; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_107; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_108; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_109; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_110; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_112; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_113; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_114; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_115; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_116; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_117; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_118; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_119; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_120; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_121; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_122; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_123; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_124; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_125; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_126; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_127; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_128; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_129; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_130; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_131; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_132; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_133; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_134; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_135; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_136; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_137; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_138; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_139; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_140; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_141; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_142; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_143; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_144; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_145; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_146; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_147; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_148; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_149; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_150; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_151; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_152; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_153; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_154; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_155; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_156; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_157; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_158; // @[FanNetwork.scala 45:34]
  reg [31:0] r_lvl_output_ff_159; // @[FanNetwork.scala 45:34]
  reg  r_lvl_output_ff_valid_0; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_1; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_2; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_3; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_4; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_5; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_6; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_7; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_8; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_9; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_10; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_11; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_12; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_13; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_14; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_15; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_16; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_17; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_18; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_19; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_20; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_21; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_22; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_23; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_24; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_25; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_26; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_27; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_28; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_29; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_30; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_31; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_32; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_33; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_34; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_35; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_36; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_37; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_38; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_39; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_40; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_41; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_42; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_43; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_44; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_45; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_46; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_47; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_48; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_49; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_50; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_51; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_52; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_53; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_54; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_55; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_56; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_57; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_58; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_59; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_60; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_61; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_62; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_63; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_64; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_65; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_66; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_67; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_68; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_69; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_70; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_71; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_72; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_73; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_74; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_75; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_76; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_77; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_78; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_79; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_80; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_81; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_82; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_83; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_84; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_85; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_86; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_87; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_88; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_89; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_90; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_91; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_92; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_93; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_94; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_95; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_96; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_97; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_98; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_99; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_100; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_101; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_102; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_103; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_104; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_105; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_106; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_107; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_108; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_109; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_110; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_111; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_112; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_113; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_114; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_115; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_116; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_117; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_118; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_119; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_120; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_121; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_122; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_123; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_124; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_125; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_126; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_127; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_128; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_129; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_130; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_131; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_132; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_133; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_134; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_135; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_136; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_137; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_138; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_139; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_140; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_141; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_142; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_143; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_144; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_145; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_146; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_147; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_148; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_149; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_150; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_151; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_152; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_153; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_154; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_155; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_156; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_157; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_158; // @[FanNetwork.scala 46:40]
  reg  r_lvl_output_ff_valid_159; // @[FanNetwork.scala 46:40]
  reg  r_valid_0; // @[FanNetwork.scala 47:26]
  reg  r_valid_1; // @[FanNetwork.scala 47:26]
  reg  r_valid_2; // @[FanNetwork.scala 47:26]
  reg  r_valid_3; // @[FanNetwork.scala 47:26]
  reg  r_valid_4; // @[FanNetwork.scala 47:26]
  reg [31:0] r_final_sum; // @[FanNetwork.scala 49:30]
  reg  r_final_add; // @[FanNetwork.scala 50:30]
  reg  r_final_add2; // @[FanNetwork.scala 51:31]
  wire  w_vn_lvl_0_valid_1 = my_adder_0_io_o_vn_valid[1]; // @[FanNetwork.scala 994:52]
  wire  w_vn_lvl_0_valid_0 = my_adder_0_io_o_vn_valid[0]; // @[FanNetwork.scala 993:52]
  wire  _T_9 = w_vn_lvl_0_valid_1 & ~w_vn_lvl_0_valid_0; // @[FanNetwork.scala 68:48]
  wire  _T_14 = ~w_vn_lvl_0_valid_1 & w_vn_lvl_0_valid_0; // @[FanNetwork.scala 73:48]
  wire [31:0] w_vn_lvl_0_0 = my_adder_0_io_o_vn[31:0]; // @[FanNetwork.scala 991:40]
  wire [31:0] w_vn_lvl_0_1 = my_adder_0_io_o_vn[63:32]; // @[FanNetwork.scala 992:40]
  wire  _GEN_6 = w_vn_lvl_0_valid_1 & ~w_vn_lvl_0_valid_0 ? 1'h0 : _T_14; // @[FanNetwork.scala 68:83 72:30]
  wire  _GEN_9 = w_vn_lvl_0_valid_1 & w_vn_lvl_0_valid_0 | _T_9; // @[FanNetwork.scala 63:77 66:30]
  wire  _GEN_10 = w_vn_lvl_0_valid_1 & w_vn_lvl_0_valid_0 | _GEN_6; // @[FanNetwork.scala 63:77 67:30]
  wire  w_vn_lvl_0_valid_3 = my_adder_2_io_o_vn_valid[1]; // @[FanNetwork.scala 1022:52]
  wire  w_vn_lvl_0_valid_2 = my_adder_2_io_o_vn_valid[0]; // @[FanNetwork.scala 1021:52]
  wire  _T_24 = w_vn_lvl_0_valid_3 & ~w_vn_lvl_0_valid_2; // @[FanNetwork.scala 90:48]
  wire  _T_29 = ~w_vn_lvl_0_valid_3 & w_vn_lvl_0_valid_2; // @[FanNetwork.scala 95:48]
  wire [31:0] w_vn_lvl_0_2 = my_adder_2_io_o_vn[31:0]; // @[FanNetwork.scala 1018:40]
  wire [31:0] w_vn_lvl_0_3 = my_adder_2_io_o_vn[63:32]; // @[FanNetwork.scala 1019:40]
  wire  _GEN_17 = w_vn_lvl_0_valid_3 & ~w_vn_lvl_0_valid_2 ? 1'h0 : _T_29; // @[FanNetwork.scala 90:83 94:34]
  wire  _GEN_20 = w_vn_lvl_0_valid_3 & w_vn_lvl_0_valid_2 | _T_24; // @[FanNetwork.scala 85:77 88:34]
  wire  _GEN_21 = w_vn_lvl_0_valid_3 & w_vn_lvl_0_valid_2 | _GEN_17; // @[FanNetwork.scala 85:77 89:34]
  wire  w_vn_lvl_0_valid_5 = my_adder_4_io_o_vn_valid[1]; // @[FanNetwork.scala 1054:52]
  wire  w_vn_lvl_0_valid_4 = my_adder_4_io_o_vn_valid[0]; // @[FanNetwork.scala 1053:52]
  wire  _T_39 = w_vn_lvl_0_valid_5 & ~w_vn_lvl_0_valid_4; // @[FanNetwork.scala 112:48]
  wire  _T_44 = ~w_vn_lvl_0_valid_5 & w_vn_lvl_0_valid_4; // @[FanNetwork.scala 117:48]
  wire [31:0] w_vn_lvl_0_4 = my_adder_4_io_o_vn[31:0]; // @[FanNetwork.scala 1050:40]
  wire [31:0] w_vn_lvl_0_5 = my_adder_4_io_o_vn[63:32]; // @[FanNetwork.scala 1051:40]
  wire  _GEN_28 = w_vn_lvl_0_valid_5 & ~w_vn_lvl_0_valid_4 ? 1'h0 : _T_44; // @[FanNetwork.scala 112:83 116:30]
  wire  _GEN_31 = w_vn_lvl_0_valid_5 & w_vn_lvl_0_valid_4 | _T_39; // @[FanNetwork.scala 107:77 110:30]
  wire  _GEN_32 = w_vn_lvl_0_valid_5 & w_vn_lvl_0_valid_4 | _GEN_28; // @[FanNetwork.scala 107:77 111:30]
  wire  w_vn_lvl_0_valid_7 = my_adder_6_io_o_vn_valid[1]; // @[FanNetwork.scala 1087:52]
  wire  w_vn_lvl_0_valid_6 = my_adder_6_io_o_vn_valid[0]; // @[FanNetwork.scala 1086:52]
  wire  _T_54 = w_vn_lvl_0_valid_7 & ~w_vn_lvl_0_valid_6; // @[FanNetwork.scala 135:48]
  wire  _T_59 = ~w_vn_lvl_0_valid_7 & w_vn_lvl_0_valid_6; // @[FanNetwork.scala 140:48]
  wire [31:0] w_vn_lvl_0_6 = my_adder_6_io_o_vn[31:0]; // @[FanNetwork.scala 1083:40]
  wire [31:0] w_vn_lvl_0_7 = my_adder_6_io_o_vn[63:32]; // @[FanNetwork.scala 1084:40]
  wire  _GEN_39 = w_vn_lvl_0_valid_7 & ~w_vn_lvl_0_valid_6 ? 1'h0 : _T_59; // @[FanNetwork.scala 135:83 139:30]
  wire  _GEN_42 = w_vn_lvl_0_valid_7 & w_vn_lvl_0_valid_6 | _T_54; // @[FanNetwork.scala 130:77 133:30]
  wire  _GEN_43 = w_vn_lvl_0_valid_7 & w_vn_lvl_0_valid_6 | _GEN_39; // @[FanNetwork.scala 130:77 134:30]
  wire  w_vn_lvl_0_valid_9 = my_adder_8_io_o_vn_valid[0]; // @[FanNetwork.scala 1120:52]
  wire  w_vn_lvl_0_valid_8 = my_adder_8_io_o_vn_valid[1]; // @[FanNetwork.scala 1119:52]
  wire  _T_66 = w_vn_lvl_0_valid_9 & ~w_vn_lvl_0_valid_8; // @[FanNetwork.scala 158:40]
  wire  _T_70 = ~w_vn_lvl_0_valid_9 & w_vn_lvl_0_valid_8; // @[FanNetwork.scala 163:41]
  wire [31:0] w_vn_lvl_0_8 = my_adder_8_io_o_vn[31:0]; // @[FanNetwork.scala 1116:40]
  wire [31:0] w_vn_lvl_0_9 = my_adder_8_io_o_vn[63:32]; // @[FanNetwork.scala 1117:40]
  wire  _GEN_50 = w_vn_lvl_0_valid_9 & ~w_vn_lvl_0_valid_8 ? 1'h0 : _T_70; // @[FanNetwork.scala 158:68 162:30]
  wire  _GEN_53 = w_vn_lvl_0_valid_9 & w_vn_lvl_0_valid_8 | _T_66; // @[FanNetwork.scala 153:61 156:30]
  wire  _GEN_54 = w_vn_lvl_0_valid_9 & w_vn_lvl_0_valid_8 | _GEN_50; // @[FanNetwork.scala 153:61 157:30]
  wire  w_vn_lvl_0_valid_11 = my_adder_10_io_o_vn_valid[1]; // @[FanNetwork.scala 1152:58]
  wire  w_vn_lvl_0_valid_10 = my_adder_10_io_o_vn_valid[0]; // @[FanNetwork.scala 1151:54]
  wire  _T_77 = w_vn_lvl_0_valid_11 & ~w_vn_lvl_0_valid_10; // @[FanNetwork.scala 181:41]
  wire  _T_81 = ~w_vn_lvl_0_valid_11 & w_vn_lvl_0_valid_10; // @[FanNetwork.scala 186:42]
  wire [31:0] w_vn_lvl_0_10 = my_adder_10_io_o_vn[31:0]; // @[FanNetwork.scala 1148:42]
  wire  _GEN_61 = w_vn_lvl_0_valid_11 & ~w_vn_lvl_0_valid_10 ? 1'h0 : _T_81; // @[FanNetwork.scala 181:70 185:31]
  wire  _GEN_64 = w_vn_lvl_0_valid_11 & w_vn_lvl_0_valid_10 | _T_77; // @[FanNetwork.scala 176:63 179:31]
  wire  _GEN_65 = w_vn_lvl_0_valid_11 & w_vn_lvl_0_valid_10 | _GEN_61; // @[FanNetwork.scala 176:63 180:31]
  wire  w_vn_lvl_0_valid_13 = my_adder_12_io_o_vn_valid[1]; // @[FanNetwork.scala 1188:58]
  wire  w_vn_lvl_0_valid_12 = my_adder_12_io_o_vn_valid[0]; // @[FanNetwork.scala 1187:54]
  wire  _T_88 = w_vn_lvl_0_valid_13 & ~w_vn_lvl_0_valid_12; // @[FanNetwork.scala 204:41]
  wire  _T_92 = ~w_vn_lvl_0_valid_13 & w_vn_lvl_0_valid_12; // @[FanNetwork.scala 209:42]
  wire [31:0] w_vn_lvl_0_12 = my_adder_12_io_o_vn[31:0]; // @[FanNetwork.scala 1184:42]
  wire [31:0] w_vn_lvl_0_13 = my_adder_12_io_o_vn[63:32]; // @[FanNetwork.scala 1185:46]
  wire  _GEN_72 = w_vn_lvl_0_valid_13 & ~w_vn_lvl_0_valid_12 ? 1'h0 : _T_92; // @[FanNetwork.scala 204:70 208:31]
  wire  _GEN_75 = w_vn_lvl_0_valid_13 & w_vn_lvl_0_valid_12 | _T_88; // @[FanNetwork.scala 199:63 202:31]
  wire  _GEN_76 = w_vn_lvl_0_valid_13 & w_vn_lvl_0_valid_12 | _GEN_72; // @[FanNetwork.scala 199:63 203:31]
  wire  w_vn_lvl_0_valid_15 = my_adder_14_io_o_vn_valid[1]; // @[FanNetwork.scala 1222:54]
  wire  w_vn_lvl_0_valid_14 = my_adder_14_io_o_vn_valid[0]; // @[FanNetwork.scala 1221:54]
  wire  _T_99 = w_vn_lvl_0_valid_15 & ~w_vn_lvl_0_valid_14; // @[FanNetwork.scala 227:41]
  wire  _T_103 = ~w_vn_lvl_0_valid_15 & w_vn_lvl_0_valid_14; // @[FanNetwork.scala 232:42]
  wire [31:0] w_vn_lvl_0_14 = my_adder_14_io_o_vn[31:0]; // @[FanNetwork.scala 1218:42]
  wire [31:0] w_vn_lvl_0_15 = my_adder_14_io_o_vn[63:32]; // @[FanNetwork.scala 1219:42]
  wire  _GEN_83 = w_vn_lvl_0_valid_15 & ~w_vn_lvl_0_valid_14 ? 1'h0 : _T_103; // @[FanNetwork.scala 227:70 231:31]
  wire  _GEN_86 = w_vn_lvl_0_valid_15 & w_vn_lvl_0_valid_14 | _T_99; // @[FanNetwork.scala 222:63 225:31]
  wire  _GEN_87 = w_vn_lvl_0_valid_15 & w_vn_lvl_0_valid_14 | _GEN_83; // @[FanNetwork.scala 222:63 226:31]
  wire  w_vn_lvl_0_valid_17 = my_adder_16_io_o_vn_valid[1]; // @[FanNetwork.scala 1256:54]
  wire  w_vn_lvl_0_valid_16 = my_adder_16_io_o_vn_valid[0]; // @[FanNetwork.scala 1255:54]
  wire  _T_110 = w_vn_lvl_0_valid_17 & ~w_vn_lvl_0_valid_16; // @[FanNetwork.scala 250:41]
  wire  _T_114 = ~w_vn_lvl_0_valid_17 & w_vn_lvl_0_valid_16; // @[FanNetwork.scala 255:42]
  wire [31:0] w_vn_lvl_0_16 = my_adder_16_io_o_vn[31:0]; // @[FanNetwork.scala 1252:42]
  wire [31:0] w_vn_lvl_0_17 = my_adder_16_io_o_vn[63:32]; // @[FanNetwork.scala 1253:42]
  wire  _GEN_94 = w_vn_lvl_0_valid_17 & ~w_vn_lvl_0_valid_16 ? 1'h0 : _T_114; // @[FanNetwork.scala 250:70 254:31]
  wire  _GEN_97 = w_vn_lvl_0_valid_17 & w_vn_lvl_0_valid_16 | _T_110; // @[FanNetwork.scala 245:63 248:31]
  wire  _GEN_98 = w_vn_lvl_0_valid_17 & w_vn_lvl_0_valid_16 | _GEN_94; // @[FanNetwork.scala 245:63 249:31]
  wire  w_vn_lvl_0_valid_19 = my_adder_18_io_o_vn_valid[1]; // @[FanNetwork.scala 1290:54]
  wire  w_vn_lvl_0_valid_18 = my_adder_18_io_o_vn_valid[0]; // @[FanNetwork.scala 1289:54]
  wire  _T_121 = w_vn_lvl_0_valid_19 & ~w_vn_lvl_0_valid_18; // @[FanNetwork.scala 273:41]
  wire  _T_125 = ~w_vn_lvl_0_valid_19 & w_vn_lvl_0_valid_18; // @[FanNetwork.scala 278:42]
  wire [31:0] w_vn_lvl_0_18 = my_adder_18_io_o_vn[31:0]; // @[FanNetwork.scala 1286:42]
  wire [31:0] w_vn_lvl_0_19 = my_adder_18_io_o_vn[63:32]; // @[FanNetwork.scala 1287:42]
  wire  _GEN_105 = w_vn_lvl_0_valid_19 & ~w_vn_lvl_0_valid_18 ? 1'h0 : _T_125; // @[FanNetwork.scala 273:70 277:31]
  wire  _GEN_108 = w_vn_lvl_0_valid_19 & w_vn_lvl_0_valid_18 | _T_121; // @[FanNetwork.scala 268:63 271:31]
  wire  _GEN_109 = w_vn_lvl_0_valid_19 & w_vn_lvl_0_valid_18 | _GEN_105; // @[FanNetwork.scala 268:63 272:31]
  wire  w_vn_lvl_0_valid_21 = my_adder_20_io_o_vn_valid[1]; // @[FanNetwork.scala 1325:54]
  wire  w_vn_lvl_0_valid_20 = my_adder_20_io_o_vn_valid[0]; // @[FanNetwork.scala 1324:54]
  wire  _T_132 = w_vn_lvl_0_valid_21 & ~w_vn_lvl_0_valid_20; // @[FanNetwork.scala 296:41]
  wire  _T_136 = ~w_vn_lvl_0_valid_21 & w_vn_lvl_0_valid_20; // @[FanNetwork.scala 301:42]
  wire [31:0] w_vn_lvl_0_20 = my_adder_20_io_o_vn[31:0]; // @[FanNetwork.scala 1321:42]
  wire [31:0] w_vn_lvl_0_21 = my_adder_20_io_o_vn[63:32]; // @[FanNetwork.scala 1322:42]
  wire  _GEN_116 = w_vn_lvl_0_valid_21 & ~w_vn_lvl_0_valid_20 ? 1'h0 : _T_136; // @[FanNetwork.scala 296:70 300:31]
  wire  _GEN_119 = w_vn_lvl_0_valid_21 & w_vn_lvl_0_valid_20 | _T_132; // @[FanNetwork.scala 291:63 294:31]
  wire  _GEN_120 = w_vn_lvl_0_valid_21 & w_vn_lvl_0_valid_20 | _GEN_116; // @[FanNetwork.scala 291:63 295:31]
  wire  w_vn_lvl_0_valid_23 = my_adder_22_io_o_vn_valid[1]; // @[FanNetwork.scala 1362:54]
  wire  w_vn_lvl_0_valid_22 = my_adder_22_io_o_vn_valid[0]; // @[FanNetwork.scala 1361:54]
  wire  _T_143 = w_vn_lvl_0_valid_23 & ~w_vn_lvl_0_valid_22; // @[FanNetwork.scala 319:41]
  wire  _T_147 = ~w_vn_lvl_0_valid_23 & w_vn_lvl_0_valid_22; // @[FanNetwork.scala 324:42]
  wire [31:0] w_vn_lvl_0_22 = my_adder_22_io_o_vn[31:0]; // @[FanNetwork.scala 1358:42]
  wire [31:0] w_vn_lvl_0_23 = my_adder_22_io_o_vn[63:32]; // @[FanNetwork.scala 1359:42]
  wire  _GEN_127 = w_vn_lvl_0_valid_23 & ~w_vn_lvl_0_valid_22 ? 1'h0 : _T_147; // @[FanNetwork.scala 319:70 323:31]
  wire  _GEN_130 = w_vn_lvl_0_valid_23 & w_vn_lvl_0_valid_22 | _T_143; // @[FanNetwork.scala 314:63 317:31]
  wire  _GEN_131 = w_vn_lvl_0_valid_23 & w_vn_lvl_0_valid_22 | _GEN_127; // @[FanNetwork.scala 314:63 318:31]
  wire  w_vn_lvl_0_valid_25 = my_adder_24_io_o_vn_valid[1]; // @[FanNetwork.scala 1394:54]
  wire  w_vn_lvl_0_valid_24 = my_adder_24_io_o_vn_valid[0]; // @[FanNetwork.scala 1393:54]
  wire  _T_154 = w_vn_lvl_0_valid_25 & ~w_vn_lvl_0_valid_24; // @[FanNetwork.scala 342:41]
  wire  _T_158 = ~w_vn_lvl_0_valid_25 & w_vn_lvl_0_valid_24; // @[FanNetwork.scala 347:42]
  wire [31:0] w_vn_lvl_0_24 = my_adder_24_io_o_vn[31:0]; // @[FanNetwork.scala 1390:42]
  wire [31:0] w_vn_lvl_0_25 = my_adder_24_io_o_vn[63:32]; // @[FanNetwork.scala 1391:42]
  wire  _GEN_138 = w_vn_lvl_0_valid_25 & ~w_vn_lvl_0_valid_24 ? 1'h0 : _T_158; // @[FanNetwork.scala 342:70 346:31]
  wire  _GEN_141 = w_vn_lvl_0_valid_25 & w_vn_lvl_0_valid_24 | _T_154; // @[FanNetwork.scala 337:63 340:31]
  wire  _GEN_142 = w_vn_lvl_0_valid_25 & w_vn_lvl_0_valid_24 | _GEN_138; // @[FanNetwork.scala 337:63 341:31]
  wire  w_vn_lvl_0_valid_27 = my_adder_26_io_o_vn_valid[1]; // @[FanNetwork.scala 1431:54]
  wire  w_vn_lvl_0_valid_26 = my_adder_26_io_o_vn_valid[0]; // @[FanNetwork.scala 1430:54]
  wire  _T_165 = w_vn_lvl_0_valid_27 & ~w_vn_lvl_0_valid_26; // @[FanNetwork.scala 365:41]
  wire  _T_169 = ~w_vn_lvl_0_valid_27 & w_vn_lvl_0_valid_26; // @[FanNetwork.scala 370:42]
  wire [31:0] w_vn_lvl_0_26 = my_adder_26_io_o_vn[31:0]; // @[FanNetwork.scala 1427:42]
  wire [31:0] w_vn_lvl_0_27 = my_adder_26_io_o_vn[63:32]; // @[FanNetwork.scala 1428:42]
  wire  _GEN_149 = w_vn_lvl_0_valid_27 & ~w_vn_lvl_0_valid_26 ? 1'h0 : _T_169; // @[FanNetwork.scala 365:70 369:31]
  wire  _GEN_152 = w_vn_lvl_0_valid_27 & w_vn_lvl_0_valid_26 | _T_165; // @[FanNetwork.scala 360:63 363:31]
  wire  _GEN_153 = w_vn_lvl_0_valid_27 & w_vn_lvl_0_valid_26 | _GEN_149; // @[FanNetwork.scala 360:63 364:31]
  wire  w_vn_lvl_0_valid_29 = my_adder_28_io_o_vn_valid[1]; // @[FanNetwork.scala 1467:54]
  wire  w_vn_lvl_0_valid_28 = my_adder_28_io_o_vn_valid[0]; // @[FanNetwork.scala 1466:54]
  wire  _T_176 = w_vn_lvl_0_valid_29 & ~w_vn_lvl_0_valid_28; // @[FanNetwork.scala 388:41]
  wire  _T_180 = ~w_vn_lvl_0_valid_29 & w_vn_lvl_0_valid_28; // @[FanNetwork.scala 393:42]
  wire [31:0] w_vn_lvl_0_28 = my_adder_28_io_o_vn[31:0]; // @[FanNetwork.scala 1463:42]
  wire [31:0] w_vn_lvl_0_29 = my_adder_28_io_o_vn[63:32]; // @[FanNetwork.scala 1464:46]
  wire  _GEN_160 = w_vn_lvl_0_valid_29 & ~w_vn_lvl_0_valid_28 ? 1'h0 : _T_180; // @[FanNetwork.scala 388:70 392:31]
  wire  _GEN_163 = w_vn_lvl_0_valid_29 & w_vn_lvl_0_valid_28 | _T_176; // @[FanNetwork.scala 383:63 386:31]
  wire  _GEN_164 = w_vn_lvl_0_valid_29 & w_vn_lvl_0_valid_28 | _GEN_160; // @[FanNetwork.scala 383:63 387:31]
  wire  w_vn_lvl_0_valid_31 = my_adder_30_io_o_vn_valid[1]; // @[FanNetwork.scala 1502:54]
  wire  w_vn_lvl_0_valid_30 = my_adder_30_io_o_vn_valid[0]; // @[FanNetwork.scala 1501:54]
  wire  _T_187 = w_vn_lvl_0_valid_31 & ~w_vn_lvl_0_valid_30; // @[FanNetwork.scala 411:40]
  wire  _T_191 = ~w_vn_lvl_0_valid_31 & w_vn_lvl_0_valid_30; // @[FanNetwork.scala 416:41]
  wire [31:0] w_vn_lvl_0_30 = my_adder_30_io_o_vn[31:0]; // @[FanNetwork.scala 1498:42]
  wire [31:0] w_vn_lvl_0_31 = my_adder_30_io_o_vn[63:32]; // @[FanNetwork.scala 1499:42]
  wire  _GEN_171 = w_vn_lvl_0_valid_31 & ~w_vn_lvl_0_valid_30 ? 1'h0 : _T_191; // @[FanNetwork.scala 411:69 415:31]
  wire  _GEN_174 = w_vn_lvl_0_valid_31 & w_vn_lvl_0_valid_30 | _T_187; // @[FanNetwork.scala 406:62 409:31]
  wire  _GEN_175 = w_vn_lvl_0_valid_31 & w_vn_lvl_0_valid_30 | _GEN_171; // @[FanNetwork.scala 406:62 410:31]
  wire  w_vn_lvl_1_valid_0 = my_adder_1_io_o_vn_valid[0]; // @[FanNetwork.scala 1006:52]
  wire [31:0] w_vn_lvl_1_0 = my_adder_1_io_o_vn[31:0]; // @[FanNetwork.scala 1004:40]
  wire  _GEN_177 = w_vn_lvl_1_valid_0 | r_lvl_output_ff_valid_1; // @[FanNetwork.scala 434:34 436:35 439:35]
  wire  w_vn_lvl_1_valid_1 = my_adder_1_io_o_vn_valid[1]; // @[FanNetwork.scala 1007:52]
  wire [31:0] w_vn_lvl_1_1 = my_adder_1_io_o_vn[63:32]; // @[FanNetwork.scala 1005:40]
  wire  _GEN_179 = w_vn_lvl_1_valid_1 | r_lvl_output_ff_valid_2; // @[FanNetwork.scala 442:34 444:35 447:35]
  wire  w_vn_lvl_1_valid_2 = my_adder_5_io_o_vn_valid[0]; // @[FanNetwork.scala 1070:52]
  wire [31:0] w_vn_lvl_1_2 = my_adder_5_io_o_vn[31:0]; // @[FanNetwork.scala 1067:40]
  wire  _GEN_181 = w_vn_lvl_1_valid_2 | r_lvl_output_ff_valid_5; // @[FanNetwork.scala 456:34 458:35 461:35]
  wire  w_vn_lvl_1_valid_3 = my_adder_5_io_o_vn_valid[1]; // @[FanNetwork.scala 1071:52]
  wire [31:0] w_vn_lvl_1_3 = my_adder_5_io_o_vn[63:32]; // @[FanNetwork.scala 1068:40]
  wire  _GEN_183 = w_vn_lvl_1_valid_3 | r_lvl_output_ff_valid_6; // @[FanNetwork.scala 464:34 466:35 469:35]
  wire  w_vn_lvl_1_valid_4 = my_adder_9_io_o_vn_valid[0]; // @[FanNetwork.scala 1135:52]
  wire [31:0] w_vn_lvl_1_4 = my_adder_9_io_o_vn[31:0]; // @[FanNetwork.scala 1132:40]
  wire  _GEN_185 = w_vn_lvl_1_valid_4 | r_lvl_output_ff_valid_9; // @[FanNetwork.scala 480:34 482:35 485:35]
  wire  w_vn_lvl_1_valid_5 = my_adder_9_io_o_vn_valid[1]; // @[FanNetwork.scala 1136:56]
  wire [31:0] w_vn_lvl_1_5 = my_adder_9_io_o_vn[63:32]; // @[FanNetwork.scala 1133:44]
  wire  _GEN_187 = w_vn_lvl_1_valid_5 | r_lvl_output_ff_valid_10; // @[FanNetwork.scala 487:34 489:35 492:35]
  wire  w_vn_lvl_1_valid_6 = my_adder_13_io_o_vn_valid[0]; // @[FanNetwork.scala 1204:53]
  wire [31:0] w_vn_lvl_1_6 = my_adder_13_io_o_vn[31:0]; // @[FanNetwork.scala 1201:41]
  wire  _GEN_189 = w_vn_lvl_1_valid_6 | r_lvl_output_ff_valid_13; // @[FanNetwork.scala 501:34 503:35 506:35]
  wire  w_vn_lvl_1_valid_7 = my_adder_13_io_o_vn_valid[1]; // @[FanNetwork.scala 1205:57]
  wire [31:0] w_vn_lvl_1_7 = my_adder_13_io_o_vn[63:32]; // @[FanNetwork.scala 1202:45]
  wire  _GEN_191 = w_vn_lvl_1_valid_7 | r_lvl_output_ff_valid_14; // @[FanNetwork.scala 509:34 511:35 514:35]
  wire  w_vn_lvl_1_valid_8 = my_adder_17_io_o_vn_valid[0]; // @[FanNetwork.scala 1272:53]
  wire [31:0] w_vn_lvl_1_8 = my_adder_17_io_o_vn[31:0]; // @[FanNetwork.scala 1269:41]
  wire  _GEN_193 = w_vn_lvl_1_valid_8 | r_lvl_output_ff_valid_17; // @[FanNetwork.scala 522:34 524:35 527:35]
  wire  w_vn_lvl_1_valid_9 = my_adder_17_io_o_vn_valid[1]; // @[FanNetwork.scala 1273:53]
  wire [31:0] w_vn_lvl_1_9 = my_adder_17_io_o_vn[63:32]; // @[FanNetwork.scala 1270:41]
  wire  _GEN_195 = w_vn_lvl_1_valid_9 | r_lvl_output_ff_valid_18; // @[FanNetwork.scala 530:34 532:35 535:35]
  wire  w_vn_lvl_1_valid_10 = my_adder_21_io_o_vn_valid[0]; // @[FanNetwork.scala 1344:54]
  wire [31:0] w_vn_lvl_1_10 = my_adder_21_io_o_vn[31:0]; // @[FanNetwork.scala 1341:42]
  wire  _GEN_197 = w_vn_lvl_1_valid_10 | r_lvl_output_ff_valid_21; // @[FanNetwork.scala 546:35 548:35 551:35]
  wire  w_vn_lvl_1_valid_11 = my_adder_21_io_o_vn_valid[1]; // @[FanNetwork.scala 1345:54]
  wire [31:0] w_vn_lvl_1_11 = my_adder_21_io_o_vn[63:32]; // @[FanNetwork.scala 1342:42]
  wire  _GEN_199 = w_vn_lvl_1_valid_11 | r_lvl_output_ff_valid_22; // @[FanNetwork.scala 554:35 556:35 559:35]
  wire  w_vn_lvl_1_valid_12 = my_adder_25_io_o_vn_valid[0]; // @[FanNetwork.scala 1411:54]
  wire [31:0] w_vn_lvl_1_12 = my_adder_25_io_o_vn[31:0];
  wire  _GEN_201 = w_vn_lvl_1_valid_12 | r_lvl_output_ff_valid_25; // @[FanNetwork.scala 568:35 570:35 573:35]
  wire  w_vn_lvl_1_valid_13 = my_adder_25_io_o_vn_valid[1]; // @[FanNetwork.scala 1412:54]
  wire [31:0] w_vn_lvl_1_13 = my_adder_25_io_o_vn[63:32]; // @[FanNetwork.scala 1409:42]
  wire  _GEN_203 = w_vn_lvl_1_valid_13 | r_lvl_output_ff_valid_26; // @[FanNetwork.scala 576:35 578:35 581:35]
  wire  w_vn_lvl_1_valid_14 = my_adder_29_io_o_vn_valid[0]; // @[FanNetwork.scala 1484:54]
  wire [31:0] w_vn_lvl_1_14 = my_adder_29_io_o_vn[31:0]; // @[FanNetwork.scala 1481:42]
  wire  _GEN_205 = w_vn_lvl_1_valid_14 | r_lvl_output_ff_valid_29; // @[FanNetwork.scala 590:43 592:35 595:31]
  wire  w_vn_lvl_1_valid_15 = my_adder_29_io_o_vn_valid[1]; // @[FanNetwork.scala 1485:54]
  wire [31:0] w_vn_lvl_1_15 = my_adder_29_io_o_vn[63:32]; // @[FanNetwork.scala 1482:42]
  wire  _GEN_207 = w_vn_lvl_1_valid_15 | r_lvl_output_ff_valid_30; // @[FanNetwork.scala 598:43 600:35 603:35]
  wire  w_vn_lvl_2_valid_0 = my_adder_3_io_o_vn_valid[0]; // @[FanNetwork.scala 1038:52]
  wire [31:0] w_vn_lvl_2_0 = my_adder_3_io_o_vn[31:0]; // @[FanNetwork.scala 1035:40]
  wire  _GEN_209 = w_vn_lvl_2_valid_0 | r_lvl_output_ff_valid_35; // @[FanNetwork.scala 619:43 621:35 624:39]
  wire  w_vn_lvl_2_valid_1 = my_adder_3_io_o_vn_valid[1]; // @[FanNetwork.scala 1039:52]
  wire [31:0] w_vn_lvl_2_1 = my_adder_3_io_o_vn[63:32]; // @[FanNetwork.scala 1036:40]
  wire  _GEN_211 = w_vn_lvl_2_valid_1 | r_lvl_output_ff_valid_36; // @[FanNetwork.scala 627:43 629:35 632:35]
  wire  w_vn_lvl_2_valid_2 = my_adder_11_io_o_vn_valid[0]; // @[FanNetwork.scala 1170:53]
  wire [31:0] w_vn_lvl_2_2 = my_adder_11_io_o_vn[31:0]; // @[FanNetwork.scala 1167:41]
  wire  _GEN_213 = w_vn_lvl_2_valid_2 | r_lvl_output_ff_valid_43; // @[FanNetwork.scala 653:43 655:35 658:35]
  wire  w_vn_lvl_2_valid_3 = my_adder_11_io_o_vn_valid[1]; // @[FanNetwork.scala 1171:57]
  wire [31:0] w_vn_lvl_2_3 = my_adder_11_io_o_vn[63:32]; // @[FanNetwork.scala 1168:45]
  wire  _GEN_215 = w_vn_lvl_2_valid_3 | r_lvl_output_ff_valid_44; // @[FanNetwork.scala 661:43 663:35 666:35]
  wire  w_vn_lvl_2_valid_4 = my_adder_19_io_o_vn_valid[0]; // @[FanNetwork.scala 1306:53]
  wire [31:0] w_vn_lvl_2_4 = my_adder_19_io_o_vn[31:0]; // @[FanNetwork.scala 1303:41]
  wire  _GEN_217 = w_vn_lvl_2_valid_4 | r_lvl_output_ff_valid_51; // @[FanNetwork.scala 687:43 689:35 692:35]
  wire  w_vn_lvl_2_valid_5 = my_adder_19_io_o_vn_valid[1]; // @[FanNetwork.scala 1307:53]
  wire [31:0] w_vn_lvl_2_5 = my_adder_19_io_o_vn[63:32]; // @[FanNetwork.scala 1304:41]
  wire  _GEN_219 = w_vn_lvl_2_valid_5 | r_lvl_output_ff_valid_52; // @[FanNetwork.scala 695:40 697:35 700:31]
  wire  w_vn_lvl_2_valid_6 = my_adder_27_io_o_vn_valid[0]; // @[FanNetwork.scala 1447:53]
  wire [31:0] w_vn_lvl_2_6 = my_adder_27_io_o_vn[31:0]; // @[FanNetwork.scala 1444:41]
  wire  _GEN_221 = w_vn_lvl_2_valid_6 | r_lvl_output_ff_valid_59; // @[FanNetwork.scala 721:40 723:35 726:35]
  wire  w_vn_lvl_2_valid_7 = my_adder_27_io_o_vn_valid[1]; // @[FanNetwork.scala 1448:53]
  wire [31:0] w_vn_lvl_2_7 = my_adder_27_io_o_vn[63:32]; // @[FanNetwork.scala 1445:41]
  wire  _GEN_223 = w_vn_lvl_2_valid_7 | r_lvl_output_ff_valid_60; // @[FanNetwork.scala 729:40 731:35 734:35]
  wire  w_vn_lvl_3_valid_0 = my_adder_7_io_o_vn_valid[0]; // @[FanNetwork.scala 1104:53]
  wire [31:0] w_vn_lvl_3_0 = my_adder_7_io_o_vn[31:0]; // @[FanNetwork.scala 1101:40]
  wire  _GEN_225 = w_vn_lvl_3_valid_0 | r_lvl_output_ff_valid_71; // @[FanNetwork.scala 769:40 771:34 774:34]
  wire  w_vn_lvl_3_valid_1 = my_adder_7_io_o_vn_valid[1]; // @[FanNetwork.scala 1105:53]
  wire [31:0] w_vn_lvl_3_1 = my_adder_7_io_o_vn[63:32]; // @[FanNetwork.scala 1102:40]
  wire  _GEN_227 = w_vn_lvl_3_valid_1 | r_lvl_output_ff_valid_72; // @[FanNetwork.scala 777:40 779:34 782:34]
  wire  w_vn_lvl_3_valid_2 = my_adder_23_io_o_vn_valid[0]; // @[FanNetwork.scala 1378:53]
  wire [31:0] w_vn_lvl_3_2 = my_adder_23_io_o_vn[31:0]; // @[FanNetwork.scala 1375:41]
  wire  _GEN_229 = w_vn_lvl_3_valid_2 | r_lvl_output_ff_valid_87; // @[FanNetwork.scala 827:40 829:36 832:36]
  wire  w_vn_lvl_3_valid_3 = my_adder_23_io_o_vn_valid[1]; // @[FanNetwork.scala 1379:53]
  wire [31:0] w_vn_lvl_3_3 = my_adder_23_io_o_vn[63:32]; // @[FanNetwork.scala 1376:41]
  wire  _GEN_231 = w_vn_lvl_3_valid_3 | r_lvl_output_ff_valid_88; // @[FanNetwork.scala 835:41 837:36 840:36]
  wire  w_vn_lvl_4_valid_0 = my_adder_15_io_o_vn_valid[0]; // @[FanNetwork.scala 1239:53]
  wire [31:0] w_vn_lvl_4_0 = my_adder_15_io_o_vn[31:0]; // @[FanNetwork.scala 1236:41]
  wire  _GEN_233 = w_vn_lvl_4_valid_0 | r_lvl_output_ff_valid_111; // @[FanNetwork.scala 910:40 912:36 915:36]
  wire  w_vn_lvl_4_valid_1 = my_adder_15_io_o_vn_valid[1]; // @[FanNetwork.scala 1240:53]
  wire [31:0] w_vn_lvl_4_1 = my_adder_15_io_o_vn[63:32]; // @[FanNetwork.scala 1237:41]
  wire  _GEN_235 = w_vn_lvl_4_valid_1 | r_lvl_output_ff_valid_112; // @[FanNetwork.scala 918:40 920:36 923:36]
  wire [3:0] _my_adder_3_io_i_sel_T = {io_i_sel_bus_1,io_i_sel_bus_0}; // @[Cat.scala 33:92]
  wire [7:0] _my_adder_7_io_i_sel_T = {io_i_sel_bus_11,io_i_sel_bus_10,io_i_sel_bus_9,io_i_sel_bus_8}; // @[Cat.scala 33:92]
  wire [3:0] _my_adder_11_io_i_sel_T = {io_i_sel_bus_3,io_i_sel_bus_2}; // @[Cat.scala 33:92]
  wire [7:0] _my_adder_15_io_i_sel_T = {io_i_sel_bus_19,io_i_sel_bus_18,io_i_sel_bus_17,io_i_sel_bus_16}; // @[Cat.scala 33:92]
  wire [3:0] _my_adder_19_io_i_sel_T = {io_i_sel_bus_5,io_i_sel_bus_4}; // @[Cat.scala 33:92]
  wire [7:0] _my_adder_23_io_i_sel_T = {io_i_sel_bus_15,io_i_sel_bus_14,io_i_sel_bus_13,io_i_sel_bus_12}; // @[Cat.scala 33:92]
  wire [3:0] _my_adder_27_io_i_sel_T = {io_i_sel_bus_7,io_i_sel_bus_6}; // @[Cat.scala 33:92]
  wire [959:0] w_fan_lvl_0_0 = {{928'd0}, my_adder_0_io_o_adder};
  wire [959:0] w_fan_lvl_0_1 = {{928'd0}, my_adder_2_io_o_adder_0};
  wire [959:0] w_fan_lvl_0_2 = {{928'd0}, my_adder_2_io_o_adder_1};
  wire [959:0] w_fan_lvl_0_3 = {{928'd0}, my_adder_4_io_o_adder_0};
  wire [959:0] w_fan_lvl_0_4 = {{928'd0}, my_adder_4_io_o_adder_1};
  wire [959:0] w_fan_lvl_0_5 = {{928'd0}, my_adder_6_io_o_adder_0};
  wire [959:0] w_fan_lvl_0_6 = {{928'd0}, my_adder_6_io_o_adder_1};
  wire [959:0] w_fan_lvl_0_7 = {{928'd0}, my_adder_8_io_o_adder_0};
  wire [959:0] w_fan_lvl_0_8 = {{928'd0}, my_adder_8_io_o_adder_1};
  wire [959:0] w_fan_lvl_0_9 = {{928'd0}, my_adder_10_io_o_adder_0};
  wire [959:0] w_fan_lvl_0_10 = {{928'd0}, my_adder_10_io_o_adder_1};
  wire [959:0] w_fan_lvl_0_11 = {{928'd0}, my_adder_12_io_o_adder_0};
  wire [959:0] w_fan_lvl_0_12 = {{928'd0}, my_adder_12_io_o_adder_1};
  wire [959:0] w_fan_lvl_0_13 = {{928'd0}, my_adder_14_io_o_adder_0};
  wire [959:0] w_fan_lvl_0_14 = {{928'd0}, my_adder_14_io_o_adder_1};
  wire [959:0] w_fan_lvl_0_15 = {{928'd0}, my_adder_16_io_o_adder_0};
  wire [959:0] w_fan_lvl_0_16 = {{928'd0}, my_adder_16_io_o_adder_1};
  wire [959:0] w_fan_lvl_0_17 = {{928'd0}, my_adder_18_io_o_adder_0};
  wire [959:0] w_fan_lvl_0_18 = {{928'd0}, my_adder_18_io_o_adder_1};
  wire [959:0] w_fan_lvl_0_19 = {{928'd0}, my_adder_20_io_o_adder_0};
  wire [959:0] w_fan_lvl_0_20 = {{928'd0}, my_adder_20_io_o_adder_1};
  wire [959:0] w_fan_lvl_0_21 = {{928'd0}, my_adder_22_io_o_adder_0};
  wire [959:0] w_fan_lvl_0_22 = {{928'd0}, my_adder_22_io_o_adder_1};
  wire [959:0] w_fan_lvl_0_23 = {{928'd0}, my_adder_24_io_o_adder_0};
  wire [959:0] w_fan_lvl_0_24 = {{928'd0}, my_adder_24_io_o_adder_1};
  wire [959:0] w_fan_lvl_0_25 = {{928'd0}, my_adder_26_io_o_adder_0};
  wire [959:0] w_fan_lvl_0_26 = {{928'd0}, my_adder_26_io_o_adder_1};
  wire [959:0] w_fan_lvl_0_27 = {{928'd0}, my_adder_28_io_o_adder_0};
  wire [959:0] w_fan_lvl_0_28 = {{928'd0}, my_adder_28_io_o_adder_1};
  wire [959:0] w_fan_lvl_0_29 = {{928'd0}, my_adder_30_io_o_adder};
  wire [479:0] w_fan_lvl_1_0 = {{448'd0}, my_adder_1_io_o_adder};
  wire [479:0] w_fan_lvl_1_1 = {{448'd0}, my_adder_5_io_o_adder_0};
  wire [479:0] w_fan_lvl_1_2 = {{448'd0}, my_adder_5_io_o_adder_1};
  wire [479:0] w_fan_lvl_1_3 = {{448'd0}, my_adder_9_io_o_adder_0};
  wire [479:0] w_fan_lvl_1_4 = {{448'd0}, my_adder_9_io_o_adder_1};
  wire [479:0] w_fan_lvl_1_5 = {{448'd0}, my_adder_13_io_o_adder_0};
  wire [479:0] w_fan_lvl_1_6 = {{448'd0}, my_adder_13_io_o_adder_1};
  wire [479:0] w_fan_lvl_1_7 = {{448'd0}, my_adder_17_io_o_adder_0};
  wire [479:0] w_fan_lvl_1_8 = {{448'd0}, my_adder_17_io_o_adder_1};
  wire [479:0] w_fan_lvl_1_9 = {{448'd0}, my_adder_21_io_o_adder_0};
  wire [479:0] w_fan_lvl_1_10 = {{448'd0}, my_adder_21_io_o_adder_1};
  wire [479:0] w_fan_lvl_1_11 = {{448'd0}, my_adder_25_io_o_adder_0};
  wire [479:0] w_fan_lvl_1_12 = {{448'd0}, my_adder_25_io_o_adder_1};
  wire [479:0] w_fan_lvl_1_13 = {{448'd0}, my_adder_29_io_o_adder};
  wire [191:0] w_fan_lvl_2_0 = {{160'd0}, my_adder_3_io_o_adder};
  wire [191:0] w_fan_lvl_2_1 = {{160'd0}, my_adder_11_io_o_adder_0};
  wire [191:0] w_fan_lvl_2_2 = {{160'd0}, my_adder_11_io_o_adder_1};
  wire [191:0] w_fan_lvl_2_3 = {{160'd0}, my_adder_19_io_o_adder_0};
  wire [191:0] w_fan_lvl_2_4 = {{160'd0}, my_adder_19_io_o_adder_1};
  wire [191:0] w_fan_lvl_2_5 = {{160'd0}, my_adder_27_io_o_adder};
  wire [63:0] w_fan_lvl_3_0 = {{32'd0}, my_adder_7_io_o_adder};
  wire [63:0] w_fan_lvl_3_1 = {{32'd0}, my_adder_23_io_o_adder};
  wire [31:0] w_fan_lvl_4_0 = my_adder_15_io_o_adder;
  wire [479:0] _WIRE_9_1 = {{448'd0}, r_fan_ff_lvl_0_to_2_1}; // @[FanNetwork.scala 1031:{42,42}]
  wire [479:0] _WIRE_9_2 = {{448'd0}, r_fan_ff_lvl_0_to_2_0}; // @[FanNetwork.scala 1031:{42,42}]
  wire [191:0] _WIRE_13_1 = {{160'd0}, r_fan_ff_lvl_1_to_3_1}; // @[FanNetwork.scala 1096:{40,40}]
  wire [191:0] _WIRE_13_2 = {{160'd0}, r_fan_ff_lvl_0_to_3_1}; // @[FanNetwork.scala 1096:{40,40}]
  wire [191:0] _WIRE_13_3 = {{160'd0}, r_fan_ff_lvl_0_to_3_0}; // @[FanNetwork.scala 1096:{40,40}]
  wire [191:0] _WIRE_13_4 = {{160'd0}, r_fan_ff_lvl_1_to_3_0}; // @[FanNetwork.scala 1096:{40,40}]
  wire [479:0] _WIRE_17_1 = {{448'd0}, r_fan_ff_lvl_0_to_2_5}; // @[FanNetwork.scala 1161:{41,41}]
  wire [479:0] _WIRE_17_2 = {{448'd0}, r_fan_ff_lvl_0_to_2_4}; // @[FanNetwork.scala 1161:{41,41}]
  wire [479:0] _WIRE_25_1 = {{448'd0}, r_fan_ff_lvl_0_to_2_9}; // @[FanNetwork.scala 1299:{42,42}]
  wire [479:0] _WIRE_25_2 = {{448'd0}, r_fan_ff_lvl_0_to_2_8}; // @[FanNetwork.scala 1299:{42,42}]
  wire [191:0] _WIRE_29_1 = {{160'd0}, r_fan_ff_lvl_1_to_3_5}; // @[FanNetwork.scala 1371:{41,41}]
  wire [191:0] _WIRE_29_2 = {{160'd0}, r_fan_ff_lvl_0_to_3_5}; // @[FanNetwork.scala 1371:{41,41}]
  wire [191:0] _WIRE_29_3 = {{160'd0}, r_fan_ff_lvl_0_to_3_4}; // @[FanNetwork.scala 1371:{41,41}]
  wire [191:0] _WIRE_29_4 = {{160'd0}, r_fan_ff_lvl_1_to_3_4}; // @[FanNetwork.scala 1371:{41,41}]
  wire [479:0] _WIRE_33_1 = {{448'd0}, r_fan_ff_lvl_0_to_2_13}; // @[FanNetwork.scala 1440:{41,41}]
  wire [479:0] _WIRE_33_2 = {{448'd0}, r_fan_ff_lvl_0_to_2_12}; // @[FanNetwork.scala 1440:{41,41}]
  wire [959:0] _GEN_239 = reset ? 960'h0 : w_fan_lvl_0_2; // @[FanNetwork.scala 29:{38,38} 53:25]
  wire [959:0] _GEN_240 = reset ? 960'h0 : w_fan_lvl_0_3; // @[FanNetwork.scala 29:{38,38} 53:25]
  wire [959:0] _GEN_241 = reset ? 960'h0 : w_fan_lvl_0_6; // @[FanNetwork.scala 29:{38,38} 53:25]
  wire [959:0] _GEN_242 = reset ? 960'h0 : w_fan_lvl_0_7; // @[FanNetwork.scala 29:{38,38} 53:25]
  wire [959:0] _GEN_243 = reset ? 960'h0 : w_fan_lvl_0_10; // @[FanNetwork.scala 29:{38,38} 53:25]
  wire [959:0] _GEN_244 = reset ? 960'h0 : w_fan_lvl_0_11; // @[FanNetwork.scala 29:{38,38} 53:25]
  wire [959:0] _GEN_245 = reset ? 960'h0 : w_fan_lvl_0_14; // @[FanNetwork.scala 29:{38,38} 53:25]
  wire [959:0] _GEN_246 = reset ? 960'h0 : w_fan_lvl_0_15; // @[FanNetwork.scala 29:{38,38} 53:25]
  wire [959:0] _GEN_247 = reset ? 960'h0 : w_fan_lvl_0_18; // @[FanNetwork.scala 29:{38,38} 53:25]
  wire [959:0] _GEN_248 = reset ? 960'h0 : w_fan_lvl_0_19; // @[FanNetwork.scala 29:{38,38} 53:25]
  wire [959:0] _GEN_249 = reset ? 960'h0 : w_fan_lvl_0_22; // @[FanNetwork.scala 29:{38,38} 53:25]
  wire [959:0] _GEN_250 = reset ? 960'h0 : w_fan_lvl_0_23; // @[FanNetwork.scala 29:{38,38} 53:25]
  wire [959:0] _GEN_251 = reset ? 960'h0 : w_fan_lvl_0_26; // @[FanNetwork.scala 29:{38,38} 53:25]
  wire [959:0] _GEN_252 = reset ? 960'h0 : w_fan_lvl_0_27; // @[FanNetwork.scala 29:{38,38} 53:25]
  wire [479:0] _GEN_253 = reset ? 480'h0 : w_fan_lvl_1_2; // @[FanNetwork.scala 31:{38,38} 57:25]
  wire [479:0] _GEN_254 = reset ? 480'h0 : w_fan_lvl_1_3; // @[FanNetwork.scala 31:{38,38} 57:25]
  wire [479:0] _GEN_255 = reset ? 480'h0 : w_fan_lvl_1_6; // @[FanNetwork.scala 31:{38,38} 57:25]
  wire [479:0] _GEN_256 = reset ? 480'h0 : w_fan_lvl_1_7; // @[FanNetwork.scala 31:{38,38} 57:25]
  wire [479:0] _GEN_257 = reset ? 480'h0 : w_fan_lvl_1_10; // @[FanNetwork.scala 31:{38,38} 57:25]
  wire [479:0] _GEN_258 = reset ? 480'h0 : w_fan_lvl_1_11; // @[FanNetwork.scala 31:{38,38} 57:25]
  wire [191:0] _GEN_259 = reset ? 192'h0 : w_fan_lvl_2_2; // @[FanNetwork.scala 32:{38,38} 58:25]
  wire [191:0] _GEN_260 = reset ? 192'h0 : w_fan_lvl_2_3; // @[FanNetwork.scala 32:{38,38} 58:25]
  EdgeAdderSwitch my_adder_0 ( // @[FanNetwork.scala 984:28]
    .clock(my_adder_0_clock),
    .reset(my_adder_0_reset),
    .io_i_valid(my_adder_0_io_i_valid),
    .io_i_data_bus_0(my_adder_0_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_0_io_i_data_bus_1),
    .io_i_add_en(my_adder_0_io_i_add_en),
    .io_i_cmd(my_adder_0_io_i_cmd),
    .io_o_vn(my_adder_0_io_o_vn),
    .io_o_vn_valid(my_adder_0_io_o_vn_valid),
    .io_o_adder(my_adder_0_io_o_adder)
  );
  EdgeAdderSwitch my_adder_1 ( // @[FanNetwork.scala 997:28]
    .clock(my_adder_1_clock),
    .reset(my_adder_1_reset),
    .io_i_valid(my_adder_1_io_i_valid),
    .io_i_data_bus_0(my_adder_1_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_1_io_i_data_bus_1),
    .io_i_add_en(my_adder_1_io_i_add_en),
    .io_i_cmd(my_adder_1_io_i_cmd),
    .io_o_vn(my_adder_1_io_o_vn),
    .io_o_vn_valid(my_adder_1_io_o_vn_valid),
    .io_o_adder(my_adder_1_io_o_adder)
  );
  AdderSwitch my_adder_2 ( // @[FanNetwork.scala 1010:28]
    .clock(my_adder_2_clock),
    .reset(my_adder_2_reset),
    .io_i_valid(my_adder_2_io_i_valid),
    .io_i_data_bus_0(my_adder_2_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_2_io_i_data_bus_1),
    .io_i_add_en(my_adder_2_io_i_add_en),
    .io_i_cmd(my_adder_2_io_i_cmd),
    .io_o_vn_valid(my_adder_2_io_o_vn_valid),
    .io_o_vn(my_adder_2_io_o_vn),
    .io_o_adder_0(my_adder_2_io_o_adder_0),
    .io_o_adder_1(my_adder_2_io_o_adder_1)
  );
  EdgeAdderSwitch_2 my_adder_3 ( // @[FanNetwork.scala 1028:28]
    .clock(my_adder_3_clock),
    .reset(my_adder_3_reset),
    .io_i_valid(my_adder_3_io_i_valid),
    .io_i_data_bus_0(my_adder_3_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_3_io_i_data_bus_1),
    .io_i_data_bus_2(my_adder_3_io_i_data_bus_2),
    .io_i_data_bus_3(my_adder_3_io_i_data_bus_3),
    .io_i_add_en(my_adder_3_io_i_add_en),
    .io_i_cmd(my_adder_3_io_i_cmd),
    .io_i_sel(my_adder_3_io_i_sel),
    .io_o_vn(my_adder_3_io_o_vn),
    .io_o_vn_valid(my_adder_3_io_o_vn_valid),
    .io_o_adder(my_adder_3_io_o_adder)
  );
  AdderSwitch my_adder_4 ( // @[FanNetwork.scala 1043:28]
    .clock(my_adder_4_clock),
    .reset(my_adder_4_reset),
    .io_i_valid(my_adder_4_io_i_valid),
    .io_i_data_bus_0(my_adder_4_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_4_io_i_data_bus_1),
    .io_i_add_en(my_adder_4_io_i_add_en),
    .io_i_cmd(my_adder_4_io_i_cmd),
    .io_o_vn_valid(my_adder_4_io_o_vn_valid),
    .io_o_vn(my_adder_4_io_o_vn),
    .io_o_adder_0(my_adder_4_io_o_adder_0),
    .io_o_adder_1(my_adder_4_io_o_adder_1)
  );
  AdderSwitch my_adder_5 ( // @[FanNetwork.scala 1060:28]
    .clock(my_adder_5_clock),
    .reset(my_adder_5_reset),
    .io_i_valid(my_adder_5_io_i_valid),
    .io_i_data_bus_0(my_adder_5_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_5_io_i_data_bus_1),
    .io_i_add_en(my_adder_5_io_i_add_en),
    .io_i_cmd(my_adder_5_io_i_cmd),
    .io_o_vn_valid(my_adder_5_io_o_vn_valid),
    .io_o_vn(my_adder_5_io_o_vn),
    .io_o_adder_0(my_adder_5_io_o_adder_0),
    .io_o_adder_1(my_adder_5_io_o_adder_1)
  );
  AdderSwitch my_adder_6 ( // @[FanNetwork.scala 1076:28]
    .clock(my_adder_6_clock),
    .reset(my_adder_6_reset),
    .io_i_valid(my_adder_6_io_i_valid),
    .io_i_data_bus_0(my_adder_6_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_6_io_i_data_bus_1),
    .io_i_add_en(my_adder_6_io_i_add_en),
    .io_i_cmd(my_adder_6_io_i_cmd),
    .io_o_vn_valid(my_adder_6_io_o_vn_valid),
    .io_o_vn(my_adder_6_io_o_vn),
    .io_o_adder_0(my_adder_6_io_o_adder_0),
    .io_o_adder_1(my_adder_6_io_o_adder_1)
  );
  EdgeAdderSwitch_3 my_adder_7 ( // @[FanNetwork.scala 1092:28]
    .clock(my_adder_7_clock),
    .reset(my_adder_7_reset),
    .io_i_valid(my_adder_7_io_i_valid),
    .io_i_data_bus_0(my_adder_7_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_7_io_i_data_bus_1),
    .io_i_data_bus_2(my_adder_7_io_i_data_bus_2),
    .io_i_data_bus_3(my_adder_7_io_i_data_bus_3),
    .io_i_data_bus_4(my_adder_7_io_i_data_bus_4),
    .io_i_data_bus_5(my_adder_7_io_i_data_bus_5),
    .io_i_add_en(my_adder_7_io_i_add_en),
    .io_i_cmd(my_adder_7_io_i_cmd),
    .io_i_sel(my_adder_7_io_i_sel),
    .io_o_vn(my_adder_7_io_o_vn),
    .io_o_vn_valid(my_adder_7_io_o_vn_valid),
    .io_o_adder(my_adder_7_io_o_adder)
  );
  AdderSwitch my_adder_8 ( // @[FanNetwork.scala 1109:28]
    .clock(my_adder_8_clock),
    .reset(my_adder_8_reset),
    .io_i_valid(my_adder_8_io_i_valid),
    .io_i_data_bus_0(my_adder_8_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_8_io_i_data_bus_1),
    .io_i_add_en(my_adder_8_io_i_add_en),
    .io_i_cmd(my_adder_8_io_i_cmd),
    .io_o_vn_valid(my_adder_8_io_o_vn_valid),
    .io_o_vn(my_adder_8_io_o_vn),
    .io_o_adder_0(my_adder_8_io_o_adder_0),
    .io_o_adder_1(my_adder_8_io_o_adder_1)
  );
  AdderSwitch my_adder_9 ( // @[FanNetwork.scala 1125:28]
    .clock(my_adder_9_clock),
    .reset(my_adder_9_reset),
    .io_i_valid(my_adder_9_io_i_valid),
    .io_i_data_bus_0(my_adder_9_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_9_io_i_data_bus_1),
    .io_i_add_en(my_adder_9_io_i_add_en),
    .io_i_cmd(my_adder_9_io_i_cmd),
    .io_o_vn_valid(my_adder_9_io_o_vn_valid),
    .io_o_vn(my_adder_9_io_o_vn),
    .io_o_adder_0(my_adder_9_io_o_adder_0),
    .io_o_adder_1(my_adder_9_io_o_adder_1)
  );
  AdderSwitch my_adder_10 ( // @[FanNetwork.scala 1141:29]
    .clock(my_adder_10_clock),
    .reset(my_adder_10_reset),
    .io_i_valid(my_adder_10_io_i_valid),
    .io_i_data_bus_0(my_adder_10_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_10_io_i_data_bus_1),
    .io_i_add_en(my_adder_10_io_i_add_en),
    .io_i_cmd(my_adder_10_io_i_cmd),
    .io_o_vn_valid(my_adder_10_io_o_vn_valid),
    .io_o_vn(my_adder_10_io_o_vn),
    .io_o_adder_0(my_adder_10_io_o_adder_0),
    .io_o_adder_1(my_adder_10_io_o_adder_1)
  );
  AdderSwitch_7 my_adder_11 ( // @[FanNetwork.scala 1158:29]
    .clock(my_adder_11_clock),
    .reset(my_adder_11_reset),
    .io_i_valid(my_adder_11_io_i_valid),
    .io_i_data_bus_0(my_adder_11_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_11_io_i_data_bus_1),
    .io_i_data_bus_2(my_adder_11_io_i_data_bus_2),
    .io_i_data_bus_3(my_adder_11_io_i_data_bus_3),
    .io_i_add_en(my_adder_11_io_i_add_en),
    .io_i_cmd(my_adder_11_io_i_cmd),
    .io_i_sel(my_adder_11_io_i_sel),
    .io_o_vn_valid(my_adder_11_io_o_vn_valid),
    .io_o_vn(my_adder_11_io_o_vn),
    .io_o_adder_0(my_adder_11_io_o_adder_0),
    .io_o_adder_1(my_adder_11_io_o_adder_1)
  );
  AdderSwitch my_adder_12 ( // @[FanNetwork.scala 1177:29]
    .clock(my_adder_12_clock),
    .reset(my_adder_12_reset),
    .io_i_valid(my_adder_12_io_i_valid),
    .io_i_data_bus_0(my_adder_12_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_12_io_i_data_bus_1),
    .io_i_add_en(my_adder_12_io_i_add_en),
    .io_i_cmd(my_adder_12_io_i_cmd),
    .io_o_vn_valid(my_adder_12_io_o_vn_valid),
    .io_o_vn(my_adder_12_io_o_vn),
    .io_o_adder_0(my_adder_12_io_o_adder_0),
    .io_o_adder_1(my_adder_12_io_o_adder_1)
  );
  AdderSwitch my_adder_13 ( // @[FanNetwork.scala 1194:29]
    .clock(my_adder_13_clock),
    .reset(my_adder_13_reset),
    .io_i_valid(my_adder_13_io_i_valid),
    .io_i_data_bus_0(my_adder_13_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_13_io_i_data_bus_1),
    .io_i_add_en(my_adder_13_io_i_add_en),
    .io_i_cmd(my_adder_13_io_i_cmd),
    .io_o_vn_valid(my_adder_13_io_o_vn_valid),
    .io_o_vn(my_adder_13_io_o_vn),
    .io_o_adder_0(my_adder_13_io_o_adder_0),
    .io_o_adder_1(my_adder_13_io_o_adder_1)
  );
  AdderSwitch my_adder_14 ( // @[FanNetwork.scala 1211:29]
    .clock(my_adder_14_clock),
    .reset(my_adder_14_reset),
    .io_i_valid(my_adder_14_io_i_valid),
    .io_i_data_bus_0(my_adder_14_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_14_io_i_data_bus_1),
    .io_i_add_en(my_adder_14_io_i_add_en),
    .io_i_cmd(my_adder_14_io_i_cmd),
    .io_o_vn_valid(my_adder_14_io_o_vn_valid),
    .io_o_vn(my_adder_14_io_o_vn),
    .io_o_adder_0(my_adder_14_io_o_adder_0),
    .io_o_adder_1(my_adder_14_io_o_adder_1)
  );
  EdgeAdderSwitch_4 my_adder_15 ( // @[FanNetwork.scala 1228:29]
    .clock(my_adder_15_clock),
    .reset(my_adder_15_reset),
    .io_i_valid(my_adder_15_io_i_valid),
    .io_i_data_bus_0(my_adder_15_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_15_io_i_data_bus_1),
    .io_i_data_bus_2(my_adder_15_io_i_data_bus_2),
    .io_i_data_bus_3(my_adder_15_io_i_data_bus_3),
    .io_i_data_bus_4(my_adder_15_io_i_data_bus_4),
    .io_i_data_bus_5(my_adder_15_io_i_data_bus_5),
    .io_i_data_bus_6(my_adder_15_io_i_data_bus_6),
    .io_i_data_bus_7(my_adder_15_io_i_data_bus_7),
    .io_i_add_en(my_adder_15_io_i_add_en),
    .io_i_cmd(my_adder_15_io_i_cmd),
    .io_i_sel(my_adder_15_io_i_sel),
    .io_o_vn(my_adder_15_io_o_vn),
    .io_o_vn_valid(my_adder_15_io_o_vn_valid),
    .io_o_adder(my_adder_15_io_o_adder)
  );
  AdderSwitch my_adder_16 ( // @[FanNetwork.scala 1245:29]
    .clock(my_adder_16_clock),
    .reset(my_adder_16_reset),
    .io_i_valid(my_adder_16_io_i_valid),
    .io_i_data_bus_0(my_adder_16_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_16_io_i_data_bus_1),
    .io_i_add_en(my_adder_16_io_i_add_en),
    .io_i_cmd(my_adder_16_io_i_cmd),
    .io_o_vn_valid(my_adder_16_io_o_vn_valid),
    .io_o_vn(my_adder_16_io_o_vn),
    .io_o_adder_0(my_adder_16_io_o_adder_0),
    .io_o_adder_1(my_adder_16_io_o_adder_1)
  );
  AdderSwitch my_adder_17 ( // @[FanNetwork.scala 1262:29]
    .clock(my_adder_17_clock),
    .reset(my_adder_17_reset),
    .io_i_valid(my_adder_17_io_i_valid),
    .io_i_data_bus_0(my_adder_17_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_17_io_i_data_bus_1),
    .io_i_add_en(my_adder_17_io_i_add_en),
    .io_i_cmd(my_adder_17_io_i_cmd),
    .io_o_vn_valid(my_adder_17_io_o_vn_valid),
    .io_o_vn(my_adder_17_io_o_vn),
    .io_o_adder_0(my_adder_17_io_o_adder_0),
    .io_o_adder_1(my_adder_17_io_o_adder_1)
  );
  AdderSwitch my_adder_18 ( // @[FanNetwork.scala 1279:29]
    .clock(my_adder_18_clock),
    .reset(my_adder_18_reset),
    .io_i_valid(my_adder_18_io_i_valid),
    .io_i_data_bus_0(my_adder_18_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_18_io_i_data_bus_1),
    .io_i_add_en(my_adder_18_io_i_add_en),
    .io_i_cmd(my_adder_18_io_i_cmd),
    .io_o_vn_valid(my_adder_18_io_o_vn_valid),
    .io_o_vn(my_adder_18_io_o_vn),
    .io_o_adder_0(my_adder_18_io_o_adder_0),
    .io_o_adder_1(my_adder_18_io_o_adder_1)
  );
  AdderSwitch_7 my_adder_19 ( // @[FanNetwork.scala 1296:29]
    .clock(my_adder_19_clock),
    .reset(my_adder_19_reset),
    .io_i_valid(my_adder_19_io_i_valid),
    .io_i_data_bus_0(my_adder_19_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_19_io_i_data_bus_1),
    .io_i_data_bus_2(my_adder_19_io_i_data_bus_2),
    .io_i_data_bus_3(my_adder_19_io_i_data_bus_3),
    .io_i_add_en(my_adder_19_io_i_add_en),
    .io_i_cmd(my_adder_19_io_i_cmd),
    .io_i_sel(my_adder_19_io_i_sel),
    .io_o_vn_valid(my_adder_19_io_o_vn_valid),
    .io_o_vn(my_adder_19_io_o_vn),
    .io_o_adder_0(my_adder_19_io_o_adder_0),
    .io_o_adder_1(my_adder_19_io_o_adder_1)
  );
  AdderSwitch my_adder_20 ( // @[FanNetwork.scala 1314:29]
    .clock(my_adder_20_clock),
    .reset(my_adder_20_reset),
    .io_i_valid(my_adder_20_io_i_valid),
    .io_i_data_bus_0(my_adder_20_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_20_io_i_data_bus_1),
    .io_i_add_en(my_adder_20_io_i_add_en),
    .io_i_cmd(my_adder_20_io_i_cmd),
    .io_o_vn_valid(my_adder_20_io_o_vn_valid),
    .io_o_vn(my_adder_20_io_o_vn),
    .io_o_adder_0(my_adder_20_io_o_adder_0),
    .io_o_adder_1(my_adder_20_io_o_adder_1)
  );
  AdderSwitch my_adder_21 ( // @[FanNetwork.scala 1333:29]
    .clock(my_adder_21_clock),
    .reset(my_adder_21_reset),
    .io_i_valid(my_adder_21_io_i_valid),
    .io_i_data_bus_0(my_adder_21_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_21_io_i_data_bus_1),
    .io_i_add_en(my_adder_21_io_i_add_en),
    .io_i_cmd(my_adder_21_io_i_cmd),
    .io_o_vn_valid(my_adder_21_io_o_vn_valid),
    .io_o_vn(my_adder_21_io_o_vn),
    .io_o_adder_0(my_adder_21_io_o_adder_0),
    .io_o_adder_1(my_adder_21_io_o_adder_1)
  );
  AdderSwitch my_adder_22 ( // @[FanNetwork.scala 1351:29]
    .clock(my_adder_22_clock),
    .reset(my_adder_22_reset),
    .io_i_valid(my_adder_22_io_i_valid),
    .io_i_data_bus_0(my_adder_22_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_22_io_i_data_bus_1),
    .io_i_add_en(my_adder_22_io_i_add_en),
    .io_i_cmd(my_adder_22_io_i_cmd),
    .io_o_vn_valid(my_adder_22_io_o_vn_valid),
    .io_o_vn(my_adder_22_io_o_vn),
    .io_o_adder_0(my_adder_22_io_o_adder_0),
    .io_o_adder_1(my_adder_22_io_o_adder_1)
  );
  EdgeAdderSwitch_3 my_adder_23 ( // @[FanNetwork.scala 1368:29]
    .clock(my_adder_23_clock),
    .reset(my_adder_23_reset),
    .io_i_valid(my_adder_23_io_i_valid),
    .io_i_data_bus_0(my_adder_23_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_23_io_i_data_bus_1),
    .io_i_data_bus_2(my_adder_23_io_i_data_bus_2),
    .io_i_data_bus_3(my_adder_23_io_i_data_bus_3),
    .io_i_data_bus_4(my_adder_23_io_i_data_bus_4),
    .io_i_data_bus_5(my_adder_23_io_i_data_bus_5),
    .io_i_add_en(my_adder_23_io_i_add_en),
    .io_i_cmd(my_adder_23_io_i_cmd),
    .io_i_sel(my_adder_23_io_i_sel),
    .io_o_vn(my_adder_23_io_o_vn),
    .io_o_vn_valid(my_adder_23_io_o_vn_valid),
    .io_o_adder(my_adder_23_io_o_adder)
  );
  AdderSwitch my_adder_24 ( // @[FanNetwork.scala 1383:29]
    .clock(my_adder_24_clock),
    .reset(my_adder_24_reset),
    .io_i_valid(my_adder_24_io_i_valid),
    .io_i_data_bus_0(my_adder_24_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_24_io_i_data_bus_1),
    .io_i_add_en(my_adder_24_io_i_add_en),
    .io_i_cmd(my_adder_24_io_i_cmd),
    .io_o_vn_valid(my_adder_24_io_o_vn_valid),
    .io_o_vn(my_adder_24_io_o_vn),
    .io_o_adder_0(my_adder_24_io_o_adder_0),
    .io_o_adder_1(my_adder_24_io_o_adder_1)
  );
  AdderSwitch my_adder_25 ( // @[FanNetwork.scala 1401:29]
    .clock(my_adder_25_clock),
    .reset(my_adder_25_reset),
    .io_i_valid(my_adder_25_io_i_valid),
    .io_i_data_bus_0(my_adder_25_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_25_io_i_data_bus_1),
    .io_i_add_en(my_adder_25_io_i_add_en),
    .io_i_cmd(my_adder_25_io_i_cmd),
    .io_o_vn_valid(my_adder_25_io_o_vn_valid),
    .io_o_vn(my_adder_25_io_o_vn),
    .io_o_adder_0(my_adder_25_io_o_adder_0),
    .io_o_adder_1(my_adder_25_io_o_adder_1)
  );
  AdderSwitch my_adder_26 ( // @[FanNetwork.scala 1420:29]
    .clock(my_adder_26_clock),
    .reset(my_adder_26_reset),
    .io_i_valid(my_adder_26_io_i_valid),
    .io_i_data_bus_0(my_adder_26_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_26_io_i_data_bus_1),
    .io_i_add_en(my_adder_26_io_i_add_en),
    .io_i_cmd(my_adder_26_io_i_cmd),
    .io_o_vn_valid(my_adder_26_io_o_vn_valid),
    .io_o_vn(my_adder_26_io_o_vn),
    .io_o_adder_0(my_adder_26_io_o_adder_0),
    .io_o_adder_1(my_adder_26_io_o_adder_1)
  );
  EdgeAdderSwitch_2 my_adder_27 ( // @[FanNetwork.scala 1437:29]
    .clock(my_adder_27_clock),
    .reset(my_adder_27_reset),
    .io_i_valid(my_adder_27_io_i_valid),
    .io_i_data_bus_0(my_adder_27_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_27_io_i_data_bus_1),
    .io_i_data_bus_2(my_adder_27_io_i_data_bus_2),
    .io_i_data_bus_3(my_adder_27_io_i_data_bus_3),
    .io_i_add_en(my_adder_27_io_i_add_en),
    .io_i_cmd(my_adder_27_io_i_cmd),
    .io_i_sel(my_adder_27_io_i_sel),
    .io_o_vn(my_adder_27_io_o_vn),
    .io_o_vn_valid(my_adder_27_io_o_vn_valid),
    .io_o_adder(my_adder_27_io_o_adder)
  );
  AdderSwitch my_adder_28 ( // @[FanNetwork.scala 1456:29]
    .clock(my_adder_28_clock),
    .reset(my_adder_28_reset),
    .io_i_valid(my_adder_28_io_i_valid),
    .io_i_data_bus_0(my_adder_28_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_28_io_i_data_bus_1),
    .io_i_add_en(my_adder_28_io_i_add_en),
    .io_i_cmd(my_adder_28_io_i_cmd),
    .io_o_vn_valid(my_adder_28_io_o_vn_valid),
    .io_o_vn(my_adder_28_io_o_vn),
    .io_o_adder_0(my_adder_28_io_o_adder_0),
    .io_o_adder_1(my_adder_28_io_o_adder_1)
  );
  EdgeAdderSwitch my_adder_29 ( // @[FanNetwork.scala 1474:29]
    .clock(my_adder_29_clock),
    .reset(my_adder_29_reset),
    .io_i_valid(my_adder_29_io_i_valid),
    .io_i_data_bus_0(my_adder_29_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_29_io_i_data_bus_1),
    .io_i_add_en(my_adder_29_io_i_add_en),
    .io_i_cmd(my_adder_29_io_i_cmd),
    .io_o_vn(my_adder_29_io_o_vn),
    .io_o_vn_valid(my_adder_29_io_o_vn_valid),
    .io_o_adder(my_adder_29_io_o_adder)
  );
  EdgeAdderSwitch my_adder_30 ( // @[FanNetwork.scala 1491:29]
    .clock(my_adder_30_clock),
    .reset(my_adder_30_reset),
    .io_i_valid(my_adder_30_io_i_valid),
    .io_i_data_bus_0(my_adder_30_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_30_io_i_data_bus_1),
    .io_i_add_en(my_adder_30_io_i_add_en),
    .io_i_cmd(my_adder_30_io_i_cmd),
    .io_o_vn(my_adder_30_io_o_vn),
    .io_o_vn_valid(my_adder_30_io_o_vn_valid),
    .io_o_adder(my_adder_30_io_o_adder)
  );
  assign io_o_valid_0 = r_lvl_output_ff_valid_128; // @[FanNetwork.scala 1638:19]
  assign io_o_valid_1 = r_lvl_output_ff_valid_129; // @[FanNetwork.scala 1639:19]
  assign io_o_valid_2 = r_lvl_output_ff_valid_130; // @[FanNetwork.scala 1640:19]
  assign io_o_valid_3 = r_lvl_output_ff_valid_131; // @[FanNetwork.scala 1641:19]
  assign io_o_valid_4 = r_lvl_output_ff_valid_132; // @[FanNetwork.scala 1642:19]
  assign io_o_valid_5 = r_lvl_output_ff_valid_133; // @[FanNetwork.scala 1643:19]
  assign io_o_valid_6 = r_lvl_output_ff_valid_134; // @[FanNetwork.scala 1644:19]
  assign io_o_valid_7 = r_lvl_output_ff_valid_135; // @[FanNetwork.scala 1645:19]
  assign io_o_valid_8 = r_lvl_output_ff_valid_136; // @[FanNetwork.scala 1646:19]
  assign io_o_valid_9 = r_lvl_output_ff_valid_137; // @[FanNetwork.scala 1647:19]
  assign io_o_valid_10 = r_lvl_output_ff_valid_138; // @[FanNetwork.scala 1648:20]
  assign io_o_valid_11 = r_lvl_output_ff_valid_139; // @[FanNetwork.scala 1649:20]
  assign io_o_valid_12 = r_lvl_output_ff_valid_140; // @[FanNetwork.scala 1650:20]
  assign io_o_valid_13 = r_lvl_output_ff_valid_141; // @[FanNetwork.scala 1651:20]
  assign io_o_valid_14 = r_lvl_output_ff_valid_142; // @[FanNetwork.scala 1652:20]
  assign io_o_valid_15 = r_final_add2 | r_lvl_output_ff_valid_143; // @[FanNetwork.scala 1653:33 1654:24 1656:25]
  assign io_o_valid_16 = r_lvl_output_ff_valid_144; // @[FanNetwork.scala 1658:20]
  assign io_o_valid_17 = r_lvl_output_ff_valid_145; // @[FanNetwork.scala 1659:20]
  assign io_o_valid_18 = r_lvl_output_ff_valid_146; // @[FanNetwork.scala 1660:20]
  assign io_o_valid_19 = r_lvl_output_ff_valid_147; // @[FanNetwork.scala 1661:20]
  assign io_o_valid_20 = r_lvl_output_ff_valid_148; // @[FanNetwork.scala 1662:20]
  assign io_o_valid_21 = r_lvl_output_ff_valid_149; // @[FanNetwork.scala 1663:20]
  assign io_o_valid_22 = r_lvl_output_ff_valid_150; // @[FanNetwork.scala 1664:20]
  assign io_o_valid_23 = r_lvl_output_ff_valid_151; // @[FanNetwork.scala 1665:20]
  assign io_o_valid_24 = r_lvl_output_ff_valid_152; // @[FanNetwork.scala 1666:20]
  assign io_o_valid_25 = r_lvl_output_ff_valid_153; // @[FanNetwork.scala 1667:20]
  assign io_o_valid_26 = r_lvl_output_ff_valid_154; // @[FanNetwork.scala 1668:20]
  assign io_o_valid_27 = r_lvl_output_ff_valid_155; // @[FanNetwork.scala 1669:20]
  assign io_o_valid_28 = r_lvl_output_ff_valid_156; // @[FanNetwork.scala 1670:20]
  assign io_o_valid_29 = r_lvl_output_ff_valid_157; // @[FanNetwork.scala 1671:20]
  assign io_o_valid_30 = r_lvl_output_ff_valid_158; // @[FanNetwork.scala 1672:20]
  assign io_o_valid_31 = r_lvl_output_ff_valid_159; // @[FanNetwork.scala 1673:20]
  assign io_o_data_bus_0 = r_lvl_output_ff_128; // @[FanNetwork.scala 1557:22]
  assign io_o_data_bus_1 = r_lvl_output_ff_129; // @[FanNetwork.scala 1558:22]
  assign io_o_data_bus_2 = r_lvl_output_ff_130; // @[FanNetwork.scala 1559:22]
  assign io_o_data_bus_3 = r_lvl_output_ff_131; // @[FanNetwork.scala 1560:22]
  assign io_o_data_bus_4 = r_lvl_output_ff_132; // @[FanNetwork.scala 1561:22]
  assign io_o_data_bus_5 = r_lvl_output_ff_133; // @[FanNetwork.scala 1562:22]
  assign io_o_data_bus_6 = r_lvl_output_ff_134; // @[FanNetwork.scala 1563:22]
  assign io_o_data_bus_7 = r_lvl_output_ff_135; // @[FanNetwork.scala 1564:22]
  assign io_o_data_bus_8 = r_lvl_output_ff_136; // @[FanNetwork.scala 1565:22]
  assign io_o_data_bus_9 = r_lvl_output_ff_137; // @[FanNetwork.scala 1566:22]
  assign io_o_data_bus_10 = r_lvl_output_ff_138; // @[FanNetwork.scala 1567:23]
  assign io_o_data_bus_11 = r_lvl_output_ff_139; // @[FanNetwork.scala 1568:23]
  assign io_o_data_bus_12 = r_lvl_output_ff_140; // @[FanNetwork.scala 1569:23]
  assign io_o_data_bus_13 = r_lvl_output_ff_141; // @[FanNetwork.scala 1570:23]
  assign io_o_data_bus_14 = r_lvl_output_ff_142; // @[FanNetwork.scala 1571:23]
  assign io_o_data_bus_15 = r_final_add2 ? r_final_sum : r_lvl_output_ff_143; // @[FanNetwork.scala 1573:33 1574:27 1576:27]
  assign io_o_data_bus_16 = r_lvl_output_ff_144; // @[FanNetwork.scala 1578:23]
  assign io_o_data_bus_17 = r_lvl_output_ff_145; // @[FanNetwork.scala 1579:23]
  assign io_o_data_bus_18 = r_lvl_output_ff_146; // @[FanNetwork.scala 1580:23]
  assign io_o_data_bus_19 = r_lvl_output_ff_147; // @[FanNetwork.scala 1581:23]
  assign io_o_data_bus_20 = r_lvl_output_ff_148; // @[FanNetwork.scala 1582:23]
  assign io_o_data_bus_21 = r_lvl_output_ff_149; // @[FanNetwork.scala 1583:23]
  assign io_o_data_bus_22 = r_lvl_output_ff_150; // @[FanNetwork.scala 1584:23]
  assign io_o_data_bus_23 = r_lvl_output_ff_151; // @[FanNetwork.scala 1585:23]
  assign io_o_data_bus_24 = r_lvl_output_ff_152; // @[FanNetwork.scala 1586:23]
  assign io_o_data_bus_25 = r_lvl_output_ff_153; // @[FanNetwork.scala 1587:23]
  assign io_o_data_bus_26 = r_lvl_output_ff_154; // @[FanNetwork.scala 1588:23]
  assign io_o_data_bus_27 = r_lvl_output_ff_155; // @[FanNetwork.scala 1589:23]
  assign io_o_data_bus_28 = r_lvl_output_ff_156; // @[FanNetwork.scala 1590:23]
  assign io_o_data_bus_29 = r_lvl_output_ff_157; // @[FanNetwork.scala 1591:23]
  assign io_o_data_bus_30 = r_lvl_output_ff_158; // @[FanNetwork.scala 1592:23]
  assign io_o_data_bus_31 = r_lvl_output_ff_159; // @[FanNetwork.scala 1593:23]
  assign io_o_adder_0 = w_fan_lvl_0_0[31:0]; // @[FanNetwork.scala 1709:19]
  assign io_o_adder_1 = w_fan_lvl_1_0[31:0]; // @[FanNetwork.scala 1710:19]
  assign io_o_adder_2 = w_fan_lvl_0_1[31:0]; // @[FanNetwork.scala 1711:19]
  assign io_o_adder_3 = w_fan_lvl_2_0[31:0]; // @[FanNetwork.scala 1712:19]
  assign io_o_adder_4 = w_fan_lvl_0_3[31:0]; // @[FanNetwork.scala 1713:19]
  assign io_o_adder_5 = w_fan_lvl_1_1[31:0]; // @[FanNetwork.scala 1714:19]
  assign io_o_adder_6 = w_fan_lvl_0_5[31:0]; // @[FanNetwork.scala 1715:19]
  assign io_o_adder_7 = w_fan_lvl_3_0[31:0]; // @[FanNetwork.scala 1716:19]
  assign io_o_adder_8 = w_fan_lvl_0_7[31:0]; // @[FanNetwork.scala 1717:19]
  assign io_o_adder_9 = w_fan_lvl_1_3[31:0]; // @[FanNetwork.scala 1718:19]
  assign io_o_adder_10 = w_fan_lvl_0_9[31:0]; // @[FanNetwork.scala 1719:20]
  assign io_o_adder_11 = w_fan_lvl_2_1[31:0]; // @[FanNetwork.scala 1720:20]
  assign io_o_adder_12 = w_fan_lvl_0_11[31:0]; // @[FanNetwork.scala 1721:20]
  assign io_o_adder_13 = w_fan_lvl_1_5[31:0]; // @[FanNetwork.scala 1722:20]
  assign io_o_adder_14 = w_fan_lvl_0_13[31:0]; // @[FanNetwork.scala 1723:20]
  assign io_o_adder_15 = my_adder_15_io_o_adder; // @[FanNetwork.scala 1724:20]
  assign io_o_adder_16 = w_fan_lvl_0_15[31:0]; // @[FanNetwork.scala 1725:20]
  assign io_o_adder_17 = w_fan_lvl_1_7[31:0]; // @[FanNetwork.scala 1726:20]
  assign io_o_adder_18 = w_fan_lvl_0_17[31:0]; // @[FanNetwork.scala 1727:20]
  assign io_o_adder_19 = w_fan_lvl_0_17[31:0]; // @[FanNetwork.scala 1728:20]
  assign io_o_adder_20 = w_fan_lvl_0_19[31:0]; // @[FanNetwork.scala 1729:20]
  assign io_o_adder_21 = w_fan_lvl_1_9[31:0]; // @[FanNetwork.scala 1730:20]
  assign io_o_adder_22 = w_fan_lvl_0_21[31:0]; // @[FanNetwork.scala 1731:20]
  assign io_o_adder_23 = w_fan_lvl_3_1[31:0]; // @[FanNetwork.scala 1732:20]
  assign io_o_adder_24 = w_fan_lvl_0_23[31:0]; // @[FanNetwork.scala 1733:20]
  assign io_o_adder_25 = w_fan_lvl_1_11[31:0]; // @[FanNetwork.scala 1734:20]
  assign io_o_adder_26 = w_fan_lvl_0_25[31:0]; // @[FanNetwork.scala 1735:20]
  assign io_o_adder_27 = w_fan_lvl_2_5[31:0]; // @[FanNetwork.scala 1736:20]
  assign io_o_adder_28 = w_fan_lvl_0_27[31:0]; // @[FanNetwork.scala 1737:20]
  assign io_o_adder_29 = w_fan_lvl_1_13[31:0]; // @[FanNetwork.scala 1738:20]
  assign io_o_adder_30 = w_fan_lvl_0_29[31:0]; // @[FanNetwork.scala 1739:20]
  assign my_adder_0_clock = clock;
  assign my_adder_0_reset = reset;
  assign my_adder_0_io_i_valid = r_valid_0; // @[FanNetwork.scala 986:27]
  assign my_adder_0_io_i_data_bus_0 = {{32'd0}, io_i_data_bus_1}; // @[FanNetwork.scala 987:30]
  assign my_adder_0_io_i_data_bus_1 = {{32'd0}, io_i_data_bus_0}; // @[FanNetwork.scala 987:30]
  assign my_adder_0_io_i_add_en = {{2'd0}, io_i_add_en_bus_0}; // @[FanNetwork.scala 988:28]
  assign my_adder_0_io_i_cmd = {{2'd0}, io_i_cmd_bus_0}; // @[FanNetwork.scala 989:25]
  assign my_adder_1_clock = clock;
  assign my_adder_1_reset = reset;
  assign my_adder_1_io_i_valid = r_valid_1; // @[FanNetwork.scala 999:27]
  assign my_adder_1_io_i_data_bus_0 = w_fan_lvl_0_1[63:0]; // @[FanNetwork.scala 1000:30]
  assign my_adder_1_io_i_data_bus_1 = w_fan_lvl_0_0[63:0]; // @[FanNetwork.scala 1000:30]
  assign my_adder_1_io_i_add_en = {{2'd0}, io_i_add_en_bus_16}; // @[FanNetwork.scala 1001:28]
  assign my_adder_1_io_i_cmd = {{2'd0}, io_i_cmd_bus_16}; // @[FanNetwork.scala 1002:26]
  assign my_adder_2_clock = clock;
  assign my_adder_2_reset = reset;
  assign my_adder_2_io_i_valid = r_valid_0; // @[FanNetwork.scala 1012:27]
  assign my_adder_2_io_i_data_bus_0 = io_i_data_bus_3; // @[FanNetwork.scala 1013:{40,40}]
  assign my_adder_2_io_i_data_bus_1 = io_i_data_bus_2; // @[FanNetwork.scala 1013:{40,40}]
  assign my_adder_2_io_i_add_en = {{2'd0}, io_i_add_en_bus_1}; // @[FanNetwork.scala 1014:28]
  assign my_adder_2_io_i_cmd = io_i_cmd_bus_1; // @[FanNetwork.scala 1015:25]
  assign my_adder_3_clock = clock;
  assign my_adder_3_reset = reset;
  assign my_adder_3_io_i_valid = r_valid_2; // @[FanNetwork.scala 1030:27]
  assign my_adder_3_io_i_data_bus_0 = w_fan_lvl_1_1[63:0]; // @[FanNetwork.scala 1031:32]
  assign my_adder_3_io_i_data_bus_1 = _WIRE_9_1[63:0]; // @[FanNetwork.scala 1031:32]
  assign my_adder_3_io_i_data_bus_2 = _WIRE_9_2[63:0]; // @[FanNetwork.scala 1031:32]
  assign my_adder_3_io_i_data_bus_3 = w_fan_lvl_1_0[63:0]; // @[FanNetwork.scala 1031:32]
  assign my_adder_3_io_i_add_en = {{2'd0}, io_i_add_en_bus_24}; // @[FanNetwork.scala 1032:28]
  assign my_adder_3_io_i_cmd = {{2'd0}, io_i_cmd_bus_24}; // @[FanNetwork.scala 1033:27]
  assign my_adder_3_io_i_sel = _my_adder_3_io_i_sel_T[1:0]; // @[FanNetwork.scala 1034:25]
  assign my_adder_4_clock = clock;
  assign my_adder_4_reset = reset;
  assign my_adder_4_io_i_valid = r_valid_0; // @[FanNetwork.scala 1045:27]
  assign my_adder_4_io_i_data_bus_0 = io_i_data_bus_5; // @[FanNetwork.scala 1046:{40,40}]
  assign my_adder_4_io_i_data_bus_1 = io_i_data_bus_4; // @[FanNetwork.scala 1046:{40,40}]
  assign my_adder_4_io_i_add_en = {{2'd0}, io_i_add_en_bus_2}; // @[FanNetwork.scala 1047:28]
  assign my_adder_4_io_i_cmd = io_i_cmd_bus_2; // @[FanNetwork.scala 1048:26]
  assign my_adder_5_clock = clock;
  assign my_adder_5_reset = reset;
  assign my_adder_5_io_i_valid = r_valid_1; // @[FanNetwork.scala 1062:27]
  assign my_adder_5_io_i_data_bus_0 = w_fan_lvl_0_5[31:0]; // @[FanNetwork.scala 1063:30]
  assign my_adder_5_io_i_data_bus_1 = w_fan_lvl_0_4[31:0]; // @[FanNetwork.scala 1063:30]
  assign my_adder_5_io_i_add_en = {{2'd0}, io_i_add_en_bus_17}; // @[FanNetwork.scala 1064:28]
  assign my_adder_5_io_i_cmd = io_i_cmd_bus_17; // @[FanNetwork.scala 1065:26]
  assign my_adder_6_clock = clock;
  assign my_adder_6_reset = reset;
  assign my_adder_6_io_i_valid = r_valid_0; // @[FanNetwork.scala 1078:27]
  assign my_adder_6_io_i_data_bus_0 = io_i_data_bus_7; // @[FanNetwork.scala 1079:{40,40}]
  assign my_adder_6_io_i_data_bus_1 = io_i_data_bus_6; // @[FanNetwork.scala 1079:{40,40}]
  assign my_adder_6_io_i_add_en = {{2'd0}, io_i_add_en_bus_3}; // @[FanNetwork.scala 1080:28]
  assign my_adder_6_io_i_cmd = io_i_cmd_bus_3; // @[FanNetwork.scala 1081:25]
  assign my_adder_7_clock = clock;
  assign my_adder_7_reset = reset;
  assign my_adder_7_io_i_valid = r_valid_3; // @[FanNetwork.scala 1094:27]
  assign my_adder_7_io_i_data_bus_0 = w_fan_lvl_2_1[63:0]; // @[FanNetwork.scala 1096:30]
  assign my_adder_7_io_i_data_bus_1 = _WIRE_13_1[63:0]; // @[FanNetwork.scala 1096:30]
  assign my_adder_7_io_i_data_bus_2 = _WIRE_13_2[63:0]; // @[FanNetwork.scala 1096:30]
  assign my_adder_7_io_i_data_bus_3 = _WIRE_13_3[63:0]; // @[FanNetwork.scala 1096:30]
  assign my_adder_7_io_i_data_bus_4 = _WIRE_13_4[63:0]; // @[FanNetwork.scala 1096:30]
  assign my_adder_7_io_i_data_bus_5 = w_fan_lvl_2_0[63:0]; // @[FanNetwork.scala 1096:30]
  assign my_adder_7_io_i_add_en = {{2'd0}, io_i_add_en_bus_28}; // @[FanNetwork.scala 1097:28]
  assign my_adder_7_io_i_cmd = {{2'd0}, io_i_cmd_bus_28}; // @[FanNetwork.scala 1098:25]
  assign my_adder_7_io_i_sel = _my_adder_7_io_i_sel_T[3:0]; // @[FanNetwork.scala 1099:21]
  assign my_adder_8_clock = clock;
  assign my_adder_8_reset = reset;
  assign my_adder_8_io_i_valid = r_valid_0; // @[FanNetwork.scala 1111:27]
  assign my_adder_8_io_i_data_bus_0 = io_i_data_bus_9; // @[FanNetwork.scala 1112:{40,40}]
  assign my_adder_8_io_i_data_bus_1 = io_i_data_bus_8; // @[FanNetwork.scala 1112:{40,40}]
  assign my_adder_8_io_i_add_en = {{2'd0}, io_i_add_en_bus_4}; // @[FanNetwork.scala 1113:28]
  assign my_adder_8_io_i_cmd = io_i_cmd_bus_4; // @[FanNetwork.scala 1114:25]
  assign my_adder_9_clock = clock;
  assign my_adder_9_reset = reset;
  assign my_adder_9_io_i_valid = r_valid_1; // @[FanNetwork.scala 1127:27]
  assign my_adder_9_io_i_data_bus_0 = w_fan_lvl_0_9[31:0]; // @[FanNetwork.scala 1128:30]
  assign my_adder_9_io_i_data_bus_1 = w_fan_lvl_0_8[31:0]; // @[FanNetwork.scala 1128:30]
  assign my_adder_9_io_i_add_en = {{2'd0}, io_i_add_en_bus_18}; // @[FanNetwork.scala 1129:28]
  assign my_adder_9_io_i_cmd = io_i_cmd_bus_18; // @[FanNetwork.scala 1130:25]
  assign my_adder_10_clock = clock;
  assign my_adder_10_reset = reset;
  assign my_adder_10_io_i_valid = r_valid_0; // @[FanNetwork.scala 1143:28]
  assign my_adder_10_io_i_data_bus_0 = io_i_data_bus_11; // @[FanNetwork.scala 1144:{41,41}]
  assign my_adder_10_io_i_data_bus_1 = io_i_data_bus_10; // @[FanNetwork.scala 1144:{41,41}]
  assign my_adder_10_io_i_add_en = {{2'd0}, io_i_add_en_bus_5}; // @[FanNetwork.scala 1145:29]
  assign my_adder_10_io_i_cmd = io_i_cmd_bus_5; // @[FanNetwork.scala 1146:27]
  assign my_adder_11_clock = clock;
  assign my_adder_11_reset = reset;
  assign my_adder_11_io_i_valid = r_valid_2; // @[FanNetwork.scala 1160:28]
  assign my_adder_11_io_i_data_bus_0 = w_fan_lvl_1_5[31:0]; // @[FanNetwork.scala 1161:31]
  assign my_adder_11_io_i_data_bus_1 = _WIRE_17_1[31:0]; // @[FanNetwork.scala 1161:31]
  assign my_adder_11_io_i_data_bus_2 = _WIRE_17_2[31:0]; // @[FanNetwork.scala 1161:31]
  assign my_adder_11_io_i_data_bus_3 = w_fan_lvl_1_4[31:0]; // @[FanNetwork.scala 1161:31]
  assign my_adder_11_io_i_add_en = {{2'd0}, io_i_add_en_bus_25}; // @[FanNetwork.scala 1163:29]
  assign my_adder_11_io_i_cmd = io_i_cmd_bus_25; // @[FanNetwork.scala 1164:26]
  assign my_adder_11_io_i_sel = _my_adder_11_io_i_sel_T[1:0]; // @[FanNetwork.scala 1165:26]
  assign my_adder_12_clock = clock;
  assign my_adder_12_reset = reset;
  assign my_adder_12_io_i_valid = r_valid_0; // @[FanNetwork.scala 1179:28]
  assign my_adder_12_io_i_data_bus_0 = io_i_data_bus_13; // @[FanNetwork.scala 1180:{41,41}]
  assign my_adder_12_io_i_data_bus_1 = io_i_data_bus_12; // @[FanNetwork.scala 1180:{41,41}]
  assign my_adder_12_io_i_add_en = {{2'd0}, io_i_add_en_bus_6}; // @[FanNetwork.scala 1181:29]
  assign my_adder_12_io_i_cmd = io_i_cmd_bus_6; // @[FanNetwork.scala 1182:27]
  assign my_adder_13_clock = clock;
  assign my_adder_13_reset = reset;
  assign my_adder_13_io_i_valid = r_valid_1; // @[FanNetwork.scala 1196:28]
  assign my_adder_13_io_i_data_bus_0 = w_fan_lvl_0_12[31:0]; // @[FanNetwork.scala 1197:31]
  assign my_adder_13_io_i_data_bus_1 = w_fan_lvl_0_11[31:0]; // @[FanNetwork.scala 1197:31]
  assign my_adder_13_io_i_add_en = {{2'd0}, io_i_add_en_bus_19}; // @[FanNetwork.scala 1198:29]
  assign my_adder_13_io_i_cmd = io_i_cmd_bus_19; // @[FanNetwork.scala 1199:26]
  assign my_adder_14_clock = clock;
  assign my_adder_14_reset = reset;
  assign my_adder_14_io_i_valid = r_valid_0; // @[FanNetwork.scala 1213:28]
  assign my_adder_14_io_i_data_bus_0 = io_i_data_bus_15; // @[FanNetwork.scala 1214:{41,41}]
  assign my_adder_14_io_i_data_bus_1 = io_i_data_bus_14; // @[FanNetwork.scala 1214:{41,41}]
  assign my_adder_14_io_i_add_en = {{2'd0}, io_i_add_en_bus_7}; // @[FanNetwork.scala 1215:29]
  assign my_adder_14_io_i_cmd = io_i_cmd_bus_7; // @[FanNetwork.scala 1216:26]
  assign my_adder_15_clock = clock;
  assign my_adder_15_reset = reset;
  assign my_adder_15_io_i_valid = r_valid_4; // @[FanNetwork.scala 1230:28]
  assign my_adder_15_io_i_data_bus_0 = {{32'd0}, my_adder_23_io_o_adder}; // @[FanNetwork.scala 1231:{41,41}]
  assign my_adder_15_io_i_data_bus_1 = {{32'd0}, r_fan_ff_lvl_2_to_4_1}; // @[FanNetwork.scala 1231:{41,41}]
  assign my_adder_15_io_i_data_bus_2 = {{32'd0}, r_fan_ff_lvl_1_to_4_1}; // @[FanNetwork.scala 1231:{41,41}]
  assign my_adder_15_io_i_data_bus_3 = {{32'd0}, r_fan_ff_lvl_0_to_4_1}; // @[FanNetwork.scala 1231:{41,41}]
  assign my_adder_15_io_i_data_bus_4 = {{32'd0}, r_fan_ff_lvl_0_to_4_0}; // @[FanNetwork.scala 1231:{41,41}]
  assign my_adder_15_io_i_data_bus_5 = {{32'd0}, r_fan_ff_lvl_1_to_4_0}; // @[FanNetwork.scala 1231:{41,41}]
  assign my_adder_15_io_i_data_bus_6 = {{32'd0}, r_fan_ff_lvl_2_to_4_0}; // @[FanNetwork.scala 1231:{41,41}]
  assign my_adder_15_io_i_data_bus_7 = {{32'd0}, my_adder_7_io_o_adder}; // @[FanNetwork.scala 1231:{41,41}]
  assign my_adder_15_io_i_add_en = {{2'd0}, io_i_add_en_bus_30}; // @[FanNetwork.scala 1233:29]
  assign my_adder_15_io_i_cmd = {{2'd0}, io_i_cmd_bus_30}; // @[FanNetwork.scala 1234:26]
  assign my_adder_15_io_i_sel = _my_adder_15_io_i_sel_T[3:0]; // @[FanNetwork.scala 1235:26]
  assign my_adder_16_clock = clock;
  assign my_adder_16_reset = reset;
  assign my_adder_16_io_i_valid = r_valid_0; // @[FanNetwork.scala 1247:28]
  assign my_adder_16_io_i_data_bus_0 = io_i_data_bus_17; // @[FanNetwork.scala 1248:{41,41}]
  assign my_adder_16_io_i_data_bus_1 = io_i_data_bus_16; // @[FanNetwork.scala 1248:{41,41}]
  assign my_adder_16_io_i_add_en = {{2'd0}, io_i_add_en_bus_8}; // @[FanNetwork.scala 1249:29]
  assign my_adder_16_io_i_cmd = io_i_cmd_bus_8; // @[FanNetwork.scala 1250:26]
  assign my_adder_17_clock = clock;
  assign my_adder_17_reset = reset;
  assign my_adder_17_io_i_valid = r_valid_1; // @[FanNetwork.scala 1264:28]
  assign my_adder_17_io_i_data_bus_0 = w_fan_lvl_0_16[31:0]; // @[FanNetwork.scala 1265:31]
  assign my_adder_17_io_i_data_bus_1 = w_fan_lvl_0_15[31:0]; // @[FanNetwork.scala 1265:31]
  assign my_adder_17_io_i_add_en = {{2'd0}, io_i_add_en_bus_20}; // @[FanNetwork.scala 1266:29]
  assign my_adder_17_io_i_cmd = io_i_cmd_bus_20; // @[FanNetwork.scala 1267:26]
  assign my_adder_18_clock = clock;
  assign my_adder_18_reset = reset;
  assign my_adder_18_io_i_valid = r_valid_0; // @[FanNetwork.scala 1281:28]
  assign my_adder_18_io_i_data_bus_0 = io_i_data_bus_19; // @[FanNetwork.scala 1282:{41,41}]
  assign my_adder_18_io_i_data_bus_1 = io_i_data_bus_18; // @[FanNetwork.scala 1282:{41,41}]
  assign my_adder_18_io_i_add_en = {{2'd0}, io_i_add_en_bus_9}; // @[FanNetwork.scala 1283:29]
  assign my_adder_18_io_i_cmd = io_i_cmd_bus_9; // @[FanNetwork.scala 1284:26]
  assign my_adder_19_clock = clock;
  assign my_adder_19_reset = reset;
  assign my_adder_19_io_i_valid = r_valid_2; // @[FanNetwork.scala 1298:28]
  assign my_adder_19_io_i_data_bus_0 = w_fan_lvl_1_9[31:0]; // @[FanNetwork.scala 1299:32]
  assign my_adder_19_io_i_data_bus_1 = _WIRE_25_1[31:0]; // @[FanNetwork.scala 1299:32]
  assign my_adder_19_io_i_data_bus_2 = _WIRE_25_2[31:0]; // @[FanNetwork.scala 1299:32]
  assign my_adder_19_io_i_data_bus_3 = w_fan_lvl_1_8[31:0]; // @[FanNetwork.scala 1299:32]
  assign my_adder_19_io_i_add_en = {{2'd0}, io_i_add_en_bus_26}; // @[FanNetwork.scala 1300:29]
  assign my_adder_19_io_i_cmd = io_i_cmd_bus_26; // @[FanNetwork.scala 1301:26]
  assign my_adder_19_io_i_sel = _my_adder_19_io_i_sel_T[1:0]; // @[FanNetwork.scala 1302:26]
  assign my_adder_20_clock = clock;
  assign my_adder_20_reset = reset;
  assign my_adder_20_io_i_valid = r_valid_0; // @[FanNetwork.scala 1316:28]
  assign my_adder_20_io_i_data_bus_0 = io_i_data_bus_21; // @[FanNetwork.scala 1317:{41,41}]
  assign my_adder_20_io_i_data_bus_1 = io_i_data_bus_20; // @[FanNetwork.scala 1317:{41,41}]
  assign my_adder_20_io_i_add_en = {{2'd0}, io_i_add_en_bus_10}; // @[FanNetwork.scala 1318:29]
  assign my_adder_20_io_i_cmd = io_i_cmd_bus_10; // @[FanNetwork.scala 1319:26]
  assign my_adder_21_clock = clock;
  assign my_adder_21_reset = reset;
  assign my_adder_21_io_i_valid = r_valid_1; // @[FanNetwork.scala 1335:28]
  assign my_adder_21_io_i_data_bus_0 = w_fan_lvl_0_20[31:0]; // @[FanNetwork.scala 1336:31]
  assign my_adder_21_io_i_data_bus_1 = w_fan_lvl_0_19[31:0]; // @[FanNetwork.scala 1336:31]
  assign my_adder_21_io_i_add_en = {{2'd0}, io_i_add_en_bus_21}; // @[FanNetwork.scala 1337:29]
  assign my_adder_21_io_i_cmd = io_i_cmd_bus_21; // @[FanNetwork.scala 1338:27]
  assign my_adder_22_clock = clock;
  assign my_adder_22_reset = reset;
  assign my_adder_22_io_i_valid = r_valid_0; // @[FanNetwork.scala 1353:28]
  assign my_adder_22_io_i_data_bus_0 = io_i_data_bus_23; // @[FanNetwork.scala 1354:{41,41}]
  assign my_adder_22_io_i_data_bus_1 = io_i_data_bus_22; // @[FanNetwork.scala 1354:{41,41}]
  assign my_adder_22_io_i_add_en = {{2'd0}, io_i_add_en_bus_11}; // @[FanNetwork.scala 1355:29]
  assign my_adder_22_io_i_cmd = io_i_cmd_bus_11; // @[FanNetwork.scala 1356:26]
  assign my_adder_23_clock = clock;
  assign my_adder_23_reset = reset;
  assign my_adder_23_io_i_valid = r_valid_3; // @[FanNetwork.scala 1370:28]
  assign my_adder_23_io_i_data_bus_0 = w_fan_lvl_2_5[63:0]; // @[FanNetwork.scala 1371:31]
  assign my_adder_23_io_i_data_bus_1 = _WIRE_29_1[63:0]; // @[FanNetwork.scala 1371:31]
  assign my_adder_23_io_i_data_bus_2 = _WIRE_29_2[63:0]; // @[FanNetwork.scala 1371:31]
  assign my_adder_23_io_i_data_bus_3 = _WIRE_29_3[63:0]; // @[FanNetwork.scala 1371:31]
  assign my_adder_23_io_i_data_bus_4 = _WIRE_29_4[63:0]; // @[FanNetwork.scala 1371:31]
  assign my_adder_23_io_i_data_bus_5 = w_fan_lvl_2_4[63:0]; // @[FanNetwork.scala 1371:31]
  assign my_adder_23_io_i_add_en = {{2'd0}, io_i_add_en_bus_29}; // @[FanNetwork.scala 1372:29]
  assign my_adder_23_io_i_cmd = {{2'd0}, io_i_cmd_bus_29}; // @[FanNetwork.scala 1373:26]
  assign my_adder_23_io_i_sel = _my_adder_23_io_i_sel_T[3:0]; // @[FanNetwork.scala 1374:26]
  assign my_adder_24_clock = clock;
  assign my_adder_24_reset = reset;
  assign my_adder_24_io_i_valid = r_valid_0; // @[FanNetwork.scala 1385:28]
  assign my_adder_24_io_i_data_bus_0 = io_i_data_bus_25; // @[FanNetwork.scala 1386:{41,41}]
  assign my_adder_24_io_i_data_bus_1 = io_i_data_bus_24; // @[FanNetwork.scala 1386:{41,41}]
  assign my_adder_24_io_i_add_en = {{2'd0}, io_i_add_en_bus_12}; // @[FanNetwork.scala 1387:29]
  assign my_adder_24_io_i_cmd = io_i_cmd_bus_12; // @[FanNetwork.scala 1388:26]
  assign my_adder_25_clock = clock;
  assign my_adder_25_reset = reset;
  assign my_adder_25_io_i_valid = r_valid_1; // @[FanNetwork.scala 1403:28]
  assign my_adder_25_io_i_data_bus_0 = w_fan_lvl_0_24[31:0]; // @[FanNetwork.scala 1404:31]
  assign my_adder_25_io_i_data_bus_1 = w_fan_lvl_0_23[31:0]; // @[FanNetwork.scala 1404:31]
  assign my_adder_25_io_i_add_en = {{2'd0}, io_i_add_en_bus_22}; // @[FanNetwork.scala 1405:29]
  assign my_adder_25_io_i_cmd = io_i_cmd_bus_22; // @[FanNetwork.scala 1406:26]
  assign my_adder_26_clock = clock;
  assign my_adder_26_reset = reset;
  assign my_adder_26_io_i_valid = r_valid_0; // @[FanNetwork.scala 1422:28]
  assign my_adder_26_io_i_data_bus_0 = io_i_data_bus_27; // @[FanNetwork.scala 1423:{41,41}]
  assign my_adder_26_io_i_data_bus_1 = io_i_data_bus_26; // @[FanNetwork.scala 1423:{41,41}]
  assign my_adder_26_io_i_add_en = {{2'd0}, io_i_add_en_bus_13}; // @[FanNetwork.scala 1424:29]
  assign my_adder_26_io_i_cmd = io_i_cmd_bus_13; // @[FanNetwork.scala 1425:26]
  assign my_adder_27_clock = clock;
  assign my_adder_27_reset = reset;
  assign my_adder_27_io_i_valid = r_valid_2; // @[FanNetwork.scala 1439:28]
  assign my_adder_27_io_i_data_bus_0 = w_fan_lvl_1_13[63:0]; // @[FanNetwork.scala 1440:31]
  assign my_adder_27_io_i_data_bus_1 = _WIRE_33_1[63:0]; // @[FanNetwork.scala 1440:31]
  assign my_adder_27_io_i_data_bus_2 = _WIRE_33_2[63:0]; // @[FanNetwork.scala 1440:31]
  assign my_adder_27_io_i_data_bus_3 = w_fan_lvl_1_12[63:0]; // @[FanNetwork.scala 1440:31]
  assign my_adder_27_io_i_add_en = {{2'd0}, io_i_add_en_bus_27}; // @[FanNetwork.scala 1441:29]
  assign my_adder_27_io_i_cmd = {{2'd0}, io_i_cmd_bus_27}; // @[FanNetwork.scala 1442:26]
  assign my_adder_27_io_i_sel = _my_adder_27_io_i_sel_T[1:0]; // @[FanNetwork.scala 1443:26]
  assign my_adder_28_clock = clock;
  assign my_adder_28_reset = reset;
  assign my_adder_28_io_i_valid = r_valid_0; // @[FanNetwork.scala 1458:28]
  assign my_adder_28_io_i_data_bus_0 = io_i_data_bus_29; // @[FanNetwork.scala 1459:{41,41}]
  assign my_adder_28_io_i_data_bus_1 = io_i_data_bus_28; // @[FanNetwork.scala 1459:{41,41}]
  assign my_adder_28_io_i_add_en = {{2'd0}, io_i_add_en_bus_14}; // @[FanNetwork.scala 1460:29]
  assign my_adder_28_io_i_cmd = io_i_cmd_bus_14; // @[FanNetwork.scala 1461:27]
  assign my_adder_29_clock = clock;
  assign my_adder_29_reset = reset;
  assign my_adder_29_io_i_valid = r_valid_1; // @[FanNetwork.scala 1476:28]
  assign my_adder_29_io_i_data_bus_0 = w_fan_lvl_0_28[63:0]; // @[FanNetwork.scala 1477:31]
  assign my_adder_29_io_i_data_bus_1 = w_fan_lvl_0_27[63:0]; // @[FanNetwork.scala 1477:31]
  assign my_adder_29_io_i_add_en = {{2'd0}, io_i_add_en_bus_23}; // @[FanNetwork.scala 1478:29]
  assign my_adder_29_io_i_cmd = {{2'd0}, io_i_cmd_bus_23}; // @[FanNetwork.scala 1479:26]
  assign my_adder_30_clock = clock;
  assign my_adder_30_reset = reset;
  assign my_adder_30_io_i_valid = r_valid_0; // @[FanNetwork.scala 1493:28]
  assign my_adder_30_io_i_data_bus_0 = {{32'd0}, io_i_data_bus_31}; // @[FanNetwork.scala 1494:31]
  assign my_adder_30_io_i_data_bus_1 = {{32'd0}, io_i_data_bus_30}; // @[FanNetwork.scala 1494:31]
  assign my_adder_30_io_i_add_en = {{2'd0}, io_i_add_en_bus_15}; // @[FanNetwork.scala 1495:29]
  assign my_adder_30_io_i_cmd = {{2'd0}, io_i_cmd_bus_15}; // @[FanNetwork.scala 1496:26]
  always @(posedge clock) begin
    if (reset) begin // @[FanNetwork.scala 27:38]
      r_fan_ff_lvl_0_to_4_0 <= 32'h0; // @[FanNetwork.scala 27:38]
    end else begin
      r_fan_ff_lvl_0_to_4_0 <= r_fan_ff_lvl_0_to_3_2; // @[FanNetwork.scala 55:25]
    end
    if (reset) begin // @[FanNetwork.scala 27:38]
      r_fan_ff_lvl_0_to_4_1 <= 32'h0; // @[FanNetwork.scala 27:38]
    end else begin
      r_fan_ff_lvl_0_to_4_1 <= r_fan_ff_lvl_0_to_3_3; // @[FanNetwork.scala 55:25]
    end
    if (reset) begin // @[FanNetwork.scala 28:38]
      r_fan_ff_lvl_0_to_3_0 <= 32'h0; // @[FanNetwork.scala 28:38]
    end else begin
      r_fan_ff_lvl_0_to_3_0 <= r_fan_ff_lvl_0_to_2_2; // @[FanNetwork.scala 54:25]
    end
    if (reset) begin // @[FanNetwork.scala 28:38]
      r_fan_ff_lvl_0_to_3_1 <= 32'h0; // @[FanNetwork.scala 28:38]
    end else begin
      r_fan_ff_lvl_0_to_3_1 <= r_fan_ff_lvl_0_to_2_3; // @[FanNetwork.scala 54:25]
    end
    if (reset) begin // @[FanNetwork.scala 28:38]
      r_fan_ff_lvl_0_to_3_2 <= 32'h0; // @[FanNetwork.scala 28:38]
    end else begin
      r_fan_ff_lvl_0_to_3_2 <= r_fan_ff_lvl_0_to_2_6; // @[FanNetwork.scala 54:25]
    end
    if (reset) begin // @[FanNetwork.scala 28:38]
      r_fan_ff_lvl_0_to_3_3 <= 32'h0; // @[FanNetwork.scala 28:38]
    end else begin
      r_fan_ff_lvl_0_to_3_3 <= r_fan_ff_lvl_0_to_2_7; // @[FanNetwork.scala 54:25]
    end
    if (reset) begin // @[FanNetwork.scala 28:38]
      r_fan_ff_lvl_0_to_3_4 <= 32'h0; // @[FanNetwork.scala 28:38]
    end else begin
      r_fan_ff_lvl_0_to_3_4 <= r_fan_ff_lvl_0_to_2_10; // @[FanNetwork.scala 54:25]
    end
    if (reset) begin // @[FanNetwork.scala 28:38]
      r_fan_ff_lvl_0_to_3_5 <= 32'h0; // @[FanNetwork.scala 28:38]
    end else begin
      r_fan_ff_lvl_0_to_3_5 <= r_fan_ff_lvl_0_to_2_11; // @[FanNetwork.scala 54:25]
    end
    r_fan_ff_lvl_0_to_2_0 <= _GEN_239[31:0]; // @[FanNetwork.scala 29:{38,38} 53:25]
    r_fan_ff_lvl_0_to_2_1 <= _GEN_240[31:0]; // @[FanNetwork.scala 29:{38,38} 53:25]
    r_fan_ff_lvl_0_to_2_2 <= _GEN_241[31:0]; // @[FanNetwork.scala 29:{38,38} 53:25]
    r_fan_ff_lvl_0_to_2_3 <= _GEN_242[31:0]; // @[FanNetwork.scala 29:{38,38} 53:25]
    r_fan_ff_lvl_0_to_2_4 <= _GEN_243[31:0]; // @[FanNetwork.scala 29:{38,38} 53:25]
    r_fan_ff_lvl_0_to_2_5 <= _GEN_244[31:0]; // @[FanNetwork.scala 29:{38,38} 53:25]
    r_fan_ff_lvl_0_to_2_6 <= _GEN_245[31:0]; // @[FanNetwork.scala 29:{38,38} 53:25]
    r_fan_ff_lvl_0_to_2_7 <= _GEN_246[31:0]; // @[FanNetwork.scala 29:{38,38} 53:25]
    r_fan_ff_lvl_0_to_2_8 <= _GEN_247[31:0]; // @[FanNetwork.scala 29:{38,38} 53:25]
    r_fan_ff_lvl_0_to_2_9 <= _GEN_248[31:0]; // @[FanNetwork.scala 29:{38,38} 53:25]
    r_fan_ff_lvl_0_to_2_10 <= _GEN_249[31:0]; // @[FanNetwork.scala 29:{38,38} 53:25]
    r_fan_ff_lvl_0_to_2_11 <= _GEN_250[31:0]; // @[FanNetwork.scala 29:{38,38} 53:25]
    r_fan_ff_lvl_0_to_2_12 <= _GEN_251[31:0]; // @[FanNetwork.scala 29:{38,38} 53:25]
    r_fan_ff_lvl_0_to_2_13 <= _GEN_252[31:0]; // @[FanNetwork.scala 29:{38,38} 53:25]
    if (reset) begin // @[FanNetwork.scala 30:38]
      r_fan_ff_lvl_1_to_4_0 <= 32'h0; // @[FanNetwork.scala 30:38]
    end else begin
      r_fan_ff_lvl_1_to_4_0 <= r_fan_ff_lvl_1_to_3_2; // @[FanNetwork.scala 56:25]
    end
    if (reset) begin // @[FanNetwork.scala 30:38]
      r_fan_ff_lvl_1_to_4_1 <= 32'h0; // @[FanNetwork.scala 30:38]
    end else begin
      r_fan_ff_lvl_1_to_4_1 <= r_fan_ff_lvl_1_to_3_3; // @[FanNetwork.scala 56:25]
    end
    r_fan_ff_lvl_1_to_3_0 <= _GEN_253[31:0]; // @[FanNetwork.scala 31:{38,38} 57:25]
    r_fan_ff_lvl_1_to_3_1 <= _GEN_254[31:0]; // @[FanNetwork.scala 31:{38,38} 57:25]
    r_fan_ff_lvl_1_to_3_2 <= _GEN_255[31:0]; // @[FanNetwork.scala 31:{38,38} 57:25]
    r_fan_ff_lvl_1_to_3_3 <= _GEN_256[31:0]; // @[FanNetwork.scala 31:{38,38} 57:25]
    r_fan_ff_lvl_1_to_3_4 <= _GEN_257[31:0]; // @[FanNetwork.scala 31:{38,38} 57:25]
    r_fan_ff_lvl_1_to_3_5 <= _GEN_258[31:0]; // @[FanNetwork.scala 31:{38,38} 57:25]
    r_fan_ff_lvl_2_to_4_0 <= _GEN_259[31:0]; // @[FanNetwork.scala 32:{38,38} 58:25]
    r_fan_ff_lvl_2_to_4_1 <= _GEN_260[31:0]; // @[FanNetwork.scala 32:{38,38} 58:25]
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_0 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_0_valid_1 & w_vn_lvl_0_valid_0) begin // @[FanNetwork.scala 63:77]
      r_lvl_output_ff_0 <= w_vn_lvl_0_0; // @[FanNetwork.scala 65:24]
    end else if (w_vn_lvl_0_valid_1 & ~w_vn_lvl_0_valid_0) begin // @[FanNetwork.scala 68:83]
      r_lvl_output_ff_0 <= 32'h0; // @[FanNetwork.scala 70:24]
    end else if (~w_vn_lvl_0_valid_1 & w_vn_lvl_0_valid_0) begin // @[FanNetwork.scala 73:83]
      r_lvl_output_ff_0 <= w_vn_lvl_0_0; // @[FanNetwork.scala 75:24]
    end else begin
      r_lvl_output_ff_0 <= 32'h0; // @[FanNetwork.scala 80:24]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_1 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_0_valid_1 & w_vn_lvl_0_valid_0) begin // @[FanNetwork.scala 63:77]
      r_lvl_output_ff_1 <= w_vn_lvl_0_1; // @[FanNetwork.scala 64:24]
    end else if (w_vn_lvl_0_valid_1 & ~w_vn_lvl_0_valid_0) begin // @[FanNetwork.scala 68:83]
      r_lvl_output_ff_1 <= w_vn_lvl_0_1; // @[FanNetwork.scala 69:24]
    end else begin
      r_lvl_output_ff_1 <= 32'h0;
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_2 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_0_valid_3 & w_vn_lvl_0_valid_2) begin // @[FanNetwork.scala 85:77]
      r_lvl_output_ff_2 <= w_vn_lvl_0_2; // @[FanNetwork.scala 87:28]
    end else if (w_vn_lvl_0_valid_3 & ~w_vn_lvl_0_valid_2) begin // @[FanNetwork.scala 90:83]
      r_lvl_output_ff_2 <= 32'h0; // @[FanNetwork.scala 92:28]
    end else if (~w_vn_lvl_0_valid_3 & w_vn_lvl_0_valid_2) begin // @[FanNetwork.scala 95:83]
      r_lvl_output_ff_2 <= w_vn_lvl_0_2; // @[FanNetwork.scala 97:28]
    end else begin
      r_lvl_output_ff_2 <= 32'h0; // @[FanNetwork.scala 102:28]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_3 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_0_valid_3 & w_vn_lvl_0_valid_2) begin // @[FanNetwork.scala 85:77]
      r_lvl_output_ff_3 <= w_vn_lvl_0_3; // @[FanNetwork.scala 86:28]
    end else if (w_vn_lvl_0_valid_3 & ~w_vn_lvl_0_valid_2) begin // @[FanNetwork.scala 90:83]
      r_lvl_output_ff_3 <= w_vn_lvl_0_3; // @[FanNetwork.scala 91:28]
    end else begin
      r_lvl_output_ff_3 <= 32'h0;
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_4 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_0_valid_5 & w_vn_lvl_0_valid_4) begin // @[FanNetwork.scala 107:77]
      r_lvl_output_ff_4 <= w_vn_lvl_0_4; // @[FanNetwork.scala 109:24]
    end else if (w_vn_lvl_0_valid_5 & ~w_vn_lvl_0_valid_4) begin // @[FanNetwork.scala 112:83]
      r_lvl_output_ff_4 <= 32'h0; // @[FanNetwork.scala 114:24]
    end else if (~w_vn_lvl_0_valid_5 & w_vn_lvl_0_valid_4) begin // @[FanNetwork.scala 117:83]
      r_lvl_output_ff_4 <= w_vn_lvl_0_4; // @[FanNetwork.scala 119:24]
    end else begin
      r_lvl_output_ff_4 <= 32'h0; // @[FanNetwork.scala 124:24]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_5 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_0_valid_5 & w_vn_lvl_0_valid_4) begin // @[FanNetwork.scala 107:77]
      r_lvl_output_ff_5 <= w_vn_lvl_0_5; // @[FanNetwork.scala 108:24]
    end else if (w_vn_lvl_0_valid_5 & ~w_vn_lvl_0_valid_4) begin // @[FanNetwork.scala 112:83]
      r_lvl_output_ff_5 <= w_vn_lvl_0_5; // @[FanNetwork.scala 113:24]
    end else begin
      r_lvl_output_ff_5 <= 32'h0;
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_6 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_0_valid_7 & w_vn_lvl_0_valid_6) begin // @[FanNetwork.scala 130:77]
      r_lvl_output_ff_6 <= w_vn_lvl_0_6; // @[FanNetwork.scala 132:24]
    end else if (w_vn_lvl_0_valid_7 & ~w_vn_lvl_0_valid_6) begin // @[FanNetwork.scala 135:83]
      r_lvl_output_ff_6 <= 32'h0; // @[FanNetwork.scala 137:24]
    end else if (~w_vn_lvl_0_valid_7 & w_vn_lvl_0_valid_6) begin // @[FanNetwork.scala 140:83]
      r_lvl_output_ff_6 <= w_vn_lvl_0_6; // @[FanNetwork.scala 142:24]
    end else begin
      r_lvl_output_ff_6 <= 32'h0; // @[FanNetwork.scala 147:24]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_7 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_0_valid_7 & w_vn_lvl_0_valid_6) begin // @[FanNetwork.scala 130:77]
      r_lvl_output_ff_7 <= w_vn_lvl_0_7; // @[FanNetwork.scala 131:24]
    end else if (w_vn_lvl_0_valid_7 & ~w_vn_lvl_0_valid_6) begin // @[FanNetwork.scala 135:83]
      r_lvl_output_ff_7 <= w_vn_lvl_0_7; // @[FanNetwork.scala 136:24]
    end else begin
      r_lvl_output_ff_7 <= 32'h0;
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_8 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_0_valid_9 & w_vn_lvl_0_valid_8) begin // @[FanNetwork.scala 153:61]
      r_lvl_output_ff_8 <= w_vn_lvl_0_8; // @[FanNetwork.scala 155:24]
    end else if (w_vn_lvl_0_valid_9 & ~w_vn_lvl_0_valid_8) begin // @[FanNetwork.scala 158:68]
      r_lvl_output_ff_8 <= 32'h0; // @[FanNetwork.scala 160:24]
    end else if (~w_vn_lvl_0_valid_9 & w_vn_lvl_0_valid_8) begin // @[FanNetwork.scala 163:68]
      r_lvl_output_ff_8 <= w_vn_lvl_0_8; // @[FanNetwork.scala 165:24]
    end else begin
      r_lvl_output_ff_8 <= 32'h0; // @[FanNetwork.scala 170:24]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_9 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_0_valid_9 & w_vn_lvl_0_valid_8) begin // @[FanNetwork.scala 153:61]
      r_lvl_output_ff_9 <= w_vn_lvl_0_9; // @[FanNetwork.scala 154:24]
    end else if (w_vn_lvl_0_valid_9 & ~w_vn_lvl_0_valid_8) begin // @[FanNetwork.scala 158:68]
      r_lvl_output_ff_9 <= w_vn_lvl_0_9; // @[FanNetwork.scala 159:24]
    end else begin
      r_lvl_output_ff_9 <= 32'h0;
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_10 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_0_valid_11 & w_vn_lvl_0_valid_10) begin // @[FanNetwork.scala 176:63]
      r_lvl_output_ff_10 <= w_vn_lvl_0_10; // @[FanNetwork.scala 178:25]
    end else if (w_vn_lvl_0_valid_11 & ~w_vn_lvl_0_valid_10) begin // @[FanNetwork.scala 181:70]
      r_lvl_output_ff_10 <= 32'h0; // @[FanNetwork.scala 183:25]
    end else if (~w_vn_lvl_0_valid_11 & w_vn_lvl_0_valid_10) begin // @[FanNetwork.scala 186:70]
      r_lvl_output_ff_10 <= w_vn_lvl_0_10; // @[FanNetwork.scala 188:25]
    end else begin
      r_lvl_output_ff_10 <= 32'h0; // @[FanNetwork.scala 193:25]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_11 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_11 <= r_lvl_output_ff_79; // @[FanNetwork.scala 803:25]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_12 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_0_valid_13 & w_vn_lvl_0_valid_12) begin // @[FanNetwork.scala 199:63]
      r_lvl_output_ff_12 <= w_vn_lvl_0_12; // @[FanNetwork.scala 201:25]
    end else if (w_vn_lvl_0_valid_13 & ~w_vn_lvl_0_valid_12) begin // @[FanNetwork.scala 204:70]
      r_lvl_output_ff_12 <= 32'h0; // @[FanNetwork.scala 206:25]
    end else if (~w_vn_lvl_0_valid_13 & w_vn_lvl_0_valid_12) begin // @[FanNetwork.scala 209:70]
      r_lvl_output_ff_12 <= w_vn_lvl_0_12; // @[FanNetwork.scala 211:25]
    end else begin
      r_lvl_output_ff_12 <= 32'h0; // @[FanNetwork.scala 216:25]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_13 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_0_valid_13 & w_vn_lvl_0_valid_12) begin // @[FanNetwork.scala 199:63]
      r_lvl_output_ff_13 <= w_vn_lvl_0_13; // @[FanNetwork.scala 200:25]
    end else if (w_vn_lvl_0_valid_13 & ~w_vn_lvl_0_valid_12) begin // @[FanNetwork.scala 204:70]
      r_lvl_output_ff_13 <= w_vn_lvl_0_13; // @[FanNetwork.scala 205:25]
    end else begin
      r_lvl_output_ff_13 <= 32'h0;
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_14 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_0_valid_15 & w_vn_lvl_0_valid_14) begin // @[FanNetwork.scala 222:63]
      r_lvl_output_ff_14 <= w_vn_lvl_0_14; // @[FanNetwork.scala 224:25]
    end else if (w_vn_lvl_0_valid_15 & ~w_vn_lvl_0_valid_14) begin // @[FanNetwork.scala 227:70]
      r_lvl_output_ff_14 <= 32'h0; // @[FanNetwork.scala 229:25]
    end else if (~w_vn_lvl_0_valid_15 & w_vn_lvl_0_valid_14) begin // @[FanNetwork.scala 232:70]
      r_lvl_output_ff_14 <= w_vn_lvl_0_14; // @[FanNetwork.scala 234:25]
    end else begin
      r_lvl_output_ff_14 <= 32'h0; // @[FanNetwork.scala 239:25]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_15 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_0_valid_15 & w_vn_lvl_0_valid_14) begin // @[FanNetwork.scala 222:63]
      r_lvl_output_ff_15 <= w_vn_lvl_0_15; // @[FanNetwork.scala 223:25]
    end else if (w_vn_lvl_0_valid_15 & ~w_vn_lvl_0_valid_14) begin // @[FanNetwork.scala 227:70]
      r_lvl_output_ff_15 <= w_vn_lvl_0_15; // @[FanNetwork.scala 228:25]
    end else begin
      r_lvl_output_ff_15 <= 32'h0;
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_16 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_0_valid_17 & w_vn_lvl_0_valid_16) begin // @[FanNetwork.scala 245:63]
      r_lvl_output_ff_16 <= w_vn_lvl_0_16; // @[FanNetwork.scala 247:25]
    end else if (w_vn_lvl_0_valid_17 & ~w_vn_lvl_0_valid_16) begin // @[FanNetwork.scala 250:70]
      r_lvl_output_ff_16 <= 32'h0; // @[FanNetwork.scala 252:25]
    end else if (~w_vn_lvl_0_valid_17 & w_vn_lvl_0_valid_16) begin // @[FanNetwork.scala 255:70]
      r_lvl_output_ff_16 <= w_vn_lvl_0_16; // @[FanNetwork.scala 257:25]
    end else begin
      r_lvl_output_ff_16 <= 32'h0; // @[FanNetwork.scala 262:25]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_17 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_0_valid_17 & w_vn_lvl_0_valid_16) begin // @[FanNetwork.scala 245:63]
      r_lvl_output_ff_17 <= w_vn_lvl_0_17; // @[FanNetwork.scala 246:25]
    end else if (w_vn_lvl_0_valid_17 & ~w_vn_lvl_0_valid_16) begin // @[FanNetwork.scala 250:70]
      r_lvl_output_ff_17 <= w_vn_lvl_0_17; // @[FanNetwork.scala 251:25]
    end else begin
      r_lvl_output_ff_17 <= 32'h0;
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_18 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_0_valid_19 & w_vn_lvl_0_valid_18) begin // @[FanNetwork.scala 268:63]
      r_lvl_output_ff_18 <= w_vn_lvl_0_18; // @[FanNetwork.scala 270:25]
    end else if (w_vn_lvl_0_valid_19 & ~w_vn_lvl_0_valid_18) begin // @[FanNetwork.scala 273:70]
      r_lvl_output_ff_18 <= 32'h0; // @[FanNetwork.scala 275:25]
    end else if (~w_vn_lvl_0_valid_19 & w_vn_lvl_0_valid_18) begin // @[FanNetwork.scala 278:70]
      r_lvl_output_ff_18 <= w_vn_lvl_0_18; // @[FanNetwork.scala 280:25]
    end else begin
      r_lvl_output_ff_18 <= 32'h0; // @[FanNetwork.scala 285:25]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_19 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_0_valid_19 & w_vn_lvl_0_valid_18) begin // @[FanNetwork.scala 268:63]
      r_lvl_output_ff_19 <= w_vn_lvl_0_19; // @[FanNetwork.scala 269:25]
    end else if (w_vn_lvl_0_valid_19 & ~w_vn_lvl_0_valid_18) begin // @[FanNetwork.scala 273:70]
      r_lvl_output_ff_19 <= w_vn_lvl_0_19; // @[FanNetwork.scala 274:25]
    end else begin
      r_lvl_output_ff_19 <= 32'h0;
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_20 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_0_valid_21 & w_vn_lvl_0_valid_20) begin // @[FanNetwork.scala 291:63]
      r_lvl_output_ff_20 <= w_vn_lvl_0_20; // @[FanNetwork.scala 293:25]
    end else if (w_vn_lvl_0_valid_21 & ~w_vn_lvl_0_valid_20) begin // @[FanNetwork.scala 296:70]
      r_lvl_output_ff_20 <= 32'h0; // @[FanNetwork.scala 298:25]
    end else if (~w_vn_lvl_0_valid_21 & w_vn_lvl_0_valid_20) begin // @[FanNetwork.scala 301:70]
      r_lvl_output_ff_20 <= w_vn_lvl_0_20; // @[FanNetwork.scala 303:25]
    end else begin
      r_lvl_output_ff_20 <= 32'h0; // @[FanNetwork.scala 308:25]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_21 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_0_valid_21 & w_vn_lvl_0_valid_20) begin // @[FanNetwork.scala 291:63]
      r_lvl_output_ff_21 <= w_vn_lvl_0_21; // @[FanNetwork.scala 292:25]
    end else if (w_vn_lvl_0_valid_21 & ~w_vn_lvl_0_valid_20) begin // @[FanNetwork.scala 296:70]
      r_lvl_output_ff_21 <= w_vn_lvl_0_21; // @[FanNetwork.scala 297:25]
    end else begin
      r_lvl_output_ff_21 <= 32'h0;
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_22 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_0_valid_23 & w_vn_lvl_0_valid_22) begin // @[FanNetwork.scala 314:63]
      r_lvl_output_ff_22 <= w_vn_lvl_0_22; // @[FanNetwork.scala 316:25]
    end else if (w_vn_lvl_0_valid_23 & ~w_vn_lvl_0_valid_22) begin // @[FanNetwork.scala 319:70]
      r_lvl_output_ff_22 <= 32'h0; // @[FanNetwork.scala 321:25]
    end else if (~w_vn_lvl_0_valid_23 & w_vn_lvl_0_valid_22) begin // @[FanNetwork.scala 324:70]
      r_lvl_output_ff_22 <= w_vn_lvl_0_22; // @[FanNetwork.scala 326:25]
    end else begin
      r_lvl_output_ff_22 <= 32'h0; // @[FanNetwork.scala 331:25]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_23 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_0_valid_23 & w_vn_lvl_0_valid_22) begin // @[FanNetwork.scala 314:63]
      r_lvl_output_ff_23 <= w_vn_lvl_0_23; // @[FanNetwork.scala 315:25]
    end else if (w_vn_lvl_0_valid_23 & ~w_vn_lvl_0_valid_22) begin // @[FanNetwork.scala 319:70]
      r_lvl_output_ff_23 <= w_vn_lvl_0_23; // @[FanNetwork.scala 320:25]
    end else begin
      r_lvl_output_ff_23 <= 32'h0;
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_24 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_0_valid_25 & w_vn_lvl_0_valid_24) begin // @[FanNetwork.scala 337:63]
      r_lvl_output_ff_24 <= w_vn_lvl_0_24; // @[FanNetwork.scala 339:25]
    end else if (w_vn_lvl_0_valid_25 & ~w_vn_lvl_0_valid_24) begin // @[FanNetwork.scala 342:70]
      r_lvl_output_ff_24 <= 32'h0; // @[FanNetwork.scala 344:25]
    end else if (~w_vn_lvl_0_valid_25 & w_vn_lvl_0_valid_24) begin // @[FanNetwork.scala 347:70]
      r_lvl_output_ff_24 <= w_vn_lvl_0_24; // @[FanNetwork.scala 349:25]
    end else begin
      r_lvl_output_ff_24 <= 32'h0; // @[FanNetwork.scala 354:25]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_25 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_0_valid_25 & w_vn_lvl_0_valid_24) begin // @[FanNetwork.scala 337:63]
      r_lvl_output_ff_25 <= w_vn_lvl_0_25; // @[FanNetwork.scala 338:25]
    end else if (w_vn_lvl_0_valid_25 & ~w_vn_lvl_0_valid_24) begin // @[FanNetwork.scala 342:70]
      r_lvl_output_ff_25 <= w_vn_lvl_0_25; // @[FanNetwork.scala 343:25]
    end else begin
      r_lvl_output_ff_25 <= 32'h0;
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_26 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_0_valid_27 & w_vn_lvl_0_valid_26) begin // @[FanNetwork.scala 360:63]
      r_lvl_output_ff_26 <= w_vn_lvl_0_26; // @[FanNetwork.scala 362:25]
    end else if (w_vn_lvl_0_valid_27 & ~w_vn_lvl_0_valid_26) begin // @[FanNetwork.scala 365:70]
      r_lvl_output_ff_26 <= 32'h0; // @[FanNetwork.scala 367:25]
    end else if (~w_vn_lvl_0_valid_27 & w_vn_lvl_0_valid_26) begin // @[FanNetwork.scala 370:70]
      r_lvl_output_ff_26 <= w_vn_lvl_0_26; // @[FanNetwork.scala 372:25]
    end else begin
      r_lvl_output_ff_26 <= 32'h0; // @[FanNetwork.scala 377:25]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_27 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_0_valid_27 & w_vn_lvl_0_valid_26) begin // @[FanNetwork.scala 360:63]
      r_lvl_output_ff_27 <= w_vn_lvl_0_27; // @[FanNetwork.scala 361:25]
    end else if (w_vn_lvl_0_valid_27 & ~w_vn_lvl_0_valid_26) begin // @[FanNetwork.scala 365:70]
      r_lvl_output_ff_27 <= w_vn_lvl_0_27; // @[FanNetwork.scala 366:25]
    end else begin
      r_lvl_output_ff_27 <= 32'h0;
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_28 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_0_valid_29 & w_vn_lvl_0_valid_28) begin // @[FanNetwork.scala 383:63]
      r_lvl_output_ff_28 <= w_vn_lvl_0_28; // @[FanNetwork.scala 385:25]
    end else if (w_vn_lvl_0_valid_29 & ~w_vn_lvl_0_valid_28) begin // @[FanNetwork.scala 388:70]
      r_lvl_output_ff_28 <= 32'h0; // @[FanNetwork.scala 390:25]
    end else if (~w_vn_lvl_0_valid_29 & w_vn_lvl_0_valid_28) begin // @[FanNetwork.scala 393:70]
      r_lvl_output_ff_28 <= w_vn_lvl_0_28; // @[FanNetwork.scala 395:25]
    end else begin
      r_lvl_output_ff_28 <= 32'h0; // @[FanNetwork.scala 400:25]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_29 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_0_valid_29 & w_vn_lvl_0_valid_28) begin // @[FanNetwork.scala 383:63]
      r_lvl_output_ff_29 <= w_vn_lvl_0_29; // @[FanNetwork.scala 384:25]
    end else if (w_vn_lvl_0_valid_29 & ~w_vn_lvl_0_valid_28) begin // @[FanNetwork.scala 388:70]
      r_lvl_output_ff_29 <= w_vn_lvl_0_29; // @[FanNetwork.scala 389:25]
    end else begin
      r_lvl_output_ff_29 <= 32'h0;
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_30 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_0_valid_31 & w_vn_lvl_0_valid_30) begin // @[FanNetwork.scala 406:62]
      r_lvl_output_ff_30 <= w_vn_lvl_0_30; // @[FanNetwork.scala 408:25]
    end else if (w_vn_lvl_0_valid_31 & ~w_vn_lvl_0_valid_30) begin // @[FanNetwork.scala 411:69]
      r_lvl_output_ff_30 <= 32'h0; // @[FanNetwork.scala 413:25]
    end else if (~w_vn_lvl_0_valid_31 & w_vn_lvl_0_valid_30) begin // @[FanNetwork.scala 416:69]
      r_lvl_output_ff_30 <= w_vn_lvl_0_30; // @[FanNetwork.scala 418:25]
    end else begin
      r_lvl_output_ff_30 <= 32'h0; // @[FanNetwork.scala 423:25]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_31 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_0_valid_31 & w_vn_lvl_0_valid_30) begin // @[FanNetwork.scala 406:62]
      r_lvl_output_ff_31 <= w_vn_lvl_0_31; // @[FanNetwork.scala 407:25]
    end else if (w_vn_lvl_0_valid_31 & ~w_vn_lvl_0_valid_30) begin // @[FanNetwork.scala 411:69]
      r_lvl_output_ff_31 <= w_vn_lvl_0_31; // @[FanNetwork.scala 412:25]
    end else begin
      r_lvl_output_ff_31 <= 32'h0;
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_32 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_32 <= r_lvl_output_ff_0; // @[FanNetwork.scala 431:25]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_33 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_1_valid_0) begin // @[FanNetwork.scala 434:34]
      r_lvl_output_ff_33 <= w_vn_lvl_1_0; // @[FanNetwork.scala 435:29]
    end else begin
      r_lvl_output_ff_33 <= r_lvl_output_ff_1; // @[FanNetwork.scala 438:29]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_34 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_1_valid_1) begin // @[FanNetwork.scala 442:34]
      r_lvl_output_ff_34 <= w_vn_lvl_1_1; // @[FanNetwork.scala 443:29]
    end else begin
      r_lvl_output_ff_34 <= r_lvl_output_ff_2; // @[FanNetwork.scala 446:29]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_35 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_35 <= r_lvl_output_ff_3; // @[FanNetwork.scala 450:25]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_36 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_36 <= r_lvl_output_ff_4; // @[FanNetwork.scala 453:27]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_37 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_1_valid_2) begin // @[FanNetwork.scala 456:34]
      r_lvl_output_ff_37 <= w_vn_lvl_1_2; // @[FanNetwork.scala 457:29]
    end else begin
      r_lvl_output_ff_37 <= r_lvl_output_ff_5; // @[FanNetwork.scala 460:29]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_38 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_1_valid_3) begin // @[FanNetwork.scala 464:34]
      r_lvl_output_ff_38 <= w_vn_lvl_1_3; // @[FanNetwork.scala 465:29]
    end else begin
      r_lvl_output_ff_38 <= r_lvl_output_ff_6; // @[FanNetwork.scala 468:29]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_39 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_39 <= r_lvl_output_ff_7; // @[FanNetwork.scala 474:25]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_40 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_40 <= r_lvl_output_ff_8; // @[FanNetwork.scala 477:25]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_41 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_1_valid_4) begin // @[FanNetwork.scala 480:34]
      r_lvl_output_ff_41 <= w_vn_lvl_1_4; // @[FanNetwork.scala 481:29]
    end else begin
      r_lvl_output_ff_41 <= r_lvl_output_ff_9; // @[FanNetwork.scala 484:29]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_42 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_1_valid_5) begin // @[FanNetwork.scala 487:34]
      r_lvl_output_ff_42 <= w_vn_lvl_1_5; // @[FanNetwork.scala 488:29]
    end else begin
      r_lvl_output_ff_42 <= r_lvl_output_ff_10; // @[FanNetwork.scala 491:29]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_43 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_43 <= r_lvl_output_ff_11; // @[FanNetwork.scala 495:25]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_44 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_44 <= r_lvl_output_ff_12; // @[FanNetwork.scala 498:25]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_45 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_1_valid_6) begin // @[FanNetwork.scala 501:34]
      r_lvl_output_ff_45 <= w_vn_lvl_1_6; // @[FanNetwork.scala 502:29]
    end else begin
      r_lvl_output_ff_45 <= r_lvl_output_ff_13; // @[FanNetwork.scala 505:29]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_46 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_1_valid_7) begin // @[FanNetwork.scala 509:34]
      r_lvl_output_ff_46 <= w_vn_lvl_1_7; // @[FanNetwork.scala 510:29]
    end else begin
      r_lvl_output_ff_46 <= r_lvl_output_ff_14; // @[FanNetwork.scala 513:29]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_47 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_47 <= r_lvl_output_ff_15; // @[FanNetwork.scala 516:25]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_48 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_48 <= r_lvl_output_ff_16; // @[FanNetwork.scala 519:25]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_49 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_1_valid_8) begin // @[FanNetwork.scala 522:34]
      r_lvl_output_ff_49 <= w_vn_lvl_1_8; // @[FanNetwork.scala 523:29]
    end else begin
      r_lvl_output_ff_49 <= r_lvl_output_ff_17; // @[FanNetwork.scala 526:29]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_50 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_1_valid_9) begin // @[FanNetwork.scala 530:34]
      r_lvl_output_ff_50 <= w_vn_lvl_1_9; // @[FanNetwork.scala 531:29]
    end else begin
      r_lvl_output_ff_50 <= r_lvl_output_ff_18; // @[FanNetwork.scala 534:29]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_51 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_51 <= r_lvl_output_ff_19; // @[FanNetwork.scala 540:25]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_52 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_52 <= r_lvl_output_ff_20; // @[FanNetwork.scala 543:25]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_53 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_1_valid_10) begin // @[FanNetwork.scala 546:35]
      r_lvl_output_ff_53 <= w_vn_lvl_1_10; // @[FanNetwork.scala 547:29]
    end else begin
      r_lvl_output_ff_53 <= r_lvl_output_ff_21; // @[FanNetwork.scala 550:29]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_54 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_1_valid_11) begin // @[FanNetwork.scala 554:35]
      r_lvl_output_ff_54 <= w_vn_lvl_1_11; // @[FanNetwork.scala 555:29]
    end else begin
      r_lvl_output_ff_54 <= r_lvl_output_ff_22; // @[FanNetwork.scala 558:29]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_55 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_55 <= r_lvl_output_ff_23; // @[FanNetwork.scala 562:25]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_56 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_56 <= r_lvl_output_ff_24; // @[FanNetwork.scala 565:25]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_57 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_1_valid_12) begin // @[FanNetwork.scala 568:35]
      r_lvl_output_ff_57 <= w_vn_lvl_1_12; // @[FanNetwork.scala 569:29]
    end else begin
      r_lvl_output_ff_57 <= r_lvl_output_ff_25; // @[FanNetwork.scala 572:29]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_58 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_1_valid_13) begin // @[FanNetwork.scala 576:35]
      r_lvl_output_ff_58 <= w_vn_lvl_1_13; // @[FanNetwork.scala 577:29]
    end else begin
      r_lvl_output_ff_58 <= r_lvl_output_ff_26; // @[FanNetwork.scala 580:29]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_59 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_59 <= r_lvl_output_ff_27; // @[FanNetwork.scala 584:25]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_60 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_60 <= r_lvl_output_ff_28; // @[FanNetwork.scala 587:25]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_61 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_1_valid_14) begin // @[FanNetwork.scala 590:43]
      r_lvl_output_ff_61 <= w_vn_lvl_1_14; // @[FanNetwork.scala 591:29]
    end else begin
      r_lvl_output_ff_61 <= r_lvl_output_ff_29; // @[FanNetwork.scala 594:29]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_62 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_1_valid_15) begin // @[FanNetwork.scala 598:43]
      r_lvl_output_ff_62 <= w_vn_lvl_1_15; // @[FanNetwork.scala 599:29]
    end else begin
      r_lvl_output_ff_62 <= r_lvl_output_ff_30; // @[FanNetwork.scala 602:29]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_63 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_63 <= r_lvl_output_ff_31; // @[FanNetwork.scala 606:25]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_64 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_64 <= r_lvl_output_ff_32; // @[FanNetwork.scala 610:26]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_65 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_65 <= r_lvl_output_ff_33; // @[FanNetwork.scala 613:25]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_66 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_66 <= r_lvl_output_ff_34; // @[FanNetwork.scala 616:25]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_67 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_2_valid_0) begin // @[FanNetwork.scala 619:43]
      r_lvl_output_ff_67 <= w_vn_lvl_2_0; // @[FanNetwork.scala 620:29]
    end else begin
      r_lvl_output_ff_67 <= r_lvl_output_ff_35; // @[FanNetwork.scala 623:33]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_68 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_2_valid_1) begin // @[FanNetwork.scala 627:43]
      r_lvl_output_ff_68 <= w_vn_lvl_2_1; // @[FanNetwork.scala 628:29]
    end else begin
      r_lvl_output_ff_68 <= r_lvl_output_ff_36; // @[FanNetwork.scala 631:29]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_69 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_69 <= r_lvl_output_ff_37; // @[FanNetwork.scala 635:25]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_70 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_70 <= r_lvl_output_ff_38; // @[FanNetwork.scala 638:25]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_71 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_71 <= r_lvl_output_ff_39; // @[FanNetwork.scala 641:25]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_72 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_72 <= r_lvl_output_ff_40; // @[FanNetwork.scala 644:25]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_73 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_73 <= r_lvl_output_ff_41; // @[FanNetwork.scala 647:25]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_74 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_74 <= r_lvl_output_ff_42; // @[FanNetwork.scala 650:25]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_75 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_2_valid_2) begin // @[FanNetwork.scala 653:43]
      r_lvl_output_ff_75 <= w_vn_lvl_2_2; // @[FanNetwork.scala 654:29]
    end else begin
      r_lvl_output_ff_75 <= r_lvl_output_ff_43; // @[FanNetwork.scala 657:29]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_76 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_2_valid_3) begin // @[FanNetwork.scala 661:43]
      r_lvl_output_ff_76 <= w_vn_lvl_2_3; // @[FanNetwork.scala 662:29]
    end else begin
      r_lvl_output_ff_76 <= r_lvl_output_ff_44; // @[FanNetwork.scala 665:29]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_77 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_77 <= r_lvl_output_ff_45; // @[FanNetwork.scala 669:25]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_78 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_78 <= r_lvl_output_ff_46; // @[FanNetwork.scala 672:25]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_79 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_79 <= r_lvl_output_ff_47; // @[FanNetwork.scala 675:25]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_80 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_80 <= r_lvl_output_ff_48; // @[FanNetwork.scala 678:25]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_81 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_81 <= r_lvl_output_ff_49; // @[FanNetwork.scala 681:25]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_82 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_82 <= r_lvl_output_ff_50; // @[FanNetwork.scala 684:25]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_83 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_2_valid_4) begin // @[FanNetwork.scala 687:43]
      r_lvl_output_ff_83 <= w_vn_lvl_2_4; // @[FanNetwork.scala 688:29]
    end else begin
      r_lvl_output_ff_83 <= r_lvl_output_ff_51; // @[FanNetwork.scala 691:29]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_84 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_2_valid_5) begin // @[FanNetwork.scala 695:40]
      r_lvl_output_ff_84 <= w_vn_lvl_2_5; // @[FanNetwork.scala 696:29]
    end else begin
      r_lvl_output_ff_84 <= r_lvl_output_ff_52; // @[FanNetwork.scala 699:29]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_85 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_85 <= r_lvl_output_ff_53; // @[FanNetwork.scala 703:25]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_86 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_86 <= r_lvl_output_ff_54; // @[FanNetwork.scala 706:25]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_87 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_87 <= r_lvl_output_ff_55; // @[FanNetwork.scala 709:25]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_88 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_88 <= r_lvl_output_ff_56; // @[FanNetwork.scala 712:25]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_89 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_89 <= r_lvl_output_ff_57; // @[FanNetwork.scala 715:25]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_90 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_90 <= r_lvl_output_ff_58; // @[FanNetwork.scala 718:25]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_91 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_2_valid_6) begin // @[FanNetwork.scala 721:40]
      r_lvl_output_ff_91 <= w_vn_lvl_2_6; // @[FanNetwork.scala 722:29]
    end else begin
      r_lvl_output_ff_91 <= r_lvl_output_ff_59; // @[FanNetwork.scala 725:29]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_92 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_2_valid_7) begin // @[FanNetwork.scala 729:40]
      r_lvl_output_ff_92 <= w_vn_lvl_2_7; // @[FanNetwork.scala 730:29]
    end else begin
      r_lvl_output_ff_92 <= r_lvl_output_ff_60; // @[FanNetwork.scala 733:29]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_93 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_93 <= r_lvl_output_ff_61; // @[FanNetwork.scala 737:25]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_94 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_94 <= r_lvl_output_ff_62; // @[FanNetwork.scala 740:25]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_95 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_95 <= r_lvl_output_ff_63; // @[FanNetwork.scala 743:25]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_96 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_96 <= r_lvl_output_ff_64; // @[FanNetwork.scala 748:25]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_97 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_97 <= r_lvl_output_ff_65; // @[FanNetwork.scala 751:25]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_98 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_98 <= r_lvl_output_ff_66; // @[FanNetwork.scala 754:25]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_99 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_99 <= r_lvl_output_ff_67; // @[FanNetwork.scala 757:25]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_100 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_100 <= r_lvl_output_ff_68; // @[FanNetwork.scala 760:26]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_101 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_101 <= r_lvl_output_ff_69; // @[FanNetwork.scala 763:26]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_102 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_102 <= r_lvl_output_ff_70; // @[FanNetwork.scala 766:26]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_103 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_3_valid_0) begin // @[FanNetwork.scala 769:40]
      r_lvl_output_ff_103 <= w_vn_lvl_3_0; // @[FanNetwork.scala 770:28]
    end else begin
      r_lvl_output_ff_103 <= r_lvl_output_ff_71; // @[FanNetwork.scala 773:28]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_104 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_3_valid_1) begin // @[FanNetwork.scala 777:40]
      r_lvl_output_ff_104 <= w_vn_lvl_3_1; // @[FanNetwork.scala 778:28]
    end else begin
      r_lvl_output_ff_104 <= r_lvl_output_ff_72; // @[FanNetwork.scala 781:28]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_105 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_105 <= r_lvl_output_ff_73; // @[FanNetwork.scala 785:26]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_106 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_106 <= r_lvl_output_ff_74; // @[FanNetwork.scala 788:26]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_107 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_107 <= r_lvl_output_ff_75; // @[FanNetwork.scala 791:26]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_108 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_108 <= r_lvl_output_ff_76; // @[FanNetwork.scala 794:26]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_109 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_109 <= r_lvl_output_ff_77; // @[FanNetwork.scala 797:26]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_110 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_110 <= r_lvl_output_ff_78; // @[FanNetwork.scala 800:26]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_112 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_112 <= r_lvl_output_ff_80; // @[FanNetwork.scala 806:26]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_113 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_113 <= r_lvl_output_ff_81; // @[FanNetwork.scala 809:26]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_114 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_114 <= r_lvl_output_ff_82; // @[FanNetwork.scala 812:26]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_115 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_115 <= r_lvl_output_ff_83; // @[FanNetwork.scala 815:26]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_116 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_116 <= r_lvl_output_ff_84; // @[FanNetwork.scala 818:26]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_117 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_117 <= r_lvl_output_ff_85; // @[FanNetwork.scala 821:26]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_118 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_118 <= r_lvl_output_ff_86; // @[FanNetwork.scala 824:26]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_119 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_3_valid_2) begin // @[FanNetwork.scala 827:40]
      r_lvl_output_ff_119 <= w_vn_lvl_3_2; // @[FanNetwork.scala 828:30]
    end else begin
      r_lvl_output_ff_119 <= r_lvl_output_ff_87; // @[FanNetwork.scala 831:30]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_120 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_3_valid_3) begin // @[FanNetwork.scala 835:41]
      r_lvl_output_ff_120 <= w_vn_lvl_3_3; // @[FanNetwork.scala 836:30]
    end else begin
      r_lvl_output_ff_120 <= r_lvl_output_ff_88; // @[FanNetwork.scala 839:30]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_121 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_121 <= r_lvl_output_ff_89; // @[FanNetwork.scala 843:26]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_122 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_122 <= r_lvl_output_ff_90; // @[FanNetwork.scala 846:26]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_123 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_123 <= r_lvl_output_ff_91; // @[FanNetwork.scala 849:26]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_124 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_124 <= r_lvl_output_ff_92; // @[FanNetwork.scala 852:26]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_125 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_125 <= r_lvl_output_ff_93; // @[FanNetwork.scala 855:26]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_126 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_126 <= r_lvl_output_ff_94; // @[FanNetwork.scala 858:26]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_127 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_127 <= r_lvl_output_ff_95; // @[FanNetwork.scala 861:26]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_128 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_128 <= r_lvl_output_ff_96; // @[FanNetwork.scala 865:26]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_129 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_129 <= r_lvl_output_ff_97; // @[FanNetwork.scala 868:26]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_130 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_130 <= r_lvl_output_ff_98; // @[FanNetwork.scala 871:26]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_131 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_131 <= r_lvl_output_ff_99; // @[FanNetwork.scala 874:26]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_132 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_132 <= r_lvl_output_ff_100; // @[FanNetwork.scala 877:26]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_133 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_133 <= r_lvl_output_ff_101; // @[FanNetwork.scala 880:26]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_134 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_134 <= r_lvl_output_ff_102; // @[FanNetwork.scala 883:26]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_135 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_135 <= r_lvl_output_ff_103; // @[FanNetwork.scala 886:26]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_136 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_136 <= r_lvl_output_ff_104; // @[FanNetwork.scala 889:26]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_137 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_137 <= r_lvl_output_ff_105; // @[FanNetwork.scala 892:26]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_138 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_138 <= r_lvl_output_ff_106; // @[FanNetwork.scala 895:26]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_139 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_139 <= r_lvl_output_ff_107; // @[FanNetwork.scala 898:26]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_140 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_140 <= r_lvl_output_ff_108; // @[FanNetwork.scala 901:26]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_141 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_141 <= r_lvl_output_ff_109; // @[FanNetwork.scala 904:26]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_142 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_142 <= r_lvl_output_ff_110; // @[FanNetwork.scala 907:26]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_143 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_4_valid_0) begin // @[FanNetwork.scala 910:40]
      r_lvl_output_ff_143 <= w_vn_lvl_4_0; // @[FanNetwork.scala 911:30]
    end else begin
      r_lvl_output_ff_143 <= 32'h0; // @[FanNetwork.scala 914:30]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_144 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else if (w_vn_lvl_4_valid_1) begin // @[FanNetwork.scala 918:40]
      r_lvl_output_ff_144 <= w_vn_lvl_4_1; // @[FanNetwork.scala 919:30]
    end else begin
      r_lvl_output_ff_144 <= r_lvl_output_ff_112; // @[FanNetwork.scala 922:30]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_145 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_145 <= r_lvl_output_ff_113; // @[FanNetwork.scala 926:26]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_146 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_146 <= r_lvl_output_ff_114; // @[FanNetwork.scala 929:26]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_147 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_147 <= r_lvl_output_ff_115; // @[FanNetwork.scala 932:26]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_148 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_148 <= r_lvl_output_ff_116; // @[FanNetwork.scala 935:26]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_149 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_149 <= r_lvl_output_ff_117; // @[FanNetwork.scala 938:26]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_150 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_150 <= r_lvl_output_ff_118; // @[FanNetwork.scala 941:26]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_151 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_151 <= r_lvl_output_ff_119; // @[FanNetwork.scala 944:26]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_152 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_152 <= r_lvl_output_ff_120; // @[FanNetwork.scala 947:26]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_153 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_153 <= r_lvl_output_ff_121; // @[FanNetwork.scala 950:26]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_154 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_154 <= r_lvl_output_ff_122; // @[FanNetwork.scala 953:26]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_155 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_155 <= r_lvl_output_ff_123; // @[FanNetwork.scala 956:26]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_156 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_156 <= r_lvl_output_ff_124; // @[FanNetwork.scala 959:26]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_157 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_157 <= r_lvl_output_ff_125; // @[FanNetwork.scala 962:26]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_158 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_158 <= r_lvl_output_ff_126; // @[FanNetwork.scala 965:26]
    end
    if (reset) begin // @[FanNetwork.scala 45:34]
      r_lvl_output_ff_159 <= 32'h0; // @[FanNetwork.scala 45:34]
    end else begin
      r_lvl_output_ff_159 <= r_lvl_output_ff_127; // @[FanNetwork.scala 968:26]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_0 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_0 <= _GEN_10;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_1 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_1 <= _GEN_9;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_2 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_2 <= _GEN_21;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_3 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_3 <= _GEN_20;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_4 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_4 <= _GEN_32;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_5 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_5 <= _GEN_31;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_6 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_6 <= _GEN_43;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_7 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_7 <= _GEN_42;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_8 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_8 <= _GEN_54;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_9 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_9 <= _GEN_53;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_10 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_10 <= _GEN_65;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_11 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_11 <= _GEN_64;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_12 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_12 <= _GEN_76;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_13 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_13 <= _GEN_75;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_14 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_14 <= _GEN_87;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_15 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_15 <= _GEN_86;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_16 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_16 <= _GEN_98;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_17 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_17 <= _GEN_97;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_18 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_18 <= _GEN_109;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_19 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_19 <= _GEN_108;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_20 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_20 <= _GEN_120;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_21 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_21 <= _GEN_119;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_22 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_22 <= _GEN_131;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_23 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_23 <= _GEN_130;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_24 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_24 <= _GEN_142;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_25 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_25 <= _GEN_141;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_26 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_26 <= _GEN_153;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_27 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_27 <= _GEN_152;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_28 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_28 <= _GEN_164;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_29 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_29 <= _GEN_163;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_30 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_30 <= _GEN_175;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_31 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_31 <= _GEN_174;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_32 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_32 <= r_lvl_output_ff_valid_0; // @[FanNetwork.scala 432:31]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_33 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_33 <= _GEN_177;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_34 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_34 <= _GEN_179;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_35 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_35 <= r_lvl_output_ff_valid_3; // @[FanNetwork.scala 451:31]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_36 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_36 <= r_lvl_output_ff_valid_4; // @[FanNetwork.scala 454:31]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_37 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_37 <= _GEN_181;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_38 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_38 <= _GEN_183;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_39 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_39 <= r_lvl_output_ff_valid_7; // @[FanNetwork.scala 475:31]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_40 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_40 <= r_lvl_output_ff_valid_8; // @[FanNetwork.scala 478:31]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_41 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_41 <= _GEN_185;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_42 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_42 <= _GEN_187;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_43 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_43 <= r_lvl_output_ff_valid_11; // @[FanNetwork.scala 496:31]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_44 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_44 <= r_lvl_output_ff_valid_12; // @[FanNetwork.scala 499:31]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_45 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_45 <= _GEN_189;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_46 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_46 <= _GEN_191;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_47 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_47 <= r_lvl_output_ff_valid_15; // @[FanNetwork.scala 517:31]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_48 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_48 <= r_lvl_output_ff_valid_16; // @[FanNetwork.scala 520:31]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_49 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_49 <= _GEN_193;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_50 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_50 <= _GEN_195;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_51 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_51 <= r_lvl_output_ff_valid_19; // @[FanNetwork.scala 541:31]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_52 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_52 <= r_lvl_output_ff_valid_20; // @[FanNetwork.scala 544:31]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_53 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_53 <= _GEN_197;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_54 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_54 <= _GEN_199;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_55 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_55 <= r_lvl_output_ff_valid_23; // @[FanNetwork.scala 563:31]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_56 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_56 <= r_lvl_output_ff_valid_24; // @[FanNetwork.scala 566:31]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_57 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_57 <= _GEN_201;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_58 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_58 <= _GEN_203;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_59 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_59 <= r_lvl_output_ff_valid_27; // @[FanNetwork.scala 585:31]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_60 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_60 <= r_lvl_output_ff_valid_28; // @[FanNetwork.scala 588:31]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_61 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_61 <= _GEN_205;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_62 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_62 <= _GEN_207;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_63 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_63 <= r_lvl_output_ff_valid_31; // @[FanNetwork.scala 607:31]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_64 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_64 <= r_lvl_output_ff_valid_32; // @[FanNetwork.scala 611:31]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_65 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_65 <= r_lvl_output_ff_valid_33; // @[FanNetwork.scala 614:31]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_66 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_66 <= r_lvl_output_ff_valid_34; // @[FanNetwork.scala 617:31]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_67 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_67 <= _GEN_209;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_68 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_68 <= _GEN_211;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_69 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_69 <= r_lvl_output_ff_valid_37; // @[FanNetwork.scala 636:31]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_70 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_70 <= r_lvl_output_ff_valid_38; // @[FanNetwork.scala 639:31]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_71 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_71 <= r_lvl_output_ff_valid_39; // @[FanNetwork.scala 642:31]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_72 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_72 <= r_lvl_output_ff_valid_40; // @[FanNetwork.scala 645:31]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_73 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_73 <= r_lvl_output_ff_valid_41; // @[FanNetwork.scala 648:31]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_74 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_74 <= r_lvl_output_ff_valid_42; // @[FanNetwork.scala 651:31]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_75 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_75 <= _GEN_213;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_76 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_76 <= _GEN_215;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_77 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_77 <= r_lvl_output_ff_valid_45; // @[FanNetwork.scala 670:31]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_78 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_78 <= r_lvl_output_ff_valid_46; // @[FanNetwork.scala 673:31]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_79 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_79 <= r_lvl_output_ff_valid_47; // @[FanNetwork.scala 676:31]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_80 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_80 <= r_lvl_output_ff_valid_48; // @[FanNetwork.scala 679:31]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_81 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_81 <= r_lvl_output_ff_valid_49; // @[FanNetwork.scala 682:31]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_82 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_82 <= r_lvl_output_ff_valid_50; // @[FanNetwork.scala 685:31]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_83 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_83 <= _GEN_217;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_84 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_84 <= _GEN_219;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_85 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_85 <= r_lvl_output_ff_valid_53; // @[FanNetwork.scala 704:31]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_86 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_86 <= r_lvl_output_ff_valid_54; // @[FanNetwork.scala 707:31]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_87 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_87 <= r_lvl_output_ff_valid_55; // @[FanNetwork.scala 710:31]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_88 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_88 <= r_lvl_output_ff_valid_56; // @[FanNetwork.scala 713:31]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_89 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_89 <= r_lvl_output_ff_valid_57; // @[FanNetwork.scala 716:31]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_90 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_90 <= r_lvl_output_ff_valid_58; // @[FanNetwork.scala 719:31]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_91 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_91 <= _GEN_221;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_92 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_92 <= _GEN_223;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_93 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_93 <= r_lvl_output_ff_valid_61; // @[FanNetwork.scala 738:31]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_94 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_94 <= r_lvl_output_ff_valid_62; // @[FanNetwork.scala 741:31]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_95 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_95 <= r_lvl_output_ff_valid_63; // @[FanNetwork.scala 744:31]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_96 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_96 <= r_lvl_output_ff_valid_64; // @[FanNetwork.scala 749:31]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_97 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_97 <= r_lvl_output_ff_valid_65; // @[FanNetwork.scala 752:31]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_98 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_98 <= r_lvl_output_ff_valid_66; // @[FanNetwork.scala 755:31]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_99 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_99 <= r_lvl_output_ff_valid_67; // @[FanNetwork.scala 758:31]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_100 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_100 <= r_lvl_output_ff_valid_68; // @[FanNetwork.scala 761:32]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_101 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_101 <= r_lvl_output_ff_valid_69; // @[FanNetwork.scala 764:32]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_102 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_102 <= r_lvl_output_ff_valid_70; // @[FanNetwork.scala 767:32]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_103 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_103 <= _GEN_225;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_104 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_104 <= _GEN_227;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_105 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_105 <= r_lvl_output_ff_valid_73; // @[FanNetwork.scala 786:32]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_106 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_106 <= r_lvl_output_ff_valid_74; // @[FanNetwork.scala 789:32]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_107 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_107 <= r_lvl_output_ff_valid_75; // @[FanNetwork.scala 792:32]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_108 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_108 <= r_lvl_output_ff_valid_76; // @[FanNetwork.scala 795:32]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_109 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_109 <= r_lvl_output_ff_valid_77; // @[FanNetwork.scala 798:32]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_110 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_110 <= r_lvl_output_ff_valid_78; // @[FanNetwork.scala 801:32]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_111 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_111 <= r_lvl_output_ff_valid_79; // @[FanNetwork.scala 804:32]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_112 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_112 <= r_lvl_output_ff_valid_80; // @[FanNetwork.scala 807:32]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_113 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_113 <= r_lvl_output_ff_valid_81; // @[FanNetwork.scala 810:32]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_114 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_114 <= r_lvl_output_ff_valid_82; // @[FanNetwork.scala 813:32]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_115 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_115 <= r_lvl_output_ff_valid_83; // @[FanNetwork.scala 816:32]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_116 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_116 <= r_lvl_output_ff_valid_84; // @[FanNetwork.scala 819:32]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_117 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_117 <= r_lvl_output_ff_valid_85; // @[FanNetwork.scala 822:32]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_118 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_118 <= r_lvl_output_ff_valid_86; // @[FanNetwork.scala 825:32]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_119 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_119 <= _GEN_229;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_120 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_120 <= _GEN_231;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_121 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_121 <= r_lvl_output_ff_valid_89; // @[FanNetwork.scala 844:32]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_122 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_122 <= r_lvl_output_ff_valid_90; // @[FanNetwork.scala 847:32]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_123 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_123 <= r_lvl_output_ff_valid_91; // @[FanNetwork.scala 850:32]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_124 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_124 <= r_lvl_output_ff_valid_92; // @[FanNetwork.scala 853:32]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_125 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_125 <= r_lvl_output_ff_valid_93; // @[FanNetwork.scala 856:32]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_126 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_126 <= r_lvl_output_ff_valid_94; // @[FanNetwork.scala 859:32]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_127 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_127 <= r_lvl_output_ff_valid_95; // @[FanNetwork.scala 862:32]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_128 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_128 <= r_lvl_output_ff_valid_96; // @[FanNetwork.scala 866:32]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_129 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_129 <= r_lvl_output_ff_valid_97; // @[FanNetwork.scala 869:32]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_130 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_130 <= r_lvl_output_ff_valid_98; // @[FanNetwork.scala 872:32]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_131 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_131 <= r_lvl_output_ff_valid_99; // @[FanNetwork.scala 875:32]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_132 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_132 <= r_lvl_output_ff_valid_100; // @[FanNetwork.scala 878:32]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_133 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_133 <= r_lvl_output_ff_valid_101; // @[FanNetwork.scala 881:32]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_134 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_134 <= r_lvl_output_ff_valid_102; // @[FanNetwork.scala 884:32]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_135 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_135 <= r_lvl_output_ff_valid_103; // @[FanNetwork.scala 887:32]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_136 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_136 <= r_lvl_output_ff_valid_104; // @[FanNetwork.scala 890:32]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_137 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_137 <= r_lvl_output_ff_valid_105; // @[FanNetwork.scala 893:32]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_138 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_138 <= r_lvl_output_ff_valid_106; // @[FanNetwork.scala 896:32]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_139 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_139 <= r_lvl_output_ff_valid_107; // @[FanNetwork.scala 899:32]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_140 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_140 <= r_lvl_output_ff_valid_108; // @[FanNetwork.scala 902:32]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_141 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_141 <= r_lvl_output_ff_valid_109; // @[FanNetwork.scala 905:32]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_142 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_142 <= r_lvl_output_ff_valid_110; // @[FanNetwork.scala 908:32]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_143 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_143 <= _GEN_233;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_144 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_144 <= _GEN_235;
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_145 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_145 <= r_lvl_output_ff_valid_113; // @[FanNetwork.scala 927:32]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_146 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_146 <= r_lvl_output_ff_valid_114; // @[FanNetwork.scala 930:32]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_147 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_147 <= r_lvl_output_ff_valid_115; // @[FanNetwork.scala 933:32]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_148 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_148 <= r_lvl_output_ff_valid_116; // @[FanNetwork.scala 936:32]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_149 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_149 <= r_lvl_output_ff_valid_117; // @[FanNetwork.scala 939:32]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_150 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_150 <= r_lvl_output_ff_valid_118; // @[FanNetwork.scala 942:32]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_151 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_151 <= r_lvl_output_ff_valid_119; // @[FanNetwork.scala 945:32]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_152 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_152 <= r_lvl_output_ff_valid_120; // @[FanNetwork.scala 948:32]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_153 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_153 <= r_lvl_output_ff_valid_121; // @[FanNetwork.scala 951:32]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_154 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_154 <= r_lvl_output_ff_valid_122; // @[FanNetwork.scala 954:32]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_155 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_155 <= r_lvl_output_ff_valid_123; // @[FanNetwork.scala 957:32]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_156 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_156 <= r_lvl_output_ff_valid_124; // @[FanNetwork.scala 960:32]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_157 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_157 <= r_lvl_output_ff_valid_125; // @[FanNetwork.scala 963:32]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_158 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_158 <= r_lvl_output_ff_valid_126; // @[FanNetwork.scala 966:32]
    end
    if (reset) begin // @[FanNetwork.scala 46:40]
      r_lvl_output_ff_valid_159 <= 1'h0; // @[FanNetwork.scala 46:40]
    end else begin
      r_lvl_output_ff_valid_159 <= r_lvl_output_ff_valid_127; // @[FanNetwork.scala 969:32]
    end
    if (reset) begin // @[FanNetwork.scala 47:26]
      r_valid_0 <= 1'h0; // @[FanNetwork.scala 47:26]
    end else begin
      r_valid_0 <= io_i_valid;
    end
    if (reset) begin // @[FanNetwork.scala 47:26]
      r_valid_1 <= 1'h0; // @[FanNetwork.scala 47:26]
    end else begin
      r_valid_1 <= r_valid_0; // @[FanNetwork.scala 980:24]
    end
    if (reset) begin // @[FanNetwork.scala 47:26]
      r_valid_2 <= 1'h0; // @[FanNetwork.scala 47:26]
    end else begin
      r_valid_2 <= r_valid_1; // @[FanNetwork.scala 980:24]
    end
    if (reset) begin // @[FanNetwork.scala 47:26]
      r_valid_3 <= 1'h0; // @[FanNetwork.scala 47:26]
    end else begin
      r_valid_3 <= r_valid_2; // @[FanNetwork.scala 980:24]
    end
    if (reset) begin // @[FanNetwork.scala 47:26]
      r_valid_4 <= 1'h0; // @[FanNetwork.scala 47:26]
    end else begin
      r_valid_4 <= r_valid_3; // @[FanNetwork.scala 980:24]
    end
    if (reset) begin // @[FanNetwork.scala 49:30]
      r_final_sum <= 32'h0; // @[FanNetwork.scala 49:30]
    end else begin
      r_final_sum <= w_fan_lvl_4_0; // @[FanNetwork.scala 1513:17]
    end
    if (reset) begin // @[FanNetwork.scala 50:30]
      r_final_add <= 1'h0; // @[FanNetwork.scala 50:30]
    end else begin
      r_final_add <= io_i_add_en_bus_30; // @[FanNetwork.scala 1511:17]
    end
    if (reset) begin // @[FanNetwork.scala 51:31]
      r_final_add2 <= 1'h0; // @[FanNetwork.scala 51:31]
    end else begin
      r_final_add2 <= r_final_add; // @[FanNetwork.scala 1512:18]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_fan_ff_lvl_0_to_4_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  r_fan_ff_lvl_0_to_4_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  r_fan_ff_lvl_0_to_3_0 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  r_fan_ff_lvl_0_to_3_1 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  r_fan_ff_lvl_0_to_3_2 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  r_fan_ff_lvl_0_to_3_3 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  r_fan_ff_lvl_0_to_3_4 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  r_fan_ff_lvl_0_to_3_5 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  r_fan_ff_lvl_0_to_2_0 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  r_fan_ff_lvl_0_to_2_1 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  r_fan_ff_lvl_0_to_2_2 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  r_fan_ff_lvl_0_to_2_3 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  r_fan_ff_lvl_0_to_2_4 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  r_fan_ff_lvl_0_to_2_5 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  r_fan_ff_lvl_0_to_2_6 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  r_fan_ff_lvl_0_to_2_7 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  r_fan_ff_lvl_0_to_2_8 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  r_fan_ff_lvl_0_to_2_9 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  r_fan_ff_lvl_0_to_2_10 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  r_fan_ff_lvl_0_to_2_11 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  r_fan_ff_lvl_0_to_2_12 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  r_fan_ff_lvl_0_to_2_13 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  r_fan_ff_lvl_1_to_4_0 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  r_fan_ff_lvl_1_to_4_1 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  r_fan_ff_lvl_1_to_3_0 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  r_fan_ff_lvl_1_to_3_1 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  r_fan_ff_lvl_1_to_3_2 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  r_fan_ff_lvl_1_to_3_3 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  r_fan_ff_lvl_1_to_3_4 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  r_fan_ff_lvl_1_to_3_5 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  r_fan_ff_lvl_2_to_4_0 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  r_fan_ff_lvl_2_to_4_1 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  r_lvl_output_ff_0 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  r_lvl_output_ff_1 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  r_lvl_output_ff_2 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  r_lvl_output_ff_3 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  r_lvl_output_ff_4 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  r_lvl_output_ff_5 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  r_lvl_output_ff_6 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  r_lvl_output_ff_7 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  r_lvl_output_ff_8 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  r_lvl_output_ff_9 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  r_lvl_output_ff_10 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  r_lvl_output_ff_11 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  r_lvl_output_ff_12 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  r_lvl_output_ff_13 = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  r_lvl_output_ff_14 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  r_lvl_output_ff_15 = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  r_lvl_output_ff_16 = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  r_lvl_output_ff_17 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  r_lvl_output_ff_18 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  r_lvl_output_ff_19 = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  r_lvl_output_ff_20 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  r_lvl_output_ff_21 = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  r_lvl_output_ff_22 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  r_lvl_output_ff_23 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  r_lvl_output_ff_24 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  r_lvl_output_ff_25 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  r_lvl_output_ff_26 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  r_lvl_output_ff_27 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  r_lvl_output_ff_28 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  r_lvl_output_ff_29 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  r_lvl_output_ff_30 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  r_lvl_output_ff_31 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  r_lvl_output_ff_32 = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  r_lvl_output_ff_33 = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  r_lvl_output_ff_34 = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  r_lvl_output_ff_35 = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  r_lvl_output_ff_36 = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  r_lvl_output_ff_37 = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  r_lvl_output_ff_38 = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  r_lvl_output_ff_39 = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  r_lvl_output_ff_40 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  r_lvl_output_ff_41 = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  r_lvl_output_ff_42 = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  r_lvl_output_ff_43 = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  r_lvl_output_ff_44 = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  r_lvl_output_ff_45 = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  r_lvl_output_ff_46 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  r_lvl_output_ff_47 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  r_lvl_output_ff_48 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  r_lvl_output_ff_49 = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  r_lvl_output_ff_50 = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  r_lvl_output_ff_51 = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  r_lvl_output_ff_52 = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  r_lvl_output_ff_53 = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  r_lvl_output_ff_54 = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  r_lvl_output_ff_55 = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  r_lvl_output_ff_56 = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  r_lvl_output_ff_57 = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  r_lvl_output_ff_58 = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  r_lvl_output_ff_59 = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  r_lvl_output_ff_60 = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  r_lvl_output_ff_61 = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  r_lvl_output_ff_62 = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  r_lvl_output_ff_63 = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  r_lvl_output_ff_64 = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  r_lvl_output_ff_65 = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  r_lvl_output_ff_66 = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  r_lvl_output_ff_67 = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  r_lvl_output_ff_68 = _RAND_100[31:0];
  _RAND_101 = {1{`RANDOM}};
  r_lvl_output_ff_69 = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  r_lvl_output_ff_70 = _RAND_102[31:0];
  _RAND_103 = {1{`RANDOM}};
  r_lvl_output_ff_71 = _RAND_103[31:0];
  _RAND_104 = {1{`RANDOM}};
  r_lvl_output_ff_72 = _RAND_104[31:0];
  _RAND_105 = {1{`RANDOM}};
  r_lvl_output_ff_73 = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  r_lvl_output_ff_74 = _RAND_106[31:0];
  _RAND_107 = {1{`RANDOM}};
  r_lvl_output_ff_75 = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  r_lvl_output_ff_76 = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  r_lvl_output_ff_77 = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  r_lvl_output_ff_78 = _RAND_110[31:0];
  _RAND_111 = {1{`RANDOM}};
  r_lvl_output_ff_79 = _RAND_111[31:0];
  _RAND_112 = {1{`RANDOM}};
  r_lvl_output_ff_80 = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  r_lvl_output_ff_81 = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  r_lvl_output_ff_82 = _RAND_114[31:0];
  _RAND_115 = {1{`RANDOM}};
  r_lvl_output_ff_83 = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  r_lvl_output_ff_84 = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  r_lvl_output_ff_85 = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  r_lvl_output_ff_86 = _RAND_118[31:0];
  _RAND_119 = {1{`RANDOM}};
  r_lvl_output_ff_87 = _RAND_119[31:0];
  _RAND_120 = {1{`RANDOM}};
  r_lvl_output_ff_88 = _RAND_120[31:0];
  _RAND_121 = {1{`RANDOM}};
  r_lvl_output_ff_89 = _RAND_121[31:0];
  _RAND_122 = {1{`RANDOM}};
  r_lvl_output_ff_90 = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  r_lvl_output_ff_91 = _RAND_123[31:0];
  _RAND_124 = {1{`RANDOM}};
  r_lvl_output_ff_92 = _RAND_124[31:0];
  _RAND_125 = {1{`RANDOM}};
  r_lvl_output_ff_93 = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  r_lvl_output_ff_94 = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  r_lvl_output_ff_95 = _RAND_127[31:0];
  _RAND_128 = {1{`RANDOM}};
  r_lvl_output_ff_96 = _RAND_128[31:0];
  _RAND_129 = {1{`RANDOM}};
  r_lvl_output_ff_97 = _RAND_129[31:0];
  _RAND_130 = {1{`RANDOM}};
  r_lvl_output_ff_98 = _RAND_130[31:0];
  _RAND_131 = {1{`RANDOM}};
  r_lvl_output_ff_99 = _RAND_131[31:0];
  _RAND_132 = {1{`RANDOM}};
  r_lvl_output_ff_100 = _RAND_132[31:0];
  _RAND_133 = {1{`RANDOM}};
  r_lvl_output_ff_101 = _RAND_133[31:0];
  _RAND_134 = {1{`RANDOM}};
  r_lvl_output_ff_102 = _RAND_134[31:0];
  _RAND_135 = {1{`RANDOM}};
  r_lvl_output_ff_103 = _RAND_135[31:0];
  _RAND_136 = {1{`RANDOM}};
  r_lvl_output_ff_104 = _RAND_136[31:0];
  _RAND_137 = {1{`RANDOM}};
  r_lvl_output_ff_105 = _RAND_137[31:0];
  _RAND_138 = {1{`RANDOM}};
  r_lvl_output_ff_106 = _RAND_138[31:0];
  _RAND_139 = {1{`RANDOM}};
  r_lvl_output_ff_107 = _RAND_139[31:0];
  _RAND_140 = {1{`RANDOM}};
  r_lvl_output_ff_108 = _RAND_140[31:0];
  _RAND_141 = {1{`RANDOM}};
  r_lvl_output_ff_109 = _RAND_141[31:0];
  _RAND_142 = {1{`RANDOM}};
  r_lvl_output_ff_110 = _RAND_142[31:0];
  _RAND_143 = {1{`RANDOM}};
  r_lvl_output_ff_112 = _RAND_143[31:0];
  _RAND_144 = {1{`RANDOM}};
  r_lvl_output_ff_113 = _RAND_144[31:0];
  _RAND_145 = {1{`RANDOM}};
  r_lvl_output_ff_114 = _RAND_145[31:0];
  _RAND_146 = {1{`RANDOM}};
  r_lvl_output_ff_115 = _RAND_146[31:0];
  _RAND_147 = {1{`RANDOM}};
  r_lvl_output_ff_116 = _RAND_147[31:0];
  _RAND_148 = {1{`RANDOM}};
  r_lvl_output_ff_117 = _RAND_148[31:0];
  _RAND_149 = {1{`RANDOM}};
  r_lvl_output_ff_118 = _RAND_149[31:0];
  _RAND_150 = {1{`RANDOM}};
  r_lvl_output_ff_119 = _RAND_150[31:0];
  _RAND_151 = {1{`RANDOM}};
  r_lvl_output_ff_120 = _RAND_151[31:0];
  _RAND_152 = {1{`RANDOM}};
  r_lvl_output_ff_121 = _RAND_152[31:0];
  _RAND_153 = {1{`RANDOM}};
  r_lvl_output_ff_122 = _RAND_153[31:0];
  _RAND_154 = {1{`RANDOM}};
  r_lvl_output_ff_123 = _RAND_154[31:0];
  _RAND_155 = {1{`RANDOM}};
  r_lvl_output_ff_124 = _RAND_155[31:0];
  _RAND_156 = {1{`RANDOM}};
  r_lvl_output_ff_125 = _RAND_156[31:0];
  _RAND_157 = {1{`RANDOM}};
  r_lvl_output_ff_126 = _RAND_157[31:0];
  _RAND_158 = {1{`RANDOM}};
  r_lvl_output_ff_127 = _RAND_158[31:0];
  _RAND_159 = {1{`RANDOM}};
  r_lvl_output_ff_128 = _RAND_159[31:0];
  _RAND_160 = {1{`RANDOM}};
  r_lvl_output_ff_129 = _RAND_160[31:0];
  _RAND_161 = {1{`RANDOM}};
  r_lvl_output_ff_130 = _RAND_161[31:0];
  _RAND_162 = {1{`RANDOM}};
  r_lvl_output_ff_131 = _RAND_162[31:0];
  _RAND_163 = {1{`RANDOM}};
  r_lvl_output_ff_132 = _RAND_163[31:0];
  _RAND_164 = {1{`RANDOM}};
  r_lvl_output_ff_133 = _RAND_164[31:0];
  _RAND_165 = {1{`RANDOM}};
  r_lvl_output_ff_134 = _RAND_165[31:0];
  _RAND_166 = {1{`RANDOM}};
  r_lvl_output_ff_135 = _RAND_166[31:0];
  _RAND_167 = {1{`RANDOM}};
  r_lvl_output_ff_136 = _RAND_167[31:0];
  _RAND_168 = {1{`RANDOM}};
  r_lvl_output_ff_137 = _RAND_168[31:0];
  _RAND_169 = {1{`RANDOM}};
  r_lvl_output_ff_138 = _RAND_169[31:0];
  _RAND_170 = {1{`RANDOM}};
  r_lvl_output_ff_139 = _RAND_170[31:0];
  _RAND_171 = {1{`RANDOM}};
  r_lvl_output_ff_140 = _RAND_171[31:0];
  _RAND_172 = {1{`RANDOM}};
  r_lvl_output_ff_141 = _RAND_172[31:0];
  _RAND_173 = {1{`RANDOM}};
  r_lvl_output_ff_142 = _RAND_173[31:0];
  _RAND_174 = {1{`RANDOM}};
  r_lvl_output_ff_143 = _RAND_174[31:0];
  _RAND_175 = {1{`RANDOM}};
  r_lvl_output_ff_144 = _RAND_175[31:0];
  _RAND_176 = {1{`RANDOM}};
  r_lvl_output_ff_145 = _RAND_176[31:0];
  _RAND_177 = {1{`RANDOM}};
  r_lvl_output_ff_146 = _RAND_177[31:0];
  _RAND_178 = {1{`RANDOM}};
  r_lvl_output_ff_147 = _RAND_178[31:0];
  _RAND_179 = {1{`RANDOM}};
  r_lvl_output_ff_148 = _RAND_179[31:0];
  _RAND_180 = {1{`RANDOM}};
  r_lvl_output_ff_149 = _RAND_180[31:0];
  _RAND_181 = {1{`RANDOM}};
  r_lvl_output_ff_150 = _RAND_181[31:0];
  _RAND_182 = {1{`RANDOM}};
  r_lvl_output_ff_151 = _RAND_182[31:0];
  _RAND_183 = {1{`RANDOM}};
  r_lvl_output_ff_152 = _RAND_183[31:0];
  _RAND_184 = {1{`RANDOM}};
  r_lvl_output_ff_153 = _RAND_184[31:0];
  _RAND_185 = {1{`RANDOM}};
  r_lvl_output_ff_154 = _RAND_185[31:0];
  _RAND_186 = {1{`RANDOM}};
  r_lvl_output_ff_155 = _RAND_186[31:0];
  _RAND_187 = {1{`RANDOM}};
  r_lvl_output_ff_156 = _RAND_187[31:0];
  _RAND_188 = {1{`RANDOM}};
  r_lvl_output_ff_157 = _RAND_188[31:0];
  _RAND_189 = {1{`RANDOM}};
  r_lvl_output_ff_158 = _RAND_189[31:0];
  _RAND_190 = {1{`RANDOM}};
  r_lvl_output_ff_159 = _RAND_190[31:0];
  _RAND_191 = {1{`RANDOM}};
  r_lvl_output_ff_valid_0 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  r_lvl_output_ff_valid_1 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  r_lvl_output_ff_valid_2 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  r_lvl_output_ff_valid_3 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  r_lvl_output_ff_valid_4 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  r_lvl_output_ff_valid_5 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  r_lvl_output_ff_valid_6 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  r_lvl_output_ff_valid_7 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  r_lvl_output_ff_valid_8 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  r_lvl_output_ff_valid_9 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  r_lvl_output_ff_valid_10 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  r_lvl_output_ff_valid_11 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  r_lvl_output_ff_valid_12 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  r_lvl_output_ff_valid_13 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  r_lvl_output_ff_valid_14 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  r_lvl_output_ff_valid_15 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  r_lvl_output_ff_valid_16 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  r_lvl_output_ff_valid_17 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  r_lvl_output_ff_valid_18 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  r_lvl_output_ff_valid_19 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  r_lvl_output_ff_valid_20 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  r_lvl_output_ff_valid_21 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  r_lvl_output_ff_valid_22 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  r_lvl_output_ff_valid_23 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  r_lvl_output_ff_valid_24 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  r_lvl_output_ff_valid_25 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  r_lvl_output_ff_valid_26 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  r_lvl_output_ff_valid_27 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  r_lvl_output_ff_valid_28 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  r_lvl_output_ff_valid_29 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  r_lvl_output_ff_valid_30 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  r_lvl_output_ff_valid_31 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  r_lvl_output_ff_valid_32 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  r_lvl_output_ff_valid_33 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  r_lvl_output_ff_valid_34 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  r_lvl_output_ff_valid_35 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  r_lvl_output_ff_valid_36 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  r_lvl_output_ff_valid_37 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  r_lvl_output_ff_valid_38 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  r_lvl_output_ff_valid_39 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  r_lvl_output_ff_valid_40 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  r_lvl_output_ff_valid_41 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  r_lvl_output_ff_valid_42 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  r_lvl_output_ff_valid_43 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  r_lvl_output_ff_valid_44 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  r_lvl_output_ff_valid_45 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  r_lvl_output_ff_valid_46 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  r_lvl_output_ff_valid_47 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  r_lvl_output_ff_valid_48 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  r_lvl_output_ff_valid_49 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  r_lvl_output_ff_valid_50 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  r_lvl_output_ff_valid_51 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  r_lvl_output_ff_valid_52 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  r_lvl_output_ff_valid_53 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  r_lvl_output_ff_valid_54 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  r_lvl_output_ff_valid_55 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  r_lvl_output_ff_valid_56 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  r_lvl_output_ff_valid_57 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  r_lvl_output_ff_valid_58 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  r_lvl_output_ff_valid_59 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  r_lvl_output_ff_valid_60 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  r_lvl_output_ff_valid_61 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  r_lvl_output_ff_valid_62 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  r_lvl_output_ff_valid_63 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  r_lvl_output_ff_valid_64 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  r_lvl_output_ff_valid_65 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  r_lvl_output_ff_valid_66 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  r_lvl_output_ff_valid_67 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  r_lvl_output_ff_valid_68 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  r_lvl_output_ff_valid_69 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  r_lvl_output_ff_valid_70 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  r_lvl_output_ff_valid_71 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  r_lvl_output_ff_valid_72 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  r_lvl_output_ff_valid_73 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  r_lvl_output_ff_valid_74 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  r_lvl_output_ff_valid_75 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  r_lvl_output_ff_valid_76 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  r_lvl_output_ff_valid_77 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  r_lvl_output_ff_valid_78 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  r_lvl_output_ff_valid_79 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  r_lvl_output_ff_valid_80 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  r_lvl_output_ff_valid_81 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  r_lvl_output_ff_valid_82 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  r_lvl_output_ff_valid_83 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  r_lvl_output_ff_valid_84 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  r_lvl_output_ff_valid_85 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  r_lvl_output_ff_valid_86 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  r_lvl_output_ff_valid_87 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  r_lvl_output_ff_valid_88 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  r_lvl_output_ff_valid_89 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  r_lvl_output_ff_valid_90 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  r_lvl_output_ff_valid_91 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  r_lvl_output_ff_valid_92 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  r_lvl_output_ff_valid_93 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  r_lvl_output_ff_valid_94 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  r_lvl_output_ff_valid_95 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  r_lvl_output_ff_valid_96 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  r_lvl_output_ff_valid_97 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  r_lvl_output_ff_valid_98 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  r_lvl_output_ff_valid_99 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  r_lvl_output_ff_valid_100 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  r_lvl_output_ff_valid_101 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  r_lvl_output_ff_valid_102 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  r_lvl_output_ff_valid_103 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  r_lvl_output_ff_valid_104 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  r_lvl_output_ff_valid_105 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  r_lvl_output_ff_valid_106 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  r_lvl_output_ff_valid_107 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  r_lvl_output_ff_valid_108 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  r_lvl_output_ff_valid_109 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  r_lvl_output_ff_valid_110 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  r_lvl_output_ff_valid_111 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  r_lvl_output_ff_valid_112 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  r_lvl_output_ff_valid_113 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  r_lvl_output_ff_valid_114 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  r_lvl_output_ff_valid_115 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  r_lvl_output_ff_valid_116 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  r_lvl_output_ff_valid_117 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  r_lvl_output_ff_valid_118 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  r_lvl_output_ff_valid_119 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  r_lvl_output_ff_valid_120 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  r_lvl_output_ff_valid_121 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  r_lvl_output_ff_valid_122 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  r_lvl_output_ff_valid_123 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  r_lvl_output_ff_valid_124 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  r_lvl_output_ff_valid_125 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  r_lvl_output_ff_valid_126 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  r_lvl_output_ff_valid_127 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  r_lvl_output_ff_valid_128 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  r_lvl_output_ff_valid_129 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  r_lvl_output_ff_valid_130 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  r_lvl_output_ff_valid_131 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  r_lvl_output_ff_valid_132 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  r_lvl_output_ff_valid_133 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  r_lvl_output_ff_valid_134 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  r_lvl_output_ff_valid_135 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  r_lvl_output_ff_valid_136 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  r_lvl_output_ff_valid_137 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  r_lvl_output_ff_valid_138 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  r_lvl_output_ff_valid_139 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  r_lvl_output_ff_valid_140 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  r_lvl_output_ff_valid_141 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  r_lvl_output_ff_valid_142 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  r_lvl_output_ff_valid_143 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  r_lvl_output_ff_valid_144 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  r_lvl_output_ff_valid_145 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  r_lvl_output_ff_valid_146 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  r_lvl_output_ff_valid_147 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  r_lvl_output_ff_valid_148 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  r_lvl_output_ff_valid_149 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  r_lvl_output_ff_valid_150 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  r_lvl_output_ff_valid_151 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  r_lvl_output_ff_valid_152 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  r_lvl_output_ff_valid_153 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  r_lvl_output_ff_valid_154 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  r_lvl_output_ff_valid_155 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  r_lvl_output_ff_valid_156 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  r_lvl_output_ff_valid_157 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  r_lvl_output_ff_valid_158 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  r_lvl_output_ff_valid_159 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  r_valid_0 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  r_valid_1 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  r_valid_2 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  r_valid_3 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  r_valid_4 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  r_final_sum = _RAND_356[31:0];
  _RAND_357 = {1{`RANDOM}};
  r_final_add = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  r_final_add2 = _RAND_358[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module flexdpecom2(
  input         clock,
  input         reset,
  output        io_o_valid_0,
  output        io_o_valid_1,
  output        io_o_valid_2,
  output        io_o_valid_3,
  output        io_o_valid_4,
  output        io_o_valid_5,
  output        io_o_valid_6,
  output        io_o_valid_7,
  output        io_o_valid_8,
  output        io_o_valid_9,
  output        io_o_valid_10,
  output        io_o_valid_11,
  output        io_o_valid_12,
  output        io_o_valid_13,
  output        io_o_valid_14,
  output        io_o_valid_15,
  output        io_o_valid_16,
  output        io_o_valid_17,
  output        io_o_valid_18,
  output        io_o_valid_19,
  output        io_o_valid_20,
  output        io_o_valid_21,
  output        io_o_valid_22,
  output        io_o_valid_23,
  output        io_o_valid_24,
  output        io_o_valid_25,
  output        io_o_valid_26,
  output        io_o_valid_27,
  output        io_o_valid_28,
  output        io_o_valid_29,
  output        io_o_valid_30,
  output        io_o_valid_31,
  output [31:0] io_o_data_bus_0,
  output [31:0] io_o_data_bus_1,
  output [31:0] io_o_data_bus_2,
  output [31:0] io_o_data_bus_3,
  output [31:0] io_o_data_bus_4,
  output [31:0] io_o_data_bus_5,
  output [31:0] io_o_data_bus_6,
  output [31:0] io_o_data_bus_7,
  output [31:0] io_o_data_bus_8,
  output [31:0] io_o_data_bus_9,
  output [31:0] io_o_data_bus_10,
  output [31:0] io_o_data_bus_11,
  output [31:0] io_o_data_bus_12,
  output [31:0] io_o_data_bus_13,
  output [31:0] io_o_data_bus_14,
  output [31:0] io_o_data_bus_15,
  output [31:0] io_o_data_bus_16,
  output [31:0] io_o_data_bus_17,
  output [31:0] io_o_data_bus_18,
  output [31:0] io_o_data_bus_19,
  output [31:0] io_o_data_bus_20,
  output [31:0] io_o_data_bus_21,
  output [31:0] io_o_data_bus_22,
  output [31:0] io_o_data_bus_23,
  output [31:0] io_o_data_bus_24,
  output [31:0] io_o_data_bus_25,
  output [31:0] io_o_data_bus_26,
  output [31:0] io_o_data_bus_27,
  output [31:0] io_o_data_bus_28,
  output [31:0] io_o_data_bus_29,
  output [31:0] io_o_data_bus_30,
  output [31:0] io_o_data_bus_31,
  output [31:0] io_o_adder_0,
  output [31:0] io_o_adder_1,
  output [31:0] io_o_adder_2,
  output [31:0] io_o_adder_3,
  output [31:0] io_o_adder_4,
  output [31:0] io_o_adder_5,
  output [31:0] io_o_adder_6,
  output [31:0] io_o_adder_7,
  output [31:0] io_o_adder_8,
  output [31:0] io_o_adder_9,
  output [31:0] io_o_adder_10,
  output [31:0] io_o_adder_11,
  output [31:0] io_o_adder_12,
  output [31:0] io_o_adder_13,
  output [31:0] io_o_adder_14,
  output [31:0] io_o_adder_15,
  output [31:0] io_o_adder_16,
  output [31:0] io_o_adder_17,
  output [31:0] io_o_adder_18,
  output [31:0] io_o_adder_19,
  output [31:0] io_o_adder_20,
  output [31:0] io_o_adder_21,
  output [31:0] io_o_adder_22,
  output [31:0] io_o_adder_23,
  output [31:0] io_o_adder_24,
  output [31:0] io_o_adder_25,
  output [31:0] io_o_adder_26,
  output [31:0] io_o_adder_27,
  output [31:0] io_o_adder_28,
  output [31:0] io_o_adder_29,
  output [31:0] io_o_adder_30
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
`endif // RANDOMIZE_REG_INIT
  wire  my_controller_clock; // @[FlexDPE.scala 40:31]
  wire  my_controller_reset; // @[FlexDPE.scala 40:31]
  wire  my_controller_io_o_reduction_add_0; // @[FlexDPE.scala 40:31]
  wire  my_controller_io_o_reduction_add_1; // @[FlexDPE.scala 40:31]
  wire  my_controller_io_o_reduction_add_2; // @[FlexDPE.scala 40:31]
  wire  my_controller_io_o_reduction_add_3; // @[FlexDPE.scala 40:31]
  wire  my_controller_io_o_reduction_add_4; // @[FlexDPE.scala 40:31]
  wire  my_controller_io_o_reduction_add_5; // @[FlexDPE.scala 40:31]
  wire  my_controller_io_o_reduction_add_6; // @[FlexDPE.scala 40:31]
  wire  my_controller_io_o_reduction_add_7; // @[FlexDPE.scala 40:31]
  wire  my_controller_io_o_reduction_add_8; // @[FlexDPE.scala 40:31]
  wire  my_controller_io_o_reduction_add_9; // @[FlexDPE.scala 40:31]
  wire  my_controller_io_o_reduction_add_10; // @[FlexDPE.scala 40:31]
  wire  my_controller_io_o_reduction_add_11; // @[FlexDPE.scala 40:31]
  wire  my_controller_io_o_reduction_add_12; // @[FlexDPE.scala 40:31]
  wire  my_controller_io_o_reduction_add_13; // @[FlexDPE.scala 40:31]
  wire  my_controller_io_o_reduction_add_14; // @[FlexDPE.scala 40:31]
  wire  my_controller_io_o_reduction_add_15; // @[FlexDPE.scala 40:31]
  wire  my_controller_io_o_reduction_add_16; // @[FlexDPE.scala 40:31]
  wire  my_controller_io_o_reduction_add_17; // @[FlexDPE.scala 40:31]
  wire  my_controller_io_o_reduction_add_18; // @[FlexDPE.scala 40:31]
  wire  my_controller_io_o_reduction_add_19; // @[FlexDPE.scala 40:31]
  wire  my_controller_io_o_reduction_add_20; // @[FlexDPE.scala 40:31]
  wire  my_controller_io_o_reduction_add_21; // @[FlexDPE.scala 40:31]
  wire  my_controller_io_o_reduction_add_22; // @[FlexDPE.scala 40:31]
  wire  my_controller_io_o_reduction_add_23; // @[FlexDPE.scala 40:31]
  wire  my_controller_io_o_reduction_add_24; // @[FlexDPE.scala 40:31]
  wire  my_controller_io_o_reduction_add_25; // @[FlexDPE.scala 40:31]
  wire  my_controller_io_o_reduction_add_26; // @[FlexDPE.scala 40:31]
  wire  my_controller_io_o_reduction_add_27; // @[FlexDPE.scala 40:31]
  wire  my_controller_io_o_reduction_add_28; // @[FlexDPE.scala 40:31]
  wire  my_controller_io_o_reduction_add_29; // @[FlexDPE.scala 40:31]
  wire  my_controller_io_o_reduction_add_30; // @[FlexDPE.scala 40:31]
  wire [2:0] my_controller_io_o_reduction_cmd_0; // @[FlexDPE.scala 40:31]
  wire [2:0] my_controller_io_o_reduction_cmd_1; // @[FlexDPE.scala 40:31]
  wire [2:0] my_controller_io_o_reduction_cmd_2; // @[FlexDPE.scala 40:31]
  wire [2:0] my_controller_io_o_reduction_cmd_3; // @[FlexDPE.scala 40:31]
  wire [2:0] my_controller_io_o_reduction_cmd_4; // @[FlexDPE.scala 40:31]
  wire [2:0] my_controller_io_o_reduction_cmd_5; // @[FlexDPE.scala 40:31]
  wire [2:0] my_controller_io_o_reduction_cmd_6; // @[FlexDPE.scala 40:31]
  wire [2:0] my_controller_io_o_reduction_cmd_7; // @[FlexDPE.scala 40:31]
  wire [2:0] my_controller_io_o_reduction_cmd_8; // @[FlexDPE.scala 40:31]
  wire [2:0] my_controller_io_o_reduction_cmd_9; // @[FlexDPE.scala 40:31]
  wire [2:0] my_controller_io_o_reduction_cmd_10; // @[FlexDPE.scala 40:31]
  wire [2:0] my_controller_io_o_reduction_cmd_11; // @[FlexDPE.scala 40:31]
  wire [2:0] my_controller_io_o_reduction_cmd_12; // @[FlexDPE.scala 40:31]
  wire [2:0] my_controller_io_o_reduction_cmd_13; // @[FlexDPE.scala 40:31]
  wire [2:0] my_controller_io_o_reduction_cmd_14; // @[FlexDPE.scala 40:31]
  wire [2:0] my_controller_io_o_reduction_cmd_15; // @[FlexDPE.scala 40:31]
  wire [2:0] my_controller_io_o_reduction_cmd_16; // @[FlexDPE.scala 40:31]
  wire [2:0] my_controller_io_o_reduction_cmd_17; // @[FlexDPE.scala 40:31]
  wire [2:0] my_controller_io_o_reduction_cmd_18; // @[FlexDPE.scala 40:31]
  wire [2:0] my_controller_io_o_reduction_cmd_19; // @[FlexDPE.scala 40:31]
  wire [2:0] my_controller_io_o_reduction_cmd_20; // @[FlexDPE.scala 40:31]
  wire [2:0] my_controller_io_o_reduction_cmd_21; // @[FlexDPE.scala 40:31]
  wire [2:0] my_controller_io_o_reduction_cmd_22; // @[FlexDPE.scala 40:31]
  wire [2:0] my_controller_io_o_reduction_cmd_23; // @[FlexDPE.scala 40:31]
  wire [2:0] my_controller_io_o_reduction_cmd_24; // @[FlexDPE.scala 40:31]
  wire [2:0] my_controller_io_o_reduction_cmd_25; // @[FlexDPE.scala 40:31]
  wire [2:0] my_controller_io_o_reduction_cmd_26; // @[FlexDPE.scala 40:31]
  wire [2:0] my_controller_io_o_reduction_cmd_27; // @[FlexDPE.scala 40:31]
  wire [2:0] my_controller_io_o_reduction_cmd_28; // @[FlexDPE.scala 40:31]
  wire [2:0] my_controller_io_o_reduction_cmd_29; // @[FlexDPE.scala 40:31]
  wire [2:0] my_controller_io_o_reduction_cmd_30; // @[FlexDPE.scala 40:31]
  wire [1:0] my_controller_io_o_reduction_sel_0; // @[FlexDPE.scala 40:31]
  wire [1:0] my_controller_io_o_reduction_sel_1; // @[FlexDPE.scala 40:31]
  wire [1:0] my_controller_io_o_reduction_sel_2; // @[FlexDPE.scala 40:31]
  wire [1:0] my_controller_io_o_reduction_sel_3; // @[FlexDPE.scala 40:31]
  wire [1:0] my_controller_io_o_reduction_sel_4; // @[FlexDPE.scala 40:31]
  wire [1:0] my_controller_io_o_reduction_sel_5; // @[FlexDPE.scala 40:31]
  wire [1:0] my_controller_io_o_reduction_sel_6; // @[FlexDPE.scala 40:31]
  wire [1:0] my_controller_io_o_reduction_sel_7; // @[FlexDPE.scala 40:31]
  wire [1:0] my_controller_io_o_reduction_sel_8; // @[FlexDPE.scala 40:31]
  wire [1:0] my_controller_io_o_reduction_sel_9; // @[FlexDPE.scala 40:31]
  wire [1:0] my_controller_io_o_reduction_sel_10; // @[FlexDPE.scala 40:31]
  wire [1:0] my_controller_io_o_reduction_sel_11; // @[FlexDPE.scala 40:31]
  wire [1:0] my_controller_io_o_reduction_sel_12; // @[FlexDPE.scala 40:31]
  wire [1:0] my_controller_io_o_reduction_sel_13; // @[FlexDPE.scala 40:31]
  wire [1:0] my_controller_io_o_reduction_sel_14; // @[FlexDPE.scala 40:31]
  wire [1:0] my_controller_io_o_reduction_sel_15; // @[FlexDPE.scala 40:31]
  wire [1:0] my_controller_io_o_reduction_sel_16; // @[FlexDPE.scala 40:31]
  wire [1:0] my_controller_io_o_reduction_sel_17; // @[FlexDPE.scala 40:31]
  wire [1:0] my_controller_io_o_reduction_sel_18; // @[FlexDPE.scala 40:31]
  wire [1:0] my_controller_io_o_reduction_sel_19; // @[FlexDPE.scala 40:31]
  wire  my_controller_io_o_reduction_valid; // @[FlexDPE.scala 40:31]
  wire  my_Benes_clock; // @[FlexDPE.scala 50:26]
  wire  my_Benes_reset; // @[FlexDPE.scala 50:26]
  wire [15:0] my_Benes_io_o_dist_bus2_0; // @[FlexDPE.scala 50:26]
  wire [15:0] my_Benes_io_o_dist_bus2_1; // @[FlexDPE.scala 50:26]
  wire [15:0] my_Benes_io_o_dist_bus2_2; // @[FlexDPE.scala 50:26]
  wire [15:0] my_Benes_io_o_dist_bus2_3; // @[FlexDPE.scala 50:26]
  wire [15:0] my_Benes_io_o_dist_bus2_4; // @[FlexDPE.scala 50:26]
  wire [15:0] my_Benes_io_o_dist_bus2_5; // @[FlexDPE.scala 50:26]
  wire [15:0] my_Benes_io_o_dist_bus2_6; // @[FlexDPE.scala 50:26]
  wire [15:0] my_Benes_io_o_dist_bus2_7; // @[FlexDPE.scala 50:26]
  wire [15:0] my_Benes_io_o_dist_bus2_8; // @[FlexDPE.scala 50:26]
  wire [15:0] my_Benes_io_o_dist_bus2_9; // @[FlexDPE.scala 50:26]
  wire [15:0] my_Benes_io_o_dist_bus2_10; // @[FlexDPE.scala 50:26]
  wire [15:0] my_Benes_io_o_dist_bus2_11; // @[FlexDPE.scala 50:26]
  wire [15:0] my_Benes_io_o_dist_bus2_12; // @[FlexDPE.scala 50:26]
  wire [15:0] my_Benes_io_o_dist_bus2_13; // @[FlexDPE.scala 50:26]
  wire [15:0] my_Benes_io_o_dist_bus2_14; // @[FlexDPE.scala 50:26]
  wire [15:0] my_Benes_io_o_dist_bus2_15; // @[FlexDPE.scala 50:26]
  wire [15:0] my_Benes_io_o_dist_bus2_16; // @[FlexDPE.scala 50:26]
  wire [15:0] my_Benes_io_o_dist_bus2_17; // @[FlexDPE.scala 50:26]
  wire [15:0] my_Benes_io_o_dist_bus2_18; // @[FlexDPE.scala 50:26]
  wire [15:0] my_Benes_io_o_dist_bus2_19; // @[FlexDPE.scala 50:26]
  wire [15:0] my_Benes_io_o_dist_bus2_20; // @[FlexDPE.scala 50:26]
  wire [15:0] my_Benes_io_o_dist_bus2_21; // @[FlexDPE.scala 50:26]
  wire [15:0] my_Benes_io_o_dist_bus2_22; // @[FlexDPE.scala 50:26]
  wire [15:0] my_Benes_io_o_dist_bus2_23; // @[FlexDPE.scala 50:26]
  wire [15:0] my_Benes_io_o_dist_bus2_24; // @[FlexDPE.scala 50:26]
  wire [15:0] my_Benes_io_o_dist_bus2_25; // @[FlexDPE.scala 50:26]
  wire [15:0] my_Benes_io_o_dist_bus2_26; // @[FlexDPE.scala 50:26]
  wire [15:0] my_Benes_io_o_dist_bus2_27; // @[FlexDPE.scala 50:26]
  wire [15:0] my_Benes_io_o_dist_bus2_28; // @[FlexDPE.scala 50:26]
  wire [15:0] my_Benes_io_o_dist_bus2_29; // @[FlexDPE.scala 50:26]
  wire [15:0] my_Benes_io_o_dist_bus2_30; // @[FlexDPE.scala 50:26]
  wire [15:0] my_Benes_io_o_dist_bus2_31; // @[FlexDPE.scala 50:26]
  wire [15:0] buffer_mult_io_buffer2_0; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_buffer2_1; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_buffer2_2; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_buffer2_3; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_buffer2_4; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_buffer2_5; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_buffer2_6; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_buffer2_7; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_buffer2_8; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_buffer2_9; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_buffer2_10; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_buffer2_11; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_buffer2_12; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_buffer2_13; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_buffer2_14; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_buffer2_15; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_buffer2_16; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_buffer2_17; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_buffer2_18; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_buffer2_19; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_buffer2_20; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_buffer2_21; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_buffer2_22; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_buffer2_23; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_buffer2_24; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_buffer2_25; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_buffer2_26; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_buffer2_27; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_buffer2_28; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_buffer2_29; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_buffer2_30; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_buffer2_31; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_out_0; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_out_1; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_out_2; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_out_3; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_out_4; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_out_5; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_out_6; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_out_7; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_out_8; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_out_9; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_out_10; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_out_11; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_out_12; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_out_13; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_out_14; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_out_15; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_out_16; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_out_17; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_out_18; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_out_19; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_out_20; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_out_21; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_out_22; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_out_23; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_out_24; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_out_25; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_out_26; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_out_27; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_out_28; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_out_29; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_out_30; // @[FlexDPE.scala 61:30]
  wire [15:0] buffer_mult_io_out_31; // @[FlexDPE.scala 61:30]
  wire  my_fan_network_clock; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_reset; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_i_valid; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_i_data_bus_0; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_i_data_bus_1; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_i_data_bus_2; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_i_data_bus_3; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_i_data_bus_4; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_i_data_bus_5; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_i_data_bus_6; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_i_data_bus_7; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_i_data_bus_8; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_i_data_bus_9; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_i_data_bus_10; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_i_data_bus_11; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_i_data_bus_12; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_i_data_bus_13; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_i_data_bus_14; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_i_data_bus_15; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_i_data_bus_16; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_i_data_bus_17; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_i_data_bus_18; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_i_data_bus_19; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_i_data_bus_20; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_i_data_bus_21; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_i_data_bus_22; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_i_data_bus_23; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_i_data_bus_24; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_i_data_bus_25; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_i_data_bus_26; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_i_data_bus_27; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_i_data_bus_28; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_i_data_bus_29; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_i_data_bus_30; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_i_data_bus_31; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_i_add_en_bus_0; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_i_add_en_bus_1; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_i_add_en_bus_2; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_i_add_en_bus_3; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_i_add_en_bus_4; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_i_add_en_bus_5; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_i_add_en_bus_6; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_i_add_en_bus_7; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_i_add_en_bus_8; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_i_add_en_bus_9; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_i_add_en_bus_10; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_i_add_en_bus_11; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_i_add_en_bus_12; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_i_add_en_bus_13; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_i_add_en_bus_14; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_i_add_en_bus_15; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_i_add_en_bus_16; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_i_add_en_bus_17; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_i_add_en_bus_18; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_i_add_en_bus_19; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_i_add_en_bus_20; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_i_add_en_bus_21; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_i_add_en_bus_22; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_i_add_en_bus_23; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_i_add_en_bus_24; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_i_add_en_bus_25; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_i_add_en_bus_26; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_i_add_en_bus_27; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_i_add_en_bus_28; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_i_add_en_bus_29; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_i_add_en_bus_30; // @[FlexDPE.scala 73:32]
  wire [2:0] my_fan_network_io_i_cmd_bus_0; // @[FlexDPE.scala 73:32]
  wire [2:0] my_fan_network_io_i_cmd_bus_1; // @[FlexDPE.scala 73:32]
  wire [2:0] my_fan_network_io_i_cmd_bus_2; // @[FlexDPE.scala 73:32]
  wire [2:0] my_fan_network_io_i_cmd_bus_3; // @[FlexDPE.scala 73:32]
  wire [2:0] my_fan_network_io_i_cmd_bus_4; // @[FlexDPE.scala 73:32]
  wire [2:0] my_fan_network_io_i_cmd_bus_5; // @[FlexDPE.scala 73:32]
  wire [2:0] my_fan_network_io_i_cmd_bus_6; // @[FlexDPE.scala 73:32]
  wire [2:0] my_fan_network_io_i_cmd_bus_7; // @[FlexDPE.scala 73:32]
  wire [2:0] my_fan_network_io_i_cmd_bus_8; // @[FlexDPE.scala 73:32]
  wire [2:0] my_fan_network_io_i_cmd_bus_9; // @[FlexDPE.scala 73:32]
  wire [2:0] my_fan_network_io_i_cmd_bus_10; // @[FlexDPE.scala 73:32]
  wire [2:0] my_fan_network_io_i_cmd_bus_11; // @[FlexDPE.scala 73:32]
  wire [2:0] my_fan_network_io_i_cmd_bus_12; // @[FlexDPE.scala 73:32]
  wire [2:0] my_fan_network_io_i_cmd_bus_13; // @[FlexDPE.scala 73:32]
  wire [2:0] my_fan_network_io_i_cmd_bus_14; // @[FlexDPE.scala 73:32]
  wire [2:0] my_fan_network_io_i_cmd_bus_15; // @[FlexDPE.scala 73:32]
  wire [2:0] my_fan_network_io_i_cmd_bus_16; // @[FlexDPE.scala 73:32]
  wire [2:0] my_fan_network_io_i_cmd_bus_17; // @[FlexDPE.scala 73:32]
  wire [2:0] my_fan_network_io_i_cmd_bus_18; // @[FlexDPE.scala 73:32]
  wire [2:0] my_fan_network_io_i_cmd_bus_19; // @[FlexDPE.scala 73:32]
  wire [2:0] my_fan_network_io_i_cmd_bus_20; // @[FlexDPE.scala 73:32]
  wire [2:0] my_fan_network_io_i_cmd_bus_21; // @[FlexDPE.scala 73:32]
  wire [2:0] my_fan_network_io_i_cmd_bus_22; // @[FlexDPE.scala 73:32]
  wire [2:0] my_fan_network_io_i_cmd_bus_23; // @[FlexDPE.scala 73:32]
  wire [2:0] my_fan_network_io_i_cmd_bus_24; // @[FlexDPE.scala 73:32]
  wire [2:0] my_fan_network_io_i_cmd_bus_25; // @[FlexDPE.scala 73:32]
  wire [2:0] my_fan_network_io_i_cmd_bus_26; // @[FlexDPE.scala 73:32]
  wire [2:0] my_fan_network_io_i_cmd_bus_27; // @[FlexDPE.scala 73:32]
  wire [2:0] my_fan_network_io_i_cmd_bus_28; // @[FlexDPE.scala 73:32]
  wire [2:0] my_fan_network_io_i_cmd_bus_29; // @[FlexDPE.scala 73:32]
  wire [2:0] my_fan_network_io_i_cmd_bus_30; // @[FlexDPE.scala 73:32]
  wire [1:0] my_fan_network_io_i_sel_bus_0; // @[FlexDPE.scala 73:32]
  wire [1:0] my_fan_network_io_i_sel_bus_1; // @[FlexDPE.scala 73:32]
  wire [1:0] my_fan_network_io_i_sel_bus_2; // @[FlexDPE.scala 73:32]
  wire [1:0] my_fan_network_io_i_sel_bus_3; // @[FlexDPE.scala 73:32]
  wire [1:0] my_fan_network_io_i_sel_bus_4; // @[FlexDPE.scala 73:32]
  wire [1:0] my_fan_network_io_i_sel_bus_5; // @[FlexDPE.scala 73:32]
  wire [1:0] my_fan_network_io_i_sel_bus_6; // @[FlexDPE.scala 73:32]
  wire [1:0] my_fan_network_io_i_sel_bus_7; // @[FlexDPE.scala 73:32]
  wire [1:0] my_fan_network_io_i_sel_bus_8; // @[FlexDPE.scala 73:32]
  wire [1:0] my_fan_network_io_i_sel_bus_9; // @[FlexDPE.scala 73:32]
  wire [1:0] my_fan_network_io_i_sel_bus_10; // @[FlexDPE.scala 73:32]
  wire [1:0] my_fan_network_io_i_sel_bus_11; // @[FlexDPE.scala 73:32]
  wire [1:0] my_fan_network_io_i_sel_bus_12; // @[FlexDPE.scala 73:32]
  wire [1:0] my_fan_network_io_i_sel_bus_13; // @[FlexDPE.scala 73:32]
  wire [1:0] my_fan_network_io_i_sel_bus_14; // @[FlexDPE.scala 73:32]
  wire [1:0] my_fan_network_io_i_sel_bus_15; // @[FlexDPE.scala 73:32]
  wire [1:0] my_fan_network_io_i_sel_bus_16; // @[FlexDPE.scala 73:32]
  wire [1:0] my_fan_network_io_i_sel_bus_17; // @[FlexDPE.scala 73:32]
  wire [1:0] my_fan_network_io_i_sel_bus_18; // @[FlexDPE.scala 73:32]
  wire [1:0] my_fan_network_io_i_sel_bus_19; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_o_valid_0; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_o_valid_1; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_o_valid_2; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_o_valid_3; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_o_valid_4; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_o_valid_5; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_o_valid_6; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_o_valid_7; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_o_valid_8; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_o_valid_9; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_o_valid_10; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_o_valid_11; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_o_valid_12; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_o_valid_13; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_o_valid_14; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_o_valid_15; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_o_valid_16; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_o_valid_17; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_o_valid_18; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_o_valid_19; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_o_valid_20; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_o_valid_21; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_o_valid_22; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_o_valid_23; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_o_valid_24; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_o_valid_25; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_o_valid_26; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_o_valid_27; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_o_valid_28; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_o_valid_29; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_o_valid_30; // @[FlexDPE.scala 73:32]
  wire  my_fan_network_io_o_valid_31; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_data_bus_0; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_data_bus_1; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_data_bus_2; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_data_bus_3; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_data_bus_4; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_data_bus_5; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_data_bus_6; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_data_bus_7; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_data_bus_8; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_data_bus_9; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_data_bus_10; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_data_bus_11; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_data_bus_12; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_data_bus_13; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_data_bus_14; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_data_bus_15; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_data_bus_16; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_data_bus_17; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_data_bus_18; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_data_bus_19; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_data_bus_20; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_data_bus_21; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_data_bus_22; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_data_bus_23; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_data_bus_24; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_data_bus_25; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_data_bus_26; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_data_bus_27; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_data_bus_28; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_data_bus_29; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_data_bus_30; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_data_bus_31; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_adder_0; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_adder_1; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_adder_2; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_adder_3; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_adder_4; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_adder_5; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_adder_6; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_adder_7; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_adder_8; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_adder_9; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_adder_10; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_adder_11; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_adder_12; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_adder_13; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_adder_14; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_adder_15; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_adder_16; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_adder_17; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_adder_18; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_adder_19; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_adder_20; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_adder_21; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_adder_22; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_adder_23; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_adder_24; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_adder_25; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_adder_26; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_adder_27; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_adder_28; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_adder_29; // @[FlexDPE.scala 73:32]
  wire [31:0] my_fan_network_io_o_adder_30; // @[FlexDPE.scala 73:32]
  reg [30:0] r_mult_0; // @[FlexDPE.scala 24:26]
  reg [30:0] r_mult_1; // @[FlexDPE.scala 24:26]
  reg [30:0] r_mult_2; // @[FlexDPE.scala 24:26]
  reg [30:0] r_mult_3; // @[FlexDPE.scala 24:26]
  reg [30:0] r_mult_4; // @[FlexDPE.scala 24:26]
  reg [30:0] r_mult_5; // @[FlexDPE.scala 24:26]
  reg [30:0] r_mult_6; // @[FlexDPE.scala 24:26]
  reg [30:0] r_mult_7; // @[FlexDPE.scala 24:26]
  reg [30:0] r_mult_8; // @[FlexDPE.scala 24:26]
  reg [30:0] r_mult_9; // @[FlexDPE.scala 24:26]
  reg [30:0] r_mult_10; // @[FlexDPE.scala 24:26]
  reg [30:0] r_mult_11; // @[FlexDPE.scala 24:26]
  reg [30:0] r_mult_12; // @[FlexDPE.scala 24:26]
  reg [30:0] r_mult_13; // @[FlexDPE.scala 24:26]
  reg [30:0] r_mult_14; // @[FlexDPE.scala 24:26]
  reg [30:0] r_mult_15; // @[FlexDPE.scala 24:26]
  reg [30:0] r_mult_16; // @[FlexDPE.scala 24:26]
  reg [30:0] r_mult_17; // @[FlexDPE.scala 24:26]
  reg [30:0] r_mult_18; // @[FlexDPE.scala 24:26]
  reg [30:0] r_mult_19; // @[FlexDPE.scala 24:26]
  reg [30:0] r_mult_20; // @[FlexDPE.scala 24:26]
  reg [30:0] r_mult_21; // @[FlexDPE.scala 24:26]
  reg [30:0] r_mult_22; // @[FlexDPE.scala 24:26]
  reg [30:0] r_mult_23; // @[FlexDPE.scala 24:26]
  reg [30:0] r_mult_24; // @[FlexDPE.scala 24:26]
  reg [30:0] r_mult_25; // @[FlexDPE.scala 24:26]
  reg [30:0] r_mult_26; // @[FlexDPE.scala 24:26]
  reg [30:0] r_mult_27; // @[FlexDPE.scala 24:26]
  reg [30:0] r_mult_28; // @[FlexDPE.scala 24:26]
  reg [30:0] r_mult_29; // @[FlexDPE.scala 24:26]
  reg [30:0] r_mult_30; // @[FlexDPE.scala 24:26]
  reg [30:0] r_mult_31; // @[FlexDPE.scala 24:26]
  fancontrol my_controller ( // @[FlexDPE.scala 40:31]
    .clock(my_controller_clock),
    .reset(my_controller_reset),
    .io_o_reduction_add_0(my_controller_io_o_reduction_add_0),
    .io_o_reduction_add_1(my_controller_io_o_reduction_add_1),
    .io_o_reduction_add_2(my_controller_io_o_reduction_add_2),
    .io_o_reduction_add_3(my_controller_io_o_reduction_add_3),
    .io_o_reduction_add_4(my_controller_io_o_reduction_add_4),
    .io_o_reduction_add_5(my_controller_io_o_reduction_add_5),
    .io_o_reduction_add_6(my_controller_io_o_reduction_add_6),
    .io_o_reduction_add_7(my_controller_io_o_reduction_add_7),
    .io_o_reduction_add_8(my_controller_io_o_reduction_add_8),
    .io_o_reduction_add_9(my_controller_io_o_reduction_add_9),
    .io_o_reduction_add_10(my_controller_io_o_reduction_add_10),
    .io_o_reduction_add_11(my_controller_io_o_reduction_add_11),
    .io_o_reduction_add_12(my_controller_io_o_reduction_add_12),
    .io_o_reduction_add_13(my_controller_io_o_reduction_add_13),
    .io_o_reduction_add_14(my_controller_io_o_reduction_add_14),
    .io_o_reduction_add_15(my_controller_io_o_reduction_add_15),
    .io_o_reduction_add_16(my_controller_io_o_reduction_add_16),
    .io_o_reduction_add_17(my_controller_io_o_reduction_add_17),
    .io_o_reduction_add_18(my_controller_io_o_reduction_add_18),
    .io_o_reduction_add_19(my_controller_io_o_reduction_add_19),
    .io_o_reduction_add_20(my_controller_io_o_reduction_add_20),
    .io_o_reduction_add_21(my_controller_io_o_reduction_add_21),
    .io_o_reduction_add_22(my_controller_io_o_reduction_add_22),
    .io_o_reduction_add_23(my_controller_io_o_reduction_add_23),
    .io_o_reduction_add_24(my_controller_io_o_reduction_add_24),
    .io_o_reduction_add_25(my_controller_io_o_reduction_add_25),
    .io_o_reduction_add_26(my_controller_io_o_reduction_add_26),
    .io_o_reduction_add_27(my_controller_io_o_reduction_add_27),
    .io_o_reduction_add_28(my_controller_io_o_reduction_add_28),
    .io_o_reduction_add_29(my_controller_io_o_reduction_add_29),
    .io_o_reduction_add_30(my_controller_io_o_reduction_add_30),
    .io_o_reduction_cmd_0(my_controller_io_o_reduction_cmd_0),
    .io_o_reduction_cmd_1(my_controller_io_o_reduction_cmd_1),
    .io_o_reduction_cmd_2(my_controller_io_o_reduction_cmd_2),
    .io_o_reduction_cmd_3(my_controller_io_o_reduction_cmd_3),
    .io_o_reduction_cmd_4(my_controller_io_o_reduction_cmd_4),
    .io_o_reduction_cmd_5(my_controller_io_o_reduction_cmd_5),
    .io_o_reduction_cmd_6(my_controller_io_o_reduction_cmd_6),
    .io_o_reduction_cmd_7(my_controller_io_o_reduction_cmd_7),
    .io_o_reduction_cmd_8(my_controller_io_o_reduction_cmd_8),
    .io_o_reduction_cmd_9(my_controller_io_o_reduction_cmd_9),
    .io_o_reduction_cmd_10(my_controller_io_o_reduction_cmd_10),
    .io_o_reduction_cmd_11(my_controller_io_o_reduction_cmd_11),
    .io_o_reduction_cmd_12(my_controller_io_o_reduction_cmd_12),
    .io_o_reduction_cmd_13(my_controller_io_o_reduction_cmd_13),
    .io_o_reduction_cmd_14(my_controller_io_o_reduction_cmd_14),
    .io_o_reduction_cmd_15(my_controller_io_o_reduction_cmd_15),
    .io_o_reduction_cmd_16(my_controller_io_o_reduction_cmd_16),
    .io_o_reduction_cmd_17(my_controller_io_o_reduction_cmd_17),
    .io_o_reduction_cmd_18(my_controller_io_o_reduction_cmd_18),
    .io_o_reduction_cmd_19(my_controller_io_o_reduction_cmd_19),
    .io_o_reduction_cmd_20(my_controller_io_o_reduction_cmd_20),
    .io_o_reduction_cmd_21(my_controller_io_o_reduction_cmd_21),
    .io_o_reduction_cmd_22(my_controller_io_o_reduction_cmd_22),
    .io_o_reduction_cmd_23(my_controller_io_o_reduction_cmd_23),
    .io_o_reduction_cmd_24(my_controller_io_o_reduction_cmd_24),
    .io_o_reduction_cmd_25(my_controller_io_o_reduction_cmd_25),
    .io_o_reduction_cmd_26(my_controller_io_o_reduction_cmd_26),
    .io_o_reduction_cmd_27(my_controller_io_o_reduction_cmd_27),
    .io_o_reduction_cmd_28(my_controller_io_o_reduction_cmd_28),
    .io_o_reduction_cmd_29(my_controller_io_o_reduction_cmd_29),
    .io_o_reduction_cmd_30(my_controller_io_o_reduction_cmd_30),
    .io_o_reduction_sel_0(my_controller_io_o_reduction_sel_0),
    .io_o_reduction_sel_1(my_controller_io_o_reduction_sel_1),
    .io_o_reduction_sel_2(my_controller_io_o_reduction_sel_2),
    .io_o_reduction_sel_3(my_controller_io_o_reduction_sel_3),
    .io_o_reduction_sel_4(my_controller_io_o_reduction_sel_4),
    .io_o_reduction_sel_5(my_controller_io_o_reduction_sel_5),
    .io_o_reduction_sel_6(my_controller_io_o_reduction_sel_6),
    .io_o_reduction_sel_7(my_controller_io_o_reduction_sel_7),
    .io_o_reduction_sel_8(my_controller_io_o_reduction_sel_8),
    .io_o_reduction_sel_9(my_controller_io_o_reduction_sel_9),
    .io_o_reduction_sel_10(my_controller_io_o_reduction_sel_10),
    .io_o_reduction_sel_11(my_controller_io_o_reduction_sel_11),
    .io_o_reduction_sel_12(my_controller_io_o_reduction_sel_12),
    .io_o_reduction_sel_13(my_controller_io_o_reduction_sel_13),
    .io_o_reduction_sel_14(my_controller_io_o_reduction_sel_14),
    .io_o_reduction_sel_15(my_controller_io_o_reduction_sel_15),
    .io_o_reduction_sel_16(my_controller_io_o_reduction_sel_16),
    .io_o_reduction_sel_17(my_controller_io_o_reduction_sel_17),
    .io_o_reduction_sel_18(my_controller_io_o_reduction_sel_18),
    .io_o_reduction_sel_19(my_controller_io_o_reduction_sel_19),
    .io_o_reduction_valid(my_controller_io_o_reduction_valid)
  );
  Benes my_Benes ( // @[FlexDPE.scala 50:26]
    .clock(my_Benes_clock),
    .reset(my_Benes_reset),
    .io_o_dist_bus2_0(my_Benes_io_o_dist_bus2_0),
    .io_o_dist_bus2_1(my_Benes_io_o_dist_bus2_1),
    .io_o_dist_bus2_2(my_Benes_io_o_dist_bus2_2),
    .io_o_dist_bus2_3(my_Benes_io_o_dist_bus2_3),
    .io_o_dist_bus2_4(my_Benes_io_o_dist_bus2_4),
    .io_o_dist_bus2_5(my_Benes_io_o_dist_bus2_5),
    .io_o_dist_bus2_6(my_Benes_io_o_dist_bus2_6),
    .io_o_dist_bus2_7(my_Benes_io_o_dist_bus2_7),
    .io_o_dist_bus2_8(my_Benes_io_o_dist_bus2_8),
    .io_o_dist_bus2_9(my_Benes_io_o_dist_bus2_9),
    .io_o_dist_bus2_10(my_Benes_io_o_dist_bus2_10),
    .io_o_dist_bus2_11(my_Benes_io_o_dist_bus2_11),
    .io_o_dist_bus2_12(my_Benes_io_o_dist_bus2_12),
    .io_o_dist_bus2_13(my_Benes_io_o_dist_bus2_13),
    .io_o_dist_bus2_14(my_Benes_io_o_dist_bus2_14),
    .io_o_dist_bus2_15(my_Benes_io_o_dist_bus2_15),
    .io_o_dist_bus2_16(my_Benes_io_o_dist_bus2_16),
    .io_o_dist_bus2_17(my_Benes_io_o_dist_bus2_17),
    .io_o_dist_bus2_18(my_Benes_io_o_dist_bus2_18),
    .io_o_dist_bus2_19(my_Benes_io_o_dist_bus2_19),
    .io_o_dist_bus2_20(my_Benes_io_o_dist_bus2_20),
    .io_o_dist_bus2_21(my_Benes_io_o_dist_bus2_21),
    .io_o_dist_bus2_22(my_Benes_io_o_dist_bus2_22),
    .io_o_dist_bus2_23(my_Benes_io_o_dist_bus2_23),
    .io_o_dist_bus2_24(my_Benes_io_o_dist_bus2_24),
    .io_o_dist_bus2_25(my_Benes_io_o_dist_bus2_25),
    .io_o_dist_bus2_26(my_Benes_io_o_dist_bus2_26),
    .io_o_dist_bus2_27(my_Benes_io_o_dist_bus2_27),
    .io_o_dist_bus2_28(my_Benes_io_o_dist_bus2_28),
    .io_o_dist_bus2_29(my_Benes_io_o_dist_bus2_29),
    .io_o_dist_bus2_30(my_Benes_io_o_dist_bus2_30),
    .io_o_dist_bus2_31(my_Benes_io_o_dist_bus2_31)
  );
  buffer_multiplication buffer_mult ( // @[FlexDPE.scala 61:30]
    .io_buffer2_0(buffer_mult_io_buffer2_0),
    .io_buffer2_1(buffer_mult_io_buffer2_1),
    .io_buffer2_2(buffer_mult_io_buffer2_2),
    .io_buffer2_3(buffer_mult_io_buffer2_3),
    .io_buffer2_4(buffer_mult_io_buffer2_4),
    .io_buffer2_5(buffer_mult_io_buffer2_5),
    .io_buffer2_6(buffer_mult_io_buffer2_6),
    .io_buffer2_7(buffer_mult_io_buffer2_7),
    .io_buffer2_8(buffer_mult_io_buffer2_8),
    .io_buffer2_9(buffer_mult_io_buffer2_9),
    .io_buffer2_10(buffer_mult_io_buffer2_10),
    .io_buffer2_11(buffer_mult_io_buffer2_11),
    .io_buffer2_12(buffer_mult_io_buffer2_12),
    .io_buffer2_13(buffer_mult_io_buffer2_13),
    .io_buffer2_14(buffer_mult_io_buffer2_14),
    .io_buffer2_15(buffer_mult_io_buffer2_15),
    .io_buffer2_16(buffer_mult_io_buffer2_16),
    .io_buffer2_17(buffer_mult_io_buffer2_17),
    .io_buffer2_18(buffer_mult_io_buffer2_18),
    .io_buffer2_19(buffer_mult_io_buffer2_19),
    .io_buffer2_20(buffer_mult_io_buffer2_20),
    .io_buffer2_21(buffer_mult_io_buffer2_21),
    .io_buffer2_22(buffer_mult_io_buffer2_22),
    .io_buffer2_23(buffer_mult_io_buffer2_23),
    .io_buffer2_24(buffer_mult_io_buffer2_24),
    .io_buffer2_25(buffer_mult_io_buffer2_25),
    .io_buffer2_26(buffer_mult_io_buffer2_26),
    .io_buffer2_27(buffer_mult_io_buffer2_27),
    .io_buffer2_28(buffer_mult_io_buffer2_28),
    .io_buffer2_29(buffer_mult_io_buffer2_29),
    .io_buffer2_30(buffer_mult_io_buffer2_30),
    .io_buffer2_31(buffer_mult_io_buffer2_31),
    .io_out_0(buffer_mult_io_out_0),
    .io_out_1(buffer_mult_io_out_1),
    .io_out_2(buffer_mult_io_out_2),
    .io_out_3(buffer_mult_io_out_3),
    .io_out_4(buffer_mult_io_out_4),
    .io_out_5(buffer_mult_io_out_5),
    .io_out_6(buffer_mult_io_out_6),
    .io_out_7(buffer_mult_io_out_7),
    .io_out_8(buffer_mult_io_out_8),
    .io_out_9(buffer_mult_io_out_9),
    .io_out_10(buffer_mult_io_out_10),
    .io_out_11(buffer_mult_io_out_11),
    .io_out_12(buffer_mult_io_out_12),
    .io_out_13(buffer_mult_io_out_13),
    .io_out_14(buffer_mult_io_out_14),
    .io_out_15(buffer_mult_io_out_15),
    .io_out_16(buffer_mult_io_out_16),
    .io_out_17(buffer_mult_io_out_17),
    .io_out_18(buffer_mult_io_out_18),
    .io_out_19(buffer_mult_io_out_19),
    .io_out_20(buffer_mult_io_out_20),
    .io_out_21(buffer_mult_io_out_21),
    .io_out_22(buffer_mult_io_out_22),
    .io_out_23(buffer_mult_io_out_23),
    .io_out_24(buffer_mult_io_out_24),
    .io_out_25(buffer_mult_io_out_25),
    .io_out_26(buffer_mult_io_out_26),
    .io_out_27(buffer_mult_io_out_27),
    .io_out_28(buffer_mult_io_out_28),
    .io_out_29(buffer_mult_io_out_29),
    .io_out_30(buffer_mult_io_out_30),
    .io_out_31(buffer_mult_io_out_31)
  );
  FanNetworkcom my_fan_network ( // @[FlexDPE.scala 73:32]
    .clock(my_fan_network_clock),
    .reset(my_fan_network_reset),
    .io_i_valid(my_fan_network_io_i_valid),
    .io_i_data_bus_0(my_fan_network_io_i_data_bus_0),
    .io_i_data_bus_1(my_fan_network_io_i_data_bus_1),
    .io_i_data_bus_2(my_fan_network_io_i_data_bus_2),
    .io_i_data_bus_3(my_fan_network_io_i_data_bus_3),
    .io_i_data_bus_4(my_fan_network_io_i_data_bus_4),
    .io_i_data_bus_5(my_fan_network_io_i_data_bus_5),
    .io_i_data_bus_6(my_fan_network_io_i_data_bus_6),
    .io_i_data_bus_7(my_fan_network_io_i_data_bus_7),
    .io_i_data_bus_8(my_fan_network_io_i_data_bus_8),
    .io_i_data_bus_9(my_fan_network_io_i_data_bus_9),
    .io_i_data_bus_10(my_fan_network_io_i_data_bus_10),
    .io_i_data_bus_11(my_fan_network_io_i_data_bus_11),
    .io_i_data_bus_12(my_fan_network_io_i_data_bus_12),
    .io_i_data_bus_13(my_fan_network_io_i_data_bus_13),
    .io_i_data_bus_14(my_fan_network_io_i_data_bus_14),
    .io_i_data_bus_15(my_fan_network_io_i_data_bus_15),
    .io_i_data_bus_16(my_fan_network_io_i_data_bus_16),
    .io_i_data_bus_17(my_fan_network_io_i_data_bus_17),
    .io_i_data_bus_18(my_fan_network_io_i_data_bus_18),
    .io_i_data_bus_19(my_fan_network_io_i_data_bus_19),
    .io_i_data_bus_20(my_fan_network_io_i_data_bus_20),
    .io_i_data_bus_21(my_fan_network_io_i_data_bus_21),
    .io_i_data_bus_22(my_fan_network_io_i_data_bus_22),
    .io_i_data_bus_23(my_fan_network_io_i_data_bus_23),
    .io_i_data_bus_24(my_fan_network_io_i_data_bus_24),
    .io_i_data_bus_25(my_fan_network_io_i_data_bus_25),
    .io_i_data_bus_26(my_fan_network_io_i_data_bus_26),
    .io_i_data_bus_27(my_fan_network_io_i_data_bus_27),
    .io_i_data_bus_28(my_fan_network_io_i_data_bus_28),
    .io_i_data_bus_29(my_fan_network_io_i_data_bus_29),
    .io_i_data_bus_30(my_fan_network_io_i_data_bus_30),
    .io_i_data_bus_31(my_fan_network_io_i_data_bus_31),
    .io_i_add_en_bus_0(my_fan_network_io_i_add_en_bus_0),
    .io_i_add_en_bus_1(my_fan_network_io_i_add_en_bus_1),
    .io_i_add_en_bus_2(my_fan_network_io_i_add_en_bus_2),
    .io_i_add_en_bus_3(my_fan_network_io_i_add_en_bus_3),
    .io_i_add_en_bus_4(my_fan_network_io_i_add_en_bus_4),
    .io_i_add_en_bus_5(my_fan_network_io_i_add_en_bus_5),
    .io_i_add_en_bus_6(my_fan_network_io_i_add_en_bus_6),
    .io_i_add_en_bus_7(my_fan_network_io_i_add_en_bus_7),
    .io_i_add_en_bus_8(my_fan_network_io_i_add_en_bus_8),
    .io_i_add_en_bus_9(my_fan_network_io_i_add_en_bus_9),
    .io_i_add_en_bus_10(my_fan_network_io_i_add_en_bus_10),
    .io_i_add_en_bus_11(my_fan_network_io_i_add_en_bus_11),
    .io_i_add_en_bus_12(my_fan_network_io_i_add_en_bus_12),
    .io_i_add_en_bus_13(my_fan_network_io_i_add_en_bus_13),
    .io_i_add_en_bus_14(my_fan_network_io_i_add_en_bus_14),
    .io_i_add_en_bus_15(my_fan_network_io_i_add_en_bus_15),
    .io_i_add_en_bus_16(my_fan_network_io_i_add_en_bus_16),
    .io_i_add_en_bus_17(my_fan_network_io_i_add_en_bus_17),
    .io_i_add_en_bus_18(my_fan_network_io_i_add_en_bus_18),
    .io_i_add_en_bus_19(my_fan_network_io_i_add_en_bus_19),
    .io_i_add_en_bus_20(my_fan_network_io_i_add_en_bus_20),
    .io_i_add_en_bus_21(my_fan_network_io_i_add_en_bus_21),
    .io_i_add_en_bus_22(my_fan_network_io_i_add_en_bus_22),
    .io_i_add_en_bus_23(my_fan_network_io_i_add_en_bus_23),
    .io_i_add_en_bus_24(my_fan_network_io_i_add_en_bus_24),
    .io_i_add_en_bus_25(my_fan_network_io_i_add_en_bus_25),
    .io_i_add_en_bus_26(my_fan_network_io_i_add_en_bus_26),
    .io_i_add_en_bus_27(my_fan_network_io_i_add_en_bus_27),
    .io_i_add_en_bus_28(my_fan_network_io_i_add_en_bus_28),
    .io_i_add_en_bus_29(my_fan_network_io_i_add_en_bus_29),
    .io_i_add_en_bus_30(my_fan_network_io_i_add_en_bus_30),
    .io_i_cmd_bus_0(my_fan_network_io_i_cmd_bus_0),
    .io_i_cmd_bus_1(my_fan_network_io_i_cmd_bus_1),
    .io_i_cmd_bus_2(my_fan_network_io_i_cmd_bus_2),
    .io_i_cmd_bus_3(my_fan_network_io_i_cmd_bus_3),
    .io_i_cmd_bus_4(my_fan_network_io_i_cmd_bus_4),
    .io_i_cmd_bus_5(my_fan_network_io_i_cmd_bus_5),
    .io_i_cmd_bus_6(my_fan_network_io_i_cmd_bus_6),
    .io_i_cmd_bus_7(my_fan_network_io_i_cmd_bus_7),
    .io_i_cmd_bus_8(my_fan_network_io_i_cmd_bus_8),
    .io_i_cmd_bus_9(my_fan_network_io_i_cmd_bus_9),
    .io_i_cmd_bus_10(my_fan_network_io_i_cmd_bus_10),
    .io_i_cmd_bus_11(my_fan_network_io_i_cmd_bus_11),
    .io_i_cmd_bus_12(my_fan_network_io_i_cmd_bus_12),
    .io_i_cmd_bus_13(my_fan_network_io_i_cmd_bus_13),
    .io_i_cmd_bus_14(my_fan_network_io_i_cmd_bus_14),
    .io_i_cmd_bus_15(my_fan_network_io_i_cmd_bus_15),
    .io_i_cmd_bus_16(my_fan_network_io_i_cmd_bus_16),
    .io_i_cmd_bus_17(my_fan_network_io_i_cmd_bus_17),
    .io_i_cmd_bus_18(my_fan_network_io_i_cmd_bus_18),
    .io_i_cmd_bus_19(my_fan_network_io_i_cmd_bus_19),
    .io_i_cmd_bus_20(my_fan_network_io_i_cmd_bus_20),
    .io_i_cmd_bus_21(my_fan_network_io_i_cmd_bus_21),
    .io_i_cmd_bus_22(my_fan_network_io_i_cmd_bus_22),
    .io_i_cmd_bus_23(my_fan_network_io_i_cmd_bus_23),
    .io_i_cmd_bus_24(my_fan_network_io_i_cmd_bus_24),
    .io_i_cmd_bus_25(my_fan_network_io_i_cmd_bus_25),
    .io_i_cmd_bus_26(my_fan_network_io_i_cmd_bus_26),
    .io_i_cmd_bus_27(my_fan_network_io_i_cmd_bus_27),
    .io_i_cmd_bus_28(my_fan_network_io_i_cmd_bus_28),
    .io_i_cmd_bus_29(my_fan_network_io_i_cmd_bus_29),
    .io_i_cmd_bus_30(my_fan_network_io_i_cmd_bus_30),
    .io_i_sel_bus_0(my_fan_network_io_i_sel_bus_0),
    .io_i_sel_bus_1(my_fan_network_io_i_sel_bus_1),
    .io_i_sel_bus_2(my_fan_network_io_i_sel_bus_2),
    .io_i_sel_bus_3(my_fan_network_io_i_sel_bus_3),
    .io_i_sel_bus_4(my_fan_network_io_i_sel_bus_4),
    .io_i_sel_bus_5(my_fan_network_io_i_sel_bus_5),
    .io_i_sel_bus_6(my_fan_network_io_i_sel_bus_6),
    .io_i_sel_bus_7(my_fan_network_io_i_sel_bus_7),
    .io_i_sel_bus_8(my_fan_network_io_i_sel_bus_8),
    .io_i_sel_bus_9(my_fan_network_io_i_sel_bus_9),
    .io_i_sel_bus_10(my_fan_network_io_i_sel_bus_10),
    .io_i_sel_bus_11(my_fan_network_io_i_sel_bus_11),
    .io_i_sel_bus_12(my_fan_network_io_i_sel_bus_12),
    .io_i_sel_bus_13(my_fan_network_io_i_sel_bus_13),
    .io_i_sel_bus_14(my_fan_network_io_i_sel_bus_14),
    .io_i_sel_bus_15(my_fan_network_io_i_sel_bus_15),
    .io_i_sel_bus_16(my_fan_network_io_i_sel_bus_16),
    .io_i_sel_bus_17(my_fan_network_io_i_sel_bus_17),
    .io_i_sel_bus_18(my_fan_network_io_i_sel_bus_18),
    .io_i_sel_bus_19(my_fan_network_io_i_sel_bus_19),
    .io_o_valid_0(my_fan_network_io_o_valid_0),
    .io_o_valid_1(my_fan_network_io_o_valid_1),
    .io_o_valid_2(my_fan_network_io_o_valid_2),
    .io_o_valid_3(my_fan_network_io_o_valid_3),
    .io_o_valid_4(my_fan_network_io_o_valid_4),
    .io_o_valid_5(my_fan_network_io_o_valid_5),
    .io_o_valid_6(my_fan_network_io_o_valid_6),
    .io_o_valid_7(my_fan_network_io_o_valid_7),
    .io_o_valid_8(my_fan_network_io_o_valid_8),
    .io_o_valid_9(my_fan_network_io_o_valid_9),
    .io_o_valid_10(my_fan_network_io_o_valid_10),
    .io_o_valid_11(my_fan_network_io_o_valid_11),
    .io_o_valid_12(my_fan_network_io_o_valid_12),
    .io_o_valid_13(my_fan_network_io_o_valid_13),
    .io_o_valid_14(my_fan_network_io_o_valid_14),
    .io_o_valid_15(my_fan_network_io_o_valid_15),
    .io_o_valid_16(my_fan_network_io_o_valid_16),
    .io_o_valid_17(my_fan_network_io_o_valid_17),
    .io_o_valid_18(my_fan_network_io_o_valid_18),
    .io_o_valid_19(my_fan_network_io_o_valid_19),
    .io_o_valid_20(my_fan_network_io_o_valid_20),
    .io_o_valid_21(my_fan_network_io_o_valid_21),
    .io_o_valid_22(my_fan_network_io_o_valid_22),
    .io_o_valid_23(my_fan_network_io_o_valid_23),
    .io_o_valid_24(my_fan_network_io_o_valid_24),
    .io_o_valid_25(my_fan_network_io_o_valid_25),
    .io_o_valid_26(my_fan_network_io_o_valid_26),
    .io_o_valid_27(my_fan_network_io_o_valid_27),
    .io_o_valid_28(my_fan_network_io_o_valid_28),
    .io_o_valid_29(my_fan_network_io_o_valid_29),
    .io_o_valid_30(my_fan_network_io_o_valid_30),
    .io_o_valid_31(my_fan_network_io_o_valid_31),
    .io_o_data_bus_0(my_fan_network_io_o_data_bus_0),
    .io_o_data_bus_1(my_fan_network_io_o_data_bus_1),
    .io_o_data_bus_2(my_fan_network_io_o_data_bus_2),
    .io_o_data_bus_3(my_fan_network_io_o_data_bus_3),
    .io_o_data_bus_4(my_fan_network_io_o_data_bus_4),
    .io_o_data_bus_5(my_fan_network_io_o_data_bus_5),
    .io_o_data_bus_6(my_fan_network_io_o_data_bus_6),
    .io_o_data_bus_7(my_fan_network_io_o_data_bus_7),
    .io_o_data_bus_8(my_fan_network_io_o_data_bus_8),
    .io_o_data_bus_9(my_fan_network_io_o_data_bus_9),
    .io_o_data_bus_10(my_fan_network_io_o_data_bus_10),
    .io_o_data_bus_11(my_fan_network_io_o_data_bus_11),
    .io_o_data_bus_12(my_fan_network_io_o_data_bus_12),
    .io_o_data_bus_13(my_fan_network_io_o_data_bus_13),
    .io_o_data_bus_14(my_fan_network_io_o_data_bus_14),
    .io_o_data_bus_15(my_fan_network_io_o_data_bus_15),
    .io_o_data_bus_16(my_fan_network_io_o_data_bus_16),
    .io_o_data_bus_17(my_fan_network_io_o_data_bus_17),
    .io_o_data_bus_18(my_fan_network_io_o_data_bus_18),
    .io_o_data_bus_19(my_fan_network_io_o_data_bus_19),
    .io_o_data_bus_20(my_fan_network_io_o_data_bus_20),
    .io_o_data_bus_21(my_fan_network_io_o_data_bus_21),
    .io_o_data_bus_22(my_fan_network_io_o_data_bus_22),
    .io_o_data_bus_23(my_fan_network_io_o_data_bus_23),
    .io_o_data_bus_24(my_fan_network_io_o_data_bus_24),
    .io_o_data_bus_25(my_fan_network_io_o_data_bus_25),
    .io_o_data_bus_26(my_fan_network_io_o_data_bus_26),
    .io_o_data_bus_27(my_fan_network_io_o_data_bus_27),
    .io_o_data_bus_28(my_fan_network_io_o_data_bus_28),
    .io_o_data_bus_29(my_fan_network_io_o_data_bus_29),
    .io_o_data_bus_30(my_fan_network_io_o_data_bus_30),
    .io_o_data_bus_31(my_fan_network_io_o_data_bus_31),
    .io_o_adder_0(my_fan_network_io_o_adder_0),
    .io_o_adder_1(my_fan_network_io_o_adder_1),
    .io_o_adder_2(my_fan_network_io_o_adder_2),
    .io_o_adder_3(my_fan_network_io_o_adder_3),
    .io_o_adder_4(my_fan_network_io_o_adder_4),
    .io_o_adder_5(my_fan_network_io_o_adder_5),
    .io_o_adder_6(my_fan_network_io_o_adder_6),
    .io_o_adder_7(my_fan_network_io_o_adder_7),
    .io_o_adder_8(my_fan_network_io_o_adder_8),
    .io_o_adder_9(my_fan_network_io_o_adder_9),
    .io_o_adder_10(my_fan_network_io_o_adder_10),
    .io_o_adder_11(my_fan_network_io_o_adder_11),
    .io_o_adder_12(my_fan_network_io_o_adder_12),
    .io_o_adder_13(my_fan_network_io_o_adder_13),
    .io_o_adder_14(my_fan_network_io_o_adder_14),
    .io_o_adder_15(my_fan_network_io_o_adder_15),
    .io_o_adder_16(my_fan_network_io_o_adder_16),
    .io_o_adder_17(my_fan_network_io_o_adder_17),
    .io_o_adder_18(my_fan_network_io_o_adder_18),
    .io_o_adder_19(my_fan_network_io_o_adder_19),
    .io_o_adder_20(my_fan_network_io_o_adder_20),
    .io_o_adder_21(my_fan_network_io_o_adder_21),
    .io_o_adder_22(my_fan_network_io_o_adder_22),
    .io_o_adder_23(my_fan_network_io_o_adder_23),
    .io_o_adder_24(my_fan_network_io_o_adder_24),
    .io_o_adder_25(my_fan_network_io_o_adder_25),
    .io_o_adder_26(my_fan_network_io_o_adder_26),
    .io_o_adder_27(my_fan_network_io_o_adder_27),
    .io_o_adder_28(my_fan_network_io_o_adder_28),
    .io_o_adder_29(my_fan_network_io_o_adder_29),
    .io_o_adder_30(my_fan_network_io_o_adder_30)
  );
  assign io_o_valid_0 = my_fan_network_io_o_valid_0; // @[FlexDPE.scala 80:16]
  assign io_o_valid_1 = my_fan_network_io_o_valid_1; // @[FlexDPE.scala 80:16]
  assign io_o_valid_2 = my_fan_network_io_o_valid_2; // @[FlexDPE.scala 80:16]
  assign io_o_valid_3 = my_fan_network_io_o_valid_3; // @[FlexDPE.scala 80:16]
  assign io_o_valid_4 = my_fan_network_io_o_valid_4; // @[FlexDPE.scala 80:16]
  assign io_o_valid_5 = my_fan_network_io_o_valid_5; // @[FlexDPE.scala 80:16]
  assign io_o_valid_6 = my_fan_network_io_o_valid_6; // @[FlexDPE.scala 80:16]
  assign io_o_valid_7 = my_fan_network_io_o_valid_7; // @[FlexDPE.scala 80:16]
  assign io_o_valid_8 = my_fan_network_io_o_valid_8; // @[FlexDPE.scala 80:16]
  assign io_o_valid_9 = my_fan_network_io_o_valid_9; // @[FlexDPE.scala 80:16]
  assign io_o_valid_10 = my_fan_network_io_o_valid_10; // @[FlexDPE.scala 80:16]
  assign io_o_valid_11 = my_fan_network_io_o_valid_11; // @[FlexDPE.scala 80:16]
  assign io_o_valid_12 = my_fan_network_io_o_valid_12; // @[FlexDPE.scala 80:16]
  assign io_o_valid_13 = my_fan_network_io_o_valid_13; // @[FlexDPE.scala 80:16]
  assign io_o_valid_14 = my_fan_network_io_o_valid_14; // @[FlexDPE.scala 80:16]
  assign io_o_valid_15 = my_fan_network_io_o_valid_15; // @[FlexDPE.scala 80:16]
  assign io_o_valid_16 = my_fan_network_io_o_valid_16; // @[FlexDPE.scala 80:16]
  assign io_o_valid_17 = my_fan_network_io_o_valid_17; // @[FlexDPE.scala 80:16]
  assign io_o_valid_18 = my_fan_network_io_o_valid_18; // @[FlexDPE.scala 80:16]
  assign io_o_valid_19 = my_fan_network_io_o_valid_19; // @[FlexDPE.scala 80:16]
  assign io_o_valid_20 = my_fan_network_io_o_valid_20; // @[FlexDPE.scala 80:16]
  assign io_o_valid_21 = my_fan_network_io_o_valid_21; // @[FlexDPE.scala 80:16]
  assign io_o_valid_22 = my_fan_network_io_o_valid_22; // @[FlexDPE.scala 80:16]
  assign io_o_valid_23 = my_fan_network_io_o_valid_23; // @[FlexDPE.scala 80:16]
  assign io_o_valid_24 = my_fan_network_io_o_valid_24; // @[FlexDPE.scala 80:16]
  assign io_o_valid_25 = my_fan_network_io_o_valid_25; // @[FlexDPE.scala 80:16]
  assign io_o_valid_26 = my_fan_network_io_o_valid_26; // @[FlexDPE.scala 80:16]
  assign io_o_valid_27 = my_fan_network_io_o_valid_27; // @[FlexDPE.scala 80:16]
  assign io_o_valid_28 = my_fan_network_io_o_valid_28; // @[FlexDPE.scala 80:16]
  assign io_o_valid_29 = my_fan_network_io_o_valid_29; // @[FlexDPE.scala 80:16]
  assign io_o_valid_30 = my_fan_network_io_o_valid_30; // @[FlexDPE.scala 80:16]
  assign io_o_valid_31 = my_fan_network_io_o_valid_31; // @[FlexDPE.scala 80:16]
  assign io_o_data_bus_0 = my_fan_network_io_o_data_bus_0; // @[FlexDPE.scala 81:19]
  assign io_o_data_bus_1 = my_fan_network_io_o_data_bus_1; // @[FlexDPE.scala 81:19]
  assign io_o_data_bus_2 = my_fan_network_io_o_data_bus_2; // @[FlexDPE.scala 81:19]
  assign io_o_data_bus_3 = my_fan_network_io_o_data_bus_3; // @[FlexDPE.scala 81:19]
  assign io_o_data_bus_4 = my_fan_network_io_o_data_bus_4; // @[FlexDPE.scala 81:19]
  assign io_o_data_bus_5 = my_fan_network_io_o_data_bus_5; // @[FlexDPE.scala 81:19]
  assign io_o_data_bus_6 = my_fan_network_io_o_data_bus_6; // @[FlexDPE.scala 81:19]
  assign io_o_data_bus_7 = my_fan_network_io_o_data_bus_7; // @[FlexDPE.scala 81:19]
  assign io_o_data_bus_8 = my_fan_network_io_o_data_bus_8; // @[FlexDPE.scala 81:19]
  assign io_o_data_bus_9 = my_fan_network_io_o_data_bus_9; // @[FlexDPE.scala 81:19]
  assign io_o_data_bus_10 = my_fan_network_io_o_data_bus_10; // @[FlexDPE.scala 81:19]
  assign io_o_data_bus_11 = my_fan_network_io_o_data_bus_11; // @[FlexDPE.scala 81:19]
  assign io_o_data_bus_12 = my_fan_network_io_o_data_bus_12; // @[FlexDPE.scala 81:19]
  assign io_o_data_bus_13 = my_fan_network_io_o_data_bus_13; // @[FlexDPE.scala 81:19]
  assign io_o_data_bus_14 = my_fan_network_io_o_data_bus_14; // @[FlexDPE.scala 81:19]
  assign io_o_data_bus_15 = my_fan_network_io_o_data_bus_15; // @[FlexDPE.scala 81:19]
  assign io_o_data_bus_16 = my_fan_network_io_o_data_bus_16; // @[FlexDPE.scala 81:19]
  assign io_o_data_bus_17 = my_fan_network_io_o_data_bus_17; // @[FlexDPE.scala 81:19]
  assign io_o_data_bus_18 = my_fan_network_io_o_data_bus_18; // @[FlexDPE.scala 81:19]
  assign io_o_data_bus_19 = my_fan_network_io_o_data_bus_19; // @[FlexDPE.scala 81:19]
  assign io_o_data_bus_20 = my_fan_network_io_o_data_bus_20; // @[FlexDPE.scala 81:19]
  assign io_o_data_bus_21 = my_fan_network_io_o_data_bus_21; // @[FlexDPE.scala 81:19]
  assign io_o_data_bus_22 = my_fan_network_io_o_data_bus_22; // @[FlexDPE.scala 81:19]
  assign io_o_data_bus_23 = my_fan_network_io_o_data_bus_23; // @[FlexDPE.scala 81:19]
  assign io_o_data_bus_24 = my_fan_network_io_o_data_bus_24; // @[FlexDPE.scala 81:19]
  assign io_o_data_bus_25 = my_fan_network_io_o_data_bus_25; // @[FlexDPE.scala 81:19]
  assign io_o_data_bus_26 = my_fan_network_io_o_data_bus_26; // @[FlexDPE.scala 81:19]
  assign io_o_data_bus_27 = my_fan_network_io_o_data_bus_27; // @[FlexDPE.scala 81:19]
  assign io_o_data_bus_28 = my_fan_network_io_o_data_bus_28; // @[FlexDPE.scala 81:19]
  assign io_o_data_bus_29 = my_fan_network_io_o_data_bus_29; // @[FlexDPE.scala 81:19]
  assign io_o_data_bus_30 = my_fan_network_io_o_data_bus_30; // @[FlexDPE.scala 81:19]
  assign io_o_data_bus_31 = my_fan_network_io_o_data_bus_31; // @[FlexDPE.scala 81:19]
  assign io_o_adder_0 = my_fan_network_io_o_adder_0; // @[FlexDPE.scala 82:16]
  assign io_o_adder_1 = my_fan_network_io_o_adder_1; // @[FlexDPE.scala 82:16]
  assign io_o_adder_2 = my_fan_network_io_o_adder_2; // @[FlexDPE.scala 82:16]
  assign io_o_adder_3 = my_fan_network_io_o_adder_3; // @[FlexDPE.scala 82:16]
  assign io_o_adder_4 = my_fan_network_io_o_adder_4; // @[FlexDPE.scala 82:16]
  assign io_o_adder_5 = my_fan_network_io_o_adder_5; // @[FlexDPE.scala 82:16]
  assign io_o_adder_6 = my_fan_network_io_o_adder_6; // @[FlexDPE.scala 82:16]
  assign io_o_adder_7 = my_fan_network_io_o_adder_7; // @[FlexDPE.scala 82:16]
  assign io_o_adder_8 = my_fan_network_io_o_adder_8; // @[FlexDPE.scala 82:16]
  assign io_o_adder_9 = my_fan_network_io_o_adder_9; // @[FlexDPE.scala 82:16]
  assign io_o_adder_10 = my_fan_network_io_o_adder_10; // @[FlexDPE.scala 82:16]
  assign io_o_adder_11 = my_fan_network_io_o_adder_11; // @[FlexDPE.scala 82:16]
  assign io_o_adder_12 = my_fan_network_io_o_adder_12; // @[FlexDPE.scala 82:16]
  assign io_o_adder_13 = my_fan_network_io_o_adder_13; // @[FlexDPE.scala 82:16]
  assign io_o_adder_14 = my_fan_network_io_o_adder_14; // @[FlexDPE.scala 82:16]
  assign io_o_adder_15 = my_fan_network_io_o_adder_15; // @[FlexDPE.scala 82:16]
  assign io_o_adder_16 = my_fan_network_io_o_adder_16; // @[FlexDPE.scala 82:16]
  assign io_o_adder_17 = my_fan_network_io_o_adder_17; // @[FlexDPE.scala 82:16]
  assign io_o_adder_18 = my_fan_network_io_o_adder_18; // @[FlexDPE.scala 82:16]
  assign io_o_adder_19 = my_fan_network_io_o_adder_19; // @[FlexDPE.scala 82:16]
  assign io_o_adder_20 = my_fan_network_io_o_adder_20; // @[FlexDPE.scala 82:16]
  assign io_o_adder_21 = my_fan_network_io_o_adder_21; // @[FlexDPE.scala 82:16]
  assign io_o_adder_22 = my_fan_network_io_o_adder_22; // @[FlexDPE.scala 82:16]
  assign io_o_adder_23 = my_fan_network_io_o_adder_23; // @[FlexDPE.scala 82:16]
  assign io_o_adder_24 = my_fan_network_io_o_adder_24; // @[FlexDPE.scala 82:16]
  assign io_o_adder_25 = my_fan_network_io_o_adder_25; // @[FlexDPE.scala 82:16]
  assign io_o_adder_26 = my_fan_network_io_o_adder_26; // @[FlexDPE.scala 82:16]
  assign io_o_adder_27 = my_fan_network_io_o_adder_27; // @[FlexDPE.scala 82:16]
  assign io_o_adder_28 = my_fan_network_io_o_adder_28; // @[FlexDPE.scala 82:16]
  assign io_o_adder_29 = my_fan_network_io_o_adder_29; // @[FlexDPE.scala 82:16]
  assign io_o_adder_30 = my_fan_network_io_o_adder_30; // @[FlexDPE.scala 82:16]
  assign my_controller_clock = clock;
  assign my_controller_reset = reset;
  assign my_Benes_clock = clock;
  assign my_Benes_reset = reset;
  assign buffer_mult_io_buffer2_0 = my_Benes_io_o_dist_bus2_0; // @[FlexDPE.scala 65:30]
  assign buffer_mult_io_buffer2_1 = my_Benes_io_o_dist_bus2_1; // @[FlexDPE.scala 65:30]
  assign buffer_mult_io_buffer2_2 = my_Benes_io_o_dist_bus2_2; // @[FlexDPE.scala 65:30]
  assign buffer_mult_io_buffer2_3 = my_Benes_io_o_dist_bus2_3; // @[FlexDPE.scala 65:30]
  assign buffer_mult_io_buffer2_4 = my_Benes_io_o_dist_bus2_4; // @[FlexDPE.scala 65:30]
  assign buffer_mult_io_buffer2_5 = my_Benes_io_o_dist_bus2_5; // @[FlexDPE.scala 65:30]
  assign buffer_mult_io_buffer2_6 = my_Benes_io_o_dist_bus2_6; // @[FlexDPE.scala 65:30]
  assign buffer_mult_io_buffer2_7 = my_Benes_io_o_dist_bus2_7; // @[FlexDPE.scala 65:30]
  assign buffer_mult_io_buffer2_8 = my_Benes_io_o_dist_bus2_8; // @[FlexDPE.scala 65:30]
  assign buffer_mult_io_buffer2_9 = my_Benes_io_o_dist_bus2_9; // @[FlexDPE.scala 65:30]
  assign buffer_mult_io_buffer2_10 = my_Benes_io_o_dist_bus2_10; // @[FlexDPE.scala 65:30]
  assign buffer_mult_io_buffer2_11 = my_Benes_io_o_dist_bus2_11; // @[FlexDPE.scala 65:30]
  assign buffer_mult_io_buffer2_12 = my_Benes_io_o_dist_bus2_12; // @[FlexDPE.scala 65:30]
  assign buffer_mult_io_buffer2_13 = my_Benes_io_o_dist_bus2_13; // @[FlexDPE.scala 65:30]
  assign buffer_mult_io_buffer2_14 = my_Benes_io_o_dist_bus2_14; // @[FlexDPE.scala 65:30]
  assign buffer_mult_io_buffer2_15 = my_Benes_io_o_dist_bus2_15; // @[FlexDPE.scala 65:30]
  assign buffer_mult_io_buffer2_16 = my_Benes_io_o_dist_bus2_16; // @[FlexDPE.scala 65:30]
  assign buffer_mult_io_buffer2_17 = my_Benes_io_o_dist_bus2_17; // @[FlexDPE.scala 65:30]
  assign buffer_mult_io_buffer2_18 = my_Benes_io_o_dist_bus2_18; // @[FlexDPE.scala 65:30]
  assign buffer_mult_io_buffer2_19 = my_Benes_io_o_dist_bus2_19; // @[FlexDPE.scala 65:30]
  assign buffer_mult_io_buffer2_20 = my_Benes_io_o_dist_bus2_20; // @[FlexDPE.scala 65:30]
  assign buffer_mult_io_buffer2_21 = my_Benes_io_o_dist_bus2_21; // @[FlexDPE.scala 65:30]
  assign buffer_mult_io_buffer2_22 = my_Benes_io_o_dist_bus2_22; // @[FlexDPE.scala 65:30]
  assign buffer_mult_io_buffer2_23 = my_Benes_io_o_dist_bus2_23; // @[FlexDPE.scala 65:30]
  assign buffer_mult_io_buffer2_24 = my_Benes_io_o_dist_bus2_24; // @[FlexDPE.scala 65:30]
  assign buffer_mult_io_buffer2_25 = my_Benes_io_o_dist_bus2_25; // @[FlexDPE.scala 65:30]
  assign buffer_mult_io_buffer2_26 = my_Benes_io_o_dist_bus2_26; // @[FlexDPE.scala 65:30]
  assign buffer_mult_io_buffer2_27 = my_Benes_io_o_dist_bus2_27; // @[FlexDPE.scala 65:30]
  assign buffer_mult_io_buffer2_28 = my_Benes_io_o_dist_bus2_28; // @[FlexDPE.scala 65:30]
  assign buffer_mult_io_buffer2_29 = my_Benes_io_o_dist_bus2_29; // @[FlexDPE.scala 65:30]
  assign buffer_mult_io_buffer2_30 = my_Benes_io_o_dist_bus2_30; // @[FlexDPE.scala 65:30]
  assign buffer_mult_io_buffer2_31 = my_Benes_io_o_dist_bus2_31; // @[FlexDPE.scala 65:30]
  assign my_fan_network_clock = clock;
  assign my_fan_network_reset = reset;
  assign my_fan_network_io_i_valid = my_controller_io_o_reduction_valid; // @[FlexDPE.scala 75:31]
  assign my_fan_network_io_i_data_bus_0 = {{1'd0}, r_mult_0}; // @[FlexDPE.scala 76:34]
  assign my_fan_network_io_i_data_bus_1 = {{1'd0}, r_mult_1}; // @[FlexDPE.scala 76:34]
  assign my_fan_network_io_i_data_bus_2 = {{1'd0}, r_mult_2}; // @[FlexDPE.scala 76:34]
  assign my_fan_network_io_i_data_bus_3 = {{1'd0}, r_mult_3}; // @[FlexDPE.scala 76:34]
  assign my_fan_network_io_i_data_bus_4 = {{1'd0}, r_mult_4}; // @[FlexDPE.scala 76:34]
  assign my_fan_network_io_i_data_bus_5 = {{1'd0}, r_mult_5}; // @[FlexDPE.scala 76:34]
  assign my_fan_network_io_i_data_bus_6 = {{1'd0}, r_mult_6}; // @[FlexDPE.scala 76:34]
  assign my_fan_network_io_i_data_bus_7 = {{1'd0}, r_mult_7}; // @[FlexDPE.scala 76:34]
  assign my_fan_network_io_i_data_bus_8 = {{1'd0}, r_mult_8}; // @[FlexDPE.scala 76:34]
  assign my_fan_network_io_i_data_bus_9 = {{1'd0}, r_mult_9}; // @[FlexDPE.scala 76:34]
  assign my_fan_network_io_i_data_bus_10 = {{1'd0}, r_mult_10}; // @[FlexDPE.scala 76:34]
  assign my_fan_network_io_i_data_bus_11 = {{1'd0}, r_mult_11}; // @[FlexDPE.scala 76:34]
  assign my_fan_network_io_i_data_bus_12 = {{1'd0}, r_mult_12}; // @[FlexDPE.scala 76:34]
  assign my_fan_network_io_i_data_bus_13 = {{1'd0}, r_mult_13}; // @[FlexDPE.scala 76:34]
  assign my_fan_network_io_i_data_bus_14 = {{1'd0}, r_mult_14}; // @[FlexDPE.scala 76:34]
  assign my_fan_network_io_i_data_bus_15 = {{1'd0}, r_mult_15}; // @[FlexDPE.scala 76:34]
  assign my_fan_network_io_i_data_bus_16 = {{1'd0}, r_mult_16}; // @[FlexDPE.scala 76:34]
  assign my_fan_network_io_i_data_bus_17 = {{1'd0}, r_mult_17}; // @[FlexDPE.scala 76:34]
  assign my_fan_network_io_i_data_bus_18 = {{1'd0}, r_mult_18}; // @[FlexDPE.scala 76:34]
  assign my_fan_network_io_i_data_bus_19 = {{1'd0}, r_mult_19}; // @[FlexDPE.scala 76:34]
  assign my_fan_network_io_i_data_bus_20 = {{1'd0}, r_mult_20}; // @[FlexDPE.scala 76:34]
  assign my_fan_network_io_i_data_bus_21 = {{1'd0}, r_mult_21}; // @[FlexDPE.scala 76:34]
  assign my_fan_network_io_i_data_bus_22 = {{1'd0}, r_mult_22}; // @[FlexDPE.scala 76:34]
  assign my_fan_network_io_i_data_bus_23 = {{1'd0}, r_mult_23}; // @[FlexDPE.scala 76:34]
  assign my_fan_network_io_i_data_bus_24 = {{1'd0}, r_mult_24}; // @[FlexDPE.scala 76:34]
  assign my_fan_network_io_i_data_bus_25 = {{1'd0}, r_mult_25}; // @[FlexDPE.scala 76:34]
  assign my_fan_network_io_i_data_bus_26 = {{1'd0}, r_mult_26}; // @[FlexDPE.scala 76:34]
  assign my_fan_network_io_i_data_bus_27 = {{1'd0}, r_mult_27}; // @[FlexDPE.scala 76:34]
  assign my_fan_network_io_i_data_bus_28 = {{1'd0}, r_mult_28}; // @[FlexDPE.scala 76:34]
  assign my_fan_network_io_i_data_bus_29 = {{1'd0}, r_mult_29}; // @[FlexDPE.scala 76:34]
  assign my_fan_network_io_i_data_bus_30 = {{1'd0}, r_mult_30}; // @[FlexDPE.scala 76:34]
  assign my_fan_network_io_i_data_bus_31 = {{1'd0}, r_mult_31}; // @[FlexDPE.scala 76:34]
  assign my_fan_network_io_i_add_en_bus_0 = my_controller_io_o_reduction_add_0; // @[FlexDPE.scala 77:36]
  assign my_fan_network_io_i_add_en_bus_1 = my_controller_io_o_reduction_add_1; // @[FlexDPE.scala 77:36]
  assign my_fan_network_io_i_add_en_bus_2 = my_controller_io_o_reduction_add_2; // @[FlexDPE.scala 77:36]
  assign my_fan_network_io_i_add_en_bus_3 = my_controller_io_o_reduction_add_3; // @[FlexDPE.scala 77:36]
  assign my_fan_network_io_i_add_en_bus_4 = my_controller_io_o_reduction_add_4; // @[FlexDPE.scala 77:36]
  assign my_fan_network_io_i_add_en_bus_5 = my_controller_io_o_reduction_add_5; // @[FlexDPE.scala 77:36]
  assign my_fan_network_io_i_add_en_bus_6 = my_controller_io_o_reduction_add_6; // @[FlexDPE.scala 77:36]
  assign my_fan_network_io_i_add_en_bus_7 = my_controller_io_o_reduction_add_7; // @[FlexDPE.scala 77:36]
  assign my_fan_network_io_i_add_en_bus_8 = my_controller_io_o_reduction_add_8; // @[FlexDPE.scala 77:36]
  assign my_fan_network_io_i_add_en_bus_9 = my_controller_io_o_reduction_add_9; // @[FlexDPE.scala 77:36]
  assign my_fan_network_io_i_add_en_bus_10 = my_controller_io_o_reduction_add_10; // @[FlexDPE.scala 77:36]
  assign my_fan_network_io_i_add_en_bus_11 = my_controller_io_o_reduction_add_11; // @[FlexDPE.scala 77:36]
  assign my_fan_network_io_i_add_en_bus_12 = my_controller_io_o_reduction_add_12; // @[FlexDPE.scala 77:36]
  assign my_fan_network_io_i_add_en_bus_13 = my_controller_io_o_reduction_add_13; // @[FlexDPE.scala 77:36]
  assign my_fan_network_io_i_add_en_bus_14 = my_controller_io_o_reduction_add_14; // @[FlexDPE.scala 77:36]
  assign my_fan_network_io_i_add_en_bus_15 = my_controller_io_o_reduction_add_15; // @[FlexDPE.scala 77:36]
  assign my_fan_network_io_i_add_en_bus_16 = my_controller_io_o_reduction_add_16; // @[FlexDPE.scala 77:36]
  assign my_fan_network_io_i_add_en_bus_17 = my_controller_io_o_reduction_add_17; // @[FlexDPE.scala 77:36]
  assign my_fan_network_io_i_add_en_bus_18 = my_controller_io_o_reduction_add_18; // @[FlexDPE.scala 77:36]
  assign my_fan_network_io_i_add_en_bus_19 = my_controller_io_o_reduction_add_19; // @[FlexDPE.scala 77:36]
  assign my_fan_network_io_i_add_en_bus_20 = my_controller_io_o_reduction_add_20; // @[FlexDPE.scala 77:36]
  assign my_fan_network_io_i_add_en_bus_21 = my_controller_io_o_reduction_add_21; // @[FlexDPE.scala 77:36]
  assign my_fan_network_io_i_add_en_bus_22 = my_controller_io_o_reduction_add_22; // @[FlexDPE.scala 77:36]
  assign my_fan_network_io_i_add_en_bus_23 = my_controller_io_o_reduction_add_23; // @[FlexDPE.scala 77:36]
  assign my_fan_network_io_i_add_en_bus_24 = my_controller_io_o_reduction_add_24; // @[FlexDPE.scala 77:36]
  assign my_fan_network_io_i_add_en_bus_25 = my_controller_io_o_reduction_add_25; // @[FlexDPE.scala 77:36]
  assign my_fan_network_io_i_add_en_bus_26 = my_controller_io_o_reduction_add_26; // @[FlexDPE.scala 77:36]
  assign my_fan_network_io_i_add_en_bus_27 = my_controller_io_o_reduction_add_27; // @[FlexDPE.scala 77:36]
  assign my_fan_network_io_i_add_en_bus_28 = my_controller_io_o_reduction_add_28; // @[FlexDPE.scala 77:36]
  assign my_fan_network_io_i_add_en_bus_29 = my_controller_io_o_reduction_add_29; // @[FlexDPE.scala 77:36]
  assign my_fan_network_io_i_add_en_bus_30 = my_controller_io_o_reduction_add_30; // @[FlexDPE.scala 77:36]
  assign my_fan_network_io_i_cmd_bus_0 = my_controller_io_o_reduction_cmd_0; // @[FlexDPE.scala 78:33]
  assign my_fan_network_io_i_cmd_bus_1 = my_controller_io_o_reduction_cmd_1; // @[FlexDPE.scala 78:33]
  assign my_fan_network_io_i_cmd_bus_2 = my_controller_io_o_reduction_cmd_2; // @[FlexDPE.scala 78:33]
  assign my_fan_network_io_i_cmd_bus_3 = my_controller_io_o_reduction_cmd_3; // @[FlexDPE.scala 78:33]
  assign my_fan_network_io_i_cmd_bus_4 = my_controller_io_o_reduction_cmd_4; // @[FlexDPE.scala 78:33]
  assign my_fan_network_io_i_cmd_bus_5 = my_controller_io_o_reduction_cmd_5; // @[FlexDPE.scala 78:33]
  assign my_fan_network_io_i_cmd_bus_6 = my_controller_io_o_reduction_cmd_6; // @[FlexDPE.scala 78:33]
  assign my_fan_network_io_i_cmd_bus_7 = my_controller_io_o_reduction_cmd_7; // @[FlexDPE.scala 78:33]
  assign my_fan_network_io_i_cmd_bus_8 = my_controller_io_o_reduction_cmd_8; // @[FlexDPE.scala 78:33]
  assign my_fan_network_io_i_cmd_bus_9 = my_controller_io_o_reduction_cmd_9; // @[FlexDPE.scala 78:33]
  assign my_fan_network_io_i_cmd_bus_10 = my_controller_io_o_reduction_cmd_10; // @[FlexDPE.scala 78:33]
  assign my_fan_network_io_i_cmd_bus_11 = my_controller_io_o_reduction_cmd_11; // @[FlexDPE.scala 78:33]
  assign my_fan_network_io_i_cmd_bus_12 = my_controller_io_o_reduction_cmd_12; // @[FlexDPE.scala 78:33]
  assign my_fan_network_io_i_cmd_bus_13 = my_controller_io_o_reduction_cmd_13; // @[FlexDPE.scala 78:33]
  assign my_fan_network_io_i_cmd_bus_14 = my_controller_io_o_reduction_cmd_14; // @[FlexDPE.scala 78:33]
  assign my_fan_network_io_i_cmd_bus_15 = my_controller_io_o_reduction_cmd_15; // @[FlexDPE.scala 78:33]
  assign my_fan_network_io_i_cmd_bus_16 = my_controller_io_o_reduction_cmd_16; // @[FlexDPE.scala 78:33]
  assign my_fan_network_io_i_cmd_bus_17 = my_controller_io_o_reduction_cmd_17; // @[FlexDPE.scala 78:33]
  assign my_fan_network_io_i_cmd_bus_18 = my_controller_io_o_reduction_cmd_18; // @[FlexDPE.scala 78:33]
  assign my_fan_network_io_i_cmd_bus_19 = my_controller_io_o_reduction_cmd_19; // @[FlexDPE.scala 78:33]
  assign my_fan_network_io_i_cmd_bus_20 = my_controller_io_o_reduction_cmd_20; // @[FlexDPE.scala 78:33]
  assign my_fan_network_io_i_cmd_bus_21 = my_controller_io_o_reduction_cmd_21; // @[FlexDPE.scala 78:33]
  assign my_fan_network_io_i_cmd_bus_22 = my_controller_io_o_reduction_cmd_22; // @[FlexDPE.scala 78:33]
  assign my_fan_network_io_i_cmd_bus_23 = my_controller_io_o_reduction_cmd_23; // @[FlexDPE.scala 78:33]
  assign my_fan_network_io_i_cmd_bus_24 = my_controller_io_o_reduction_cmd_24; // @[FlexDPE.scala 78:33]
  assign my_fan_network_io_i_cmd_bus_25 = my_controller_io_o_reduction_cmd_25; // @[FlexDPE.scala 78:33]
  assign my_fan_network_io_i_cmd_bus_26 = my_controller_io_o_reduction_cmd_26; // @[FlexDPE.scala 78:33]
  assign my_fan_network_io_i_cmd_bus_27 = my_controller_io_o_reduction_cmd_27; // @[FlexDPE.scala 78:33]
  assign my_fan_network_io_i_cmd_bus_28 = my_controller_io_o_reduction_cmd_28; // @[FlexDPE.scala 78:33]
  assign my_fan_network_io_i_cmd_bus_29 = my_controller_io_o_reduction_cmd_29; // @[FlexDPE.scala 78:33]
  assign my_fan_network_io_i_cmd_bus_30 = my_controller_io_o_reduction_cmd_30; // @[FlexDPE.scala 78:33]
  assign my_fan_network_io_i_sel_bus_0 = my_controller_io_o_reduction_sel_0; // @[FlexDPE.scala 79:33]
  assign my_fan_network_io_i_sel_bus_1 = my_controller_io_o_reduction_sel_1; // @[FlexDPE.scala 79:33]
  assign my_fan_network_io_i_sel_bus_2 = my_controller_io_o_reduction_sel_2; // @[FlexDPE.scala 79:33]
  assign my_fan_network_io_i_sel_bus_3 = my_controller_io_o_reduction_sel_3; // @[FlexDPE.scala 79:33]
  assign my_fan_network_io_i_sel_bus_4 = my_controller_io_o_reduction_sel_4; // @[FlexDPE.scala 79:33]
  assign my_fan_network_io_i_sel_bus_5 = my_controller_io_o_reduction_sel_5; // @[FlexDPE.scala 79:33]
  assign my_fan_network_io_i_sel_bus_6 = my_controller_io_o_reduction_sel_6; // @[FlexDPE.scala 79:33]
  assign my_fan_network_io_i_sel_bus_7 = my_controller_io_o_reduction_sel_7; // @[FlexDPE.scala 79:33]
  assign my_fan_network_io_i_sel_bus_8 = my_controller_io_o_reduction_sel_8; // @[FlexDPE.scala 79:33]
  assign my_fan_network_io_i_sel_bus_9 = my_controller_io_o_reduction_sel_9; // @[FlexDPE.scala 79:33]
  assign my_fan_network_io_i_sel_bus_10 = my_controller_io_o_reduction_sel_10; // @[FlexDPE.scala 79:33]
  assign my_fan_network_io_i_sel_bus_11 = my_controller_io_o_reduction_sel_11; // @[FlexDPE.scala 79:33]
  assign my_fan_network_io_i_sel_bus_12 = my_controller_io_o_reduction_sel_12; // @[FlexDPE.scala 79:33]
  assign my_fan_network_io_i_sel_bus_13 = my_controller_io_o_reduction_sel_13; // @[FlexDPE.scala 79:33]
  assign my_fan_network_io_i_sel_bus_14 = my_controller_io_o_reduction_sel_14; // @[FlexDPE.scala 79:33]
  assign my_fan_network_io_i_sel_bus_15 = my_controller_io_o_reduction_sel_15; // @[FlexDPE.scala 79:33]
  assign my_fan_network_io_i_sel_bus_16 = my_controller_io_o_reduction_sel_16; // @[FlexDPE.scala 79:33]
  assign my_fan_network_io_i_sel_bus_17 = my_controller_io_o_reduction_sel_17; // @[FlexDPE.scala 79:33]
  assign my_fan_network_io_i_sel_bus_18 = my_controller_io_o_reduction_sel_18; // @[FlexDPE.scala 79:33]
  assign my_fan_network_io_i_sel_bus_19 = my_controller_io_o_reduction_sel_19; // @[FlexDPE.scala 79:33]
  always @(posedge clock) begin
    if (reset) begin // @[FlexDPE.scala 24:26]
      r_mult_0 <= 31'h0; // @[FlexDPE.scala 24:26]
    end else begin
      r_mult_0 <= {{15'd0}, buffer_mult_io_out_0}; // @[FlexDPE.scala 67:14]
    end
    if (reset) begin // @[FlexDPE.scala 24:26]
      r_mult_1 <= 31'h0; // @[FlexDPE.scala 24:26]
    end else begin
      r_mult_1 <= {{15'd0}, buffer_mult_io_out_1}; // @[FlexDPE.scala 67:14]
    end
    if (reset) begin // @[FlexDPE.scala 24:26]
      r_mult_2 <= 31'h0; // @[FlexDPE.scala 24:26]
    end else begin
      r_mult_2 <= {{15'd0}, buffer_mult_io_out_2}; // @[FlexDPE.scala 67:14]
    end
    if (reset) begin // @[FlexDPE.scala 24:26]
      r_mult_3 <= 31'h0; // @[FlexDPE.scala 24:26]
    end else begin
      r_mult_3 <= {{15'd0}, buffer_mult_io_out_3}; // @[FlexDPE.scala 67:14]
    end
    if (reset) begin // @[FlexDPE.scala 24:26]
      r_mult_4 <= 31'h0; // @[FlexDPE.scala 24:26]
    end else begin
      r_mult_4 <= {{15'd0}, buffer_mult_io_out_4}; // @[FlexDPE.scala 67:14]
    end
    if (reset) begin // @[FlexDPE.scala 24:26]
      r_mult_5 <= 31'h0; // @[FlexDPE.scala 24:26]
    end else begin
      r_mult_5 <= {{15'd0}, buffer_mult_io_out_5}; // @[FlexDPE.scala 67:14]
    end
    if (reset) begin // @[FlexDPE.scala 24:26]
      r_mult_6 <= 31'h0; // @[FlexDPE.scala 24:26]
    end else begin
      r_mult_6 <= {{15'd0}, buffer_mult_io_out_6}; // @[FlexDPE.scala 67:14]
    end
    if (reset) begin // @[FlexDPE.scala 24:26]
      r_mult_7 <= 31'h0; // @[FlexDPE.scala 24:26]
    end else begin
      r_mult_7 <= {{15'd0}, buffer_mult_io_out_7}; // @[FlexDPE.scala 67:14]
    end
    if (reset) begin // @[FlexDPE.scala 24:26]
      r_mult_8 <= 31'h0; // @[FlexDPE.scala 24:26]
    end else begin
      r_mult_8 <= {{15'd0}, buffer_mult_io_out_8}; // @[FlexDPE.scala 67:14]
    end
    if (reset) begin // @[FlexDPE.scala 24:26]
      r_mult_9 <= 31'h0; // @[FlexDPE.scala 24:26]
    end else begin
      r_mult_9 <= {{15'd0}, buffer_mult_io_out_9}; // @[FlexDPE.scala 67:14]
    end
    if (reset) begin // @[FlexDPE.scala 24:26]
      r_mult_10 <= 31'h0; // @[FlexDPE.scala 24:26]
    end else begin
      r_mult_10 <= {{15'd0}, buffer_mult_io_out_10}; // @[FlexDPE.scala 67:14]
    end
    if (reset) begin // @[FlexDPE.scala 24:26]
      r_mult_11 <= 31'h0; // @[FlexDPE.scala 24:26]
    end else begin
      r_mult_11 <= {{15'd0}, buffer_mult_io_out_11}; // @[FlexDPE.scala 67:14]
    end
    if (reset) begin // @[FlexDPE.scala 24:26]
      r_mult_12 <= 31'h0; // @[FlexDPE.scala 24:26]
    end else begin
      r_mult_12 <= {{15'd0}, buffer_mult_io_out_12}; // @[FlexDPE.scala 67:14]
    end
    if (reset) begin // @[FlexDPE.scala 24:26]
      r_mult_13 <= 31'h0; // @[FlexDPE.scala 24:26]
    end else begin
      r_mult_13 <= {{15'd0}, buffer_mult_io_out_13}; // @[FlexDPE.scala 67:14]
    end
    if (reset) begin // @[FlexDPE.scala 24:26]
      r_mult_14 <= 31'h0; // @[FlexDPE.scala 24:26]
    end else begin
      r_mult_14 <= {{15'd0}, buffer_mult_io_out_14}; // @[FlexDPE.scala 67:14]
    end
    if (reset) begin // @[FlexDPE.scala 24:26]
      r_mult_15 <= 31'h0; // @[FlexDPE.scala 24:26]
    end else begin
      r_mult_15 <= {{15'd0}, buffer_mult_io_out_15}; // @[FlexDPE.scala 67:14]
    end
    if (reset) begin // @[FlexDPE.scala 24:26]
      r_mult_16 <= 31'h0; // @[FlexDPE.scala 24:26]
    end else begin
      r_mult_16 <= {{15'd0}, buffer_mult_io_out_16}; // @[FlexDPE.scala 67:14]
    end
    if (reset) begin // @[FlexDPE.scala 24:26]
      r_mult_17 <= 31'h0; // @[FlexDPE.scala 24:26]
    end else begin
      r_mult_17 <= {{15'd0}, buffer_mult_io_out_17}; // @[FlexDPE.scala 67:14]
    end
    if (reset) begin // @[FlexDPE.scala 24:26]
      r_mult_18 <= 31'h0; // @[FlexDPE.scala 24:26]
    end else begin
      r_mult_18 <= {{15'd0}, buffer_mult_io_out_18}; // @[FlexDPE.scala 67:14]
    end
    if (reset) begin // @[FlexDPE.scala 24:26]
      r_mult_19 <= 31'h0; // @[FlexDPE.scala 24:26]
    end else begin
      r_mult_19 <= {{15'd0}, buffer_mult_io_out_19}; // @[FlexDPE.scala 67:14]
    end
    if (reset) begin // @[FlexDPE.scala 24:26]
      r_mult_20 <= 31'h0; // @[FlexDPE.scala 24:26]
    end else begin
      r_mult_20 <= {{15'd0}, buffer_mult_io_out_20}; // @[FlexDPE.scala 67:14]
    end
    if (reset) begin // @[FlexDPE.scala 24:26]
      r_mult_21 <= 31'h0; // @[FlexDPE.scala 24:26]
    end else begin
      r_mult_21 <= {{15'd0}, buffer_mult_io_out_21}; // @[FlexDPE.scala 67:14]
    end
    if (reset) begin // @[FlexDPE.scala 24:26]
      r_mult_22 <= 31'h0; // @[FlexDPE.scala 24:26]
    end else begin
      r_mult_22 <= {{15'd0}, buffer_mult_io_out_22}; // @[FlexDPE.scala 67:14]
    end
    if (reset) begin // @[FlexDPE.scala 24:26]
      r_mult_23 <= 31'h0; // @[FlexDPE.scala 24:26]
    end else begin
      r_mult_23 <= {{15'd0}, buffer_mult_io_out_23}; // @[FlexDPE.scala 67:14]
    end
    if (reset) begin // @[FlexDPE.scala 24:26]
      r_mult_24 <= 31'h0; // @[FlexDPE.scala 24:26]
    end else begin
      r_mult_24 <= {{15'd0}, buffer_mult_io_out_24}; // @[FlexDPE.scala 67:14]
    end
    if (reset) begin // @[FlexDPE.scala 24:26]
      r_mult_25 <= 31'h0; // @[FlexDPE.scala 24:26]
    end else begin
      r_mult_25 <= {{15'd0}, buffer_mult_io_out_25}; // @[FlexDPE.scala 67:14]
    end
    if (reset) begin // @[FlexDPE.scala 24:26]
      r_mult_26 <= 31'h0; // @[FlexDPE.scala 24:26]
    end else begin
      r_mult_26 <= {{15'd0}, buffer_mult_io_out_26}; // @[FlexDPE.scala 67:14]
    end
    if (reset) begin // @[FlexDPE.scala 24:26]
      r_mult_27 <= 31'h0; // @[FlexDPE.scala 24:26]
    end else begin
      r_mult_27 <= {{15'd0}, buffer_mult_io_out_27}; // @[FlexDPE.scala 67:14]
    end
    if (reset) begin // @[FlexDPE.scala 24:26]
      r_mult_28 <= 31'h0; // @[FlexDPE.scala 24:26]
    end else begin
      r_mult_28 <= {{15'd0}, buffer_mult_io_out_28}; // @[FlexDPE.scala 67:14]
    end
    if (reset) begin // @[FlexDPE.scala 24:26]
      r_mult_29 <= 31'h0; // @[FlexDPE.scala 24:26]
    end else begin
      r_mult_29 <= {{15'd0}, buffer_mult_io_out_29}; // @[FlexDPE.scala 67:14]
    end
    if (reset) begin // @[FlexDPE.scala 24:26]
      r_mult_30 <= 31'h0; // @[FlexDPE.scala 24:26]
    end else begin
      r_mult_30 <= {{15'd0}, buffer_mult_io_out_30}; // @[FlexDPE.scala 67:14]
    end
    if (reset) begin // @[FlexDPE.scala 24:26]
      r_mult_31 <= 31'h0; // @[FlexDPE.scala 24:26]
    end else begin
      r_mult_31 <= {{15'd0}, buffer_mult_io_out_31}; // @[FlexDPE.scala 67:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_mult_0 = _RAND_0[30:0];
  _RAND_1 = {1{`RANDOM}};
  r_mult_1 = _RAND_1[30:0];
  _RAND_2 = {1{`RANDOM}};
  r_mult_2 = _RAND_2[30:0];
  _RAND_3 = {1{`RANDOM}};
  r_mult_3 = _RAND_3[30:0];
  _RAND_4 = {1{`RANDOM}};
  r_mult_4 = _RAND_4[30:0];
  _RAND_5 = {1{`RANDOM}};
  r_mult_5 = _RAND_5[30:0];
  _RAND_6 = {1{`RANDOM}};
  r_mult_6 = _RAND_6[30:0];
  _RAND_7 = {1{`RANDOM}};
  r_mult_7 = _RAND_7[30:0];
  _RAND_8 = {1{`RANDOM}};
  r_mult_8 = _RAND_8[30:0];
  _RAND_9 = {1{`RANDOM}};
  r_mult_9 = _RAND_9[30:0];
  _RAND_10 = {1{`RANDOM}};
  r_mult_10 = _RAND_10[30:0];
  _RAND_11 = {1{`RANDOM}};
  r_mult_11 = _RAND_11[30:0];
  _RAND_12 = {1{`RANDOM}};
  r_mult_12 = _RAND_12[30:0];
  _RAND_13 = {1{`RANDOM}};
  r_mult_13 = _RAND_13[30:0];
  _RAND_14 = {1{`RANDOM}};
  r_mult_14 = _RAND_14[30:0];
  _RAND_15 = {1{`RANDOM}};
  r_mult_15 = _RAND_15[30:0];
  _RAND_16 = {1{`RANDOM}};
  r_mult_16 = _RAND_16[30:0];
  _RAND_17 = {1{`RANDOM}};
  r_mult_17 = _RAND_17[30:0];
  _RAND_18 = {1{`RANDOM}};
  r_mult_18 = _RAND_18[30:0];
  _RAND_19 = {1{`RANDOM}};
  r_mult_19 = _RAND_19[30:0];
  _RAND_20 = {1{`RANDOM}};
  r_mult_20 = _RAND_20[30:0];
  _RAND_21 = {1{`RANDOM}};
  r_mult_21 = _RAND_21[30:0];
  _RAND_22 = {1{`RANDOM}};
  r_mult_22 = _RAND_22[30:0];
  _RAND_23 = {1{`RANDOM}};
  r_mult_23 = _RAND_23[30:0];
  _RAND_24 = {1{`RANDOM}};
  r_mult_24 = _RAND_24[30:0];
  _RAND_25 = {1{`RANDOM}};
  r_mult_25 = _RAND_25[30:0];
  _RAND_26 = {1{`RANDOM}};
  r_mult_26 = _RAND_26[30:0];
  _RAND_27 = {1{`RANDOM}};
  r_mult_27 = _RAND_27[30:0];
  _RAND_28 = {1{`RANDOM}};
  r_mult_28 = _RAND_28[30:0];
  _RAND_29 = {1{`RANDOM}};
  r_mult_29 = _RAND_29[30:0];
  _RAND_30 = {1{`RANDOM}};
  r_mult_30 = _RAND_30[30:0];
  _RAND_31 = {1{`RANDOM}};
  r_mult_31 = _RAND_31[30:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FDPEWrapper(
  input         clock,
  input         reset,
  output        io_o_valid_0,
  output        io_o_valid_1,
  output        io_o_valid_2,
  output        io_o_valid_3,
  output        io_o_valid_4,
  output        io_o_valid_5,
  output        io_o_valid_6,
  output        io_o_valid_7,
  output        io_o_valid_8,
  output        io_o_valid_9,
  output        io_o_valid_10,
  output        io_o_valid_11,
  output        io_o_valid_12,
  output        io_o_valid_13,
  output        io_o_valid_14,
  output        io_o_valid_15,
  output        io_o_valid_16,
  output        io_o_valid_17,
  output        io_o_valid_18,
  output        io_o_valid_19,
  output        io_o_valid_20,
  output        io_o_valid_21,
  output        io_o_valid_22,
  output        io_o_valid_23,
  output        io_o_valid_24,
  output        io_o_valid_25,
  output        io_o_valid_26,
  output        io_o_valid_27,
  output        io_o_valid_28,
  output        io_o_valid_29,
  output        io_o_valid_30,
  output        io_o_valid_31,
  output [15:0] io_o_data_bus_0,
  output [15:0] io_o_data_bus_1,
  output [15:0] io_o_data_bus_2,
  output [15:0] io_o_data_bus_3,
  output [15:0] io_o_data_bus_4,
  output [15:0] io_o_data_bus_5,
  output [15:0] io_o_data_bus_6,
  output [15:0] io_o_data_bus_7,
  output [15:0] io_o_data_bus_8,
  output [15:0] io_o_data_bus_9,
  output [15:0] io_o_data_bus_10,
  output [15:0] io_o_data_bus_11,
  output [15:0] io_o_data_bus_12,
  output [15:0] io_o_data_bus_13,
  output [15:0] io_o_data_bus_14,
  output [15:0] io_o_data_bus_15,
  output [15:0] io_o_data_bus_16,
  output [15:0] io_o_data_bus_17,
  output [15:0] io_o_data_bus_18,
  output [15:0] io_o_data_bus_19,
  output [15:0] io_o_data_bus_20,
  output [15:0] io_o_data_bus_21,
  output [15:0] io_o_data_bus_22,
  output [15:0] io_o_data_bus_23,
  output [15:0] io_o_data_bus_24,
  output [15:0] io_o_data_bus_25,
  output [15:0] io_o_data_bus_26,
  output [15:0] io_o_data_bus_27,
  output [15:0] io_o_data_bus_28,
  output [15:0] io_o_data_bus_29,
  output [15:0] io_o_data_bus_30,
  output [15:0] io_o_data_bus_31,
  output [15:0] io_o_adder_0,
  output [15:0] io_o_adder_1,
  output [15:0] io_o_adder_2,
  output [15:0] io_o_adder_3,
  output [15:0] io_o_adder_4,
  output [15:0] io_o_adder_5,
  output [15:0] io_o_adder_6,
  output [15:0] io_o_adder_7,
  output [15:0] io_o_adder_8,
  output [15:0] io_o_adder_9,
  output [15:0] io_o_adder_10,
  output [15:0] io_o_adder_11,
  output [15:0] io_o_adder_12,
  output [15:0] io_o_adder_13,
  output [15:0] io_o_adder_14,
  output [15:0] io_o_adder_15,
  output [15:0] io_o_adder_16,
  output [15:0] io_o_adder_17,
  output [15:0] io_o_adder_18,
  output [15:0] io_o_adder_19,
  output [15:0] io_o_adder_20,
  output [15:0] io_o_adder_21,
  output [15:0] io_o_adder_22,
  output [15:0] io_o_adder_23,
  output [15:0] io_o_adder_24,
  output [15:0] io_o_adder_25,
  output [15:0] io_o_adder_26,
  output [15:0] io_o_adder_27,
  output [15:0] io_o_adder_28,
  output [15:0] io_o_adder_29,
  output [15:0] io_o_adder_30,
  output [15:0] io_o_adder_31
);
  wire  FDPE_clock; // @[FDPEWrapper.scala 15:22]
  wire  FDPE_reset; // @[FDPEWrapper.scala 15:22]
  wire  FDPE_io_o_valid_0; // @[FDPEWrapper.scala 15:22]
  wire  FDPE_io_o_valid_1; // @[FDPEWrapper.scala 15:22]
  wire  FDPE_io_o_valid_2; // @[FDPEWrapper.scala 15:22]
  wire  FDPE_io_o_valid_3; // @[FDPEWrapper.scala 15:22]
  wire  FDPE_io_o_valid_4; // @[FDPEWrapper.scala 15:22]
  wire  FDPE_io_o_valid_5; // @[FDPEWrapper.scala 15:22]
  wire  FDPE_io_o_valid_6; // @[FDPEWrapper.scala 15:22]
  wire  FDPE_io_o_valid_7; // @[FDPEWrapper.scala 15:22]
  wire  FDPE_io_o_valid_8; // @[FDPEWrapper.scala 15:22]
  wire  FDPE_io_o_valid_9; // @[FDPEWrapper.scala 15:22]
  wire  FDPE_io_o_valid_10; // @[FDPEWrapper.scala 15:22]
  wire  FDPE_io_o_valid_11; // @[FDPEWrapper.scala 15:22]
  wire  FDPE_io_o_valid_12; // @[FDPEWrapper.scala 15:22]
  wire  FDPE_io_o_valid_13; // @[FDPEWrapper.scala 15:22]
  wire  FDPE_io_o_valid_14; // @[FDPEWrapper.scala 15:22]
  wire  FDPE_io_o_valid_15; // @[FDPEWrapper.scala 15:22]
  wire  FDPE_io_o_valid_16; // @[FDPEWrapper.scala 15:22]
  wire  FDPE_io_o_valid_17; // @[FDPEWrapper.scala 15:22]
  wire  FDPE_io_o_valid_18; // @[FDPEWrapper.scala 15:22]
  wire  FDPE_io_o_valid_19; // @[FDPEWrapper.scala 15:22]
  wire  FDPE_io_o_valid_20; // @[FDPEWrapper.scala 15:22]
  wire  FDPE_io_o_valid_21; // @[FDPEWrapper.scala 15:22]
  wire  FDPE_io_o_valid_22; // @[FDPEWrapper.scala 15:22]
  wire  FDPE_io_o_valid_23; // @[FDPEWrapper.scala 15:22]
  wire  FDPE_io_o_valid_24; // @[FDPEWrapper.scala 15:22]
  wire  FDPE_io_o_valid_25; // @[FDPEWrapper.scala 15:22]
  wire  FDPE_io_o_valid_26; // @[FDPEWrapper.scala 15:22]
  wire  FDPE_io_o_valid_27; // @[FDPEWrapper.scala 15:22]
  wire  FDPE_io_o_valid_28; // @[FDPEWrapper.scala 15:22]
  wire  FDPE_io_o_valid_29; // @[FDPEWrapper.scala 15:22]
  wire  FDPE_io_o_valid_30; // @[FDPEWrapper.scala 15:22]
  wire  FDPE_io_o_valid_31; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_data_bus_0; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_data_bus_1; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_data_bus_2; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_data_bus_3; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_data_bus_4; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_data_bus_5; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_data_bus_6; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_data_bus_7; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_data_bus_8; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_data_bus_9; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_data_bus_10; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_data_bus_11; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_data_bus_12; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_data_bus_13; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_data_bus_14; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_data_bus_15; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_data_bus_16; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_data_bus_17; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_data_bus_18; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_data_bus_19; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_data_bus_20; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_data_bus_21; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_data_bus_22; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_data_bus_23; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_data_bus_24; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_data_bus_25; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_data_bus_26; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_data_bus_27; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_data_bus_28; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_data_bus_29; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_data_bus_30; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_data_bus_31; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_adder_0; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_adder_1; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_adder_2; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_adder_3; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_adder_4; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_adder_5; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_adder_6; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_adder_7; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_adder_8; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_adder_9; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_adder_10; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_adder_11; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_adder_12; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_adder_13; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_adder_14; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_adder_15; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_adder_16; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_adder_17; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_adder_18; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_adder_19; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_adder_20; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_adder_21; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_adder_22; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_adder_23; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_adder_24; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_adder_25; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_adder_26; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_adder_27; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_adder_28; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_adder_29; // @[FDPEWrapper.scala 15:22]
  wire [31:0] FDPE_io_o_adder_30; // @[FDPEWrapper.scala 15:22]
  flexdpecom2 FDPE ( // @[FDPEWrapper.scala 15:22]
    .clock(FDPE_clock),
    .reset(FDPE_reset),
    .io_o_valid_0(FDPE_io_o_valid_0),
    .io_o_valid_1(FDPE_io_o_valid_1),
    .io_o_valid_2(FDPE_io_o_valid_2),
    .io_o_valid_3(FDPE_io_o_valid_3),
    .io_o_valid_4(FDPE_io_o_valid_4),
    .io_o_valid_5(FDPE_io_o_valid_5),
    .io_o_valid_6(FDPE_io_o_valid_6),
    .io_o_valid_7(FDPE_io_o_valid_7),
    .io_o_valid_8(FDPE_io_o_valid_8),
    .io_o_valid_9(FDPE_io_o_valid_9),
    .io_o_valid_10(FDPE_io_o_valid_10),
    .io_o_valid_11(FDPE_io_o_valid_11),
    .io_o_valid_12(FDPE_io_o_valid_12),
    .io_o_valid_13(FDPE_io_o_valid_13),
    .io_o_valid_14(FDPE_io_o_valid_14),
    .io_o_valid_15(FDPE_io_o_valid_15),
    .io_o_valid_16(FDPE_io_o_valid_16),
    .io_o_valid_17(FDPE_io_o_valid_17),
    .io_o_valid_18(FDPE_io_o_valid_18),
    .io_o_valid_19(FDPE_io_o_valid_19),
    .io_o_valid_20(FDPE_io_o_valid_20),
    .io_o_valid_21(FDPE_io_o_valid_21),
    .io_o_valid_22(FDPE_io_o_valid_22),
    .io_o_valid_23(FDPE_io_o_valid_23),
    .io_o_valid_24(FDPE_io_o_valid_24),
    .io_o_valid_25(FDPE_io_o_valid_25),
    .io_o_valid_26(FDPE_io_o_valid_26),
    .io_o_valid_27(FDPE_io_o_valid_27),
    .io_o_valid_28(FDPE_io_o_valid_28),
    .io_o_valid_29(FDPE_io_o_valid_29),
    .io_o_valid_30(FDPE_io_o_valid_30),
    .io_o_valid_31(FDPE_io_o_valid_31),
    .io_o_data_bus_0(FDPE_io_o_data_bus_0),
    .io_o_data_bus_1(FDPE_io_o_data_bus_1),
    .io_o_data_bus_2(FDPE_io_o_data_bus_2),
    .io_o_data_bus_3(FDPE_io_o_data_bus_3),
    .io_o_data_bus_4(FDPE_io_o_data_bus_4),
    .io_o_data_bus_5(FDPE_io_o_data_bus_5),
    .io_o_data_bus_6(FDPE_io_o_data_bus_6),
    .io_o_data_bus_7(FDPE_io_o_data_bus_7),
    .io_o_data_bus_8(FDPE_io_o_data_bus_8),
    .io_o_data_bus_9(FDPE_io_o_data_bus_9),
    .io_o_data_bus_10(FDPE_io_o_data_bus_10),
    .io_o_data_bus_11(FDPE_io_o_data_bus_11),
    .io_o_data_bus_12(FDPE_io_o_data_bus_12),
    .io_o_data_bus_13(FDPE_io_o_data_bus_13),
    .io_o_data_bus_14(FDPE_io_o_data_bus_14),
    .io_o_data_bus_15(FDPE_io_o_data_bus_15),
    .io_o_data_bus_16(FDPE_io_o_data_bus_16),
    .io_o_data_bus_17(FDPE_io_o_data_bus_17),
    .io_o_data_bus_18(FDPE_io_o_data_bus_18),
    .io_o_data_bus_19(FDPE_io_o_data_bus_19),
    .io_o_data_bus_20(FDPE_io_o_data_bus_20),
    .io_o_data_bus_21(FDPE_io_o_data_bus_21),
    .io_o_data_bus_22(FDPE_io_o_data_bus_22),
    .io_o_data_bus_23(FDPE_io_o_data_bus_23),
    .io_o_data_bus_24(FDPE_io_o_data_bus_24),
    .io_o_data_bus_25(FDPE_io_o_data_bus_25),
    .io_o_data_bus_26(FDPE_io_o_data_bus_26),
    .io_o_data_bus_27(FDPE_io_o_data_bus_27),
    .io_o_data_bus_28(FDPE_io_o_data_bus_28),
    .io_o_data_bus_29(FDPE_io_o_data_bus_29),
    .io_o_data_bus_30(FDPE_io_o_data_bus_30),
    .io_o_data_bus_31(FDPE_io_o_data_bus_31),
    .io_o_adder_0(FDPE_io_o_adder_0),
    .io_o_adder_1(FDPE_io_o_adder_1),
    .io_o_adder_2(FDPE_io_o_adder_2),
    .io_o_adder_3(FDPE_io_o_adder_3),
    .io_o_adder_4(FDPE_io_o_adder_4),
    .io_o_adder_5(FDPE_io_o_adder_5),
    .io_o_adder_6(FDPE_io_o_adder_6),
    .io_o_adder_7(FDPE_io_o_adder_7),
    .io_o_adder_8(FDPE_io_o_adder_8),
    .io_o_adder_9(FDPE_io_o_adder_9),
    .io_o_adder_10(FDPE_io_o_adder_10),
    .io_o_adder_11(FDPE_io_o_adder_11),
    .io_o_adder_12(FDPE_io_o_adder_12),
    .io_o_adder_13(FDPE_io_o_adder_13),
    .io_o_adder_14(FDPE_io_o_adder_14),
    .io_o_adder_15(FDPE_io_o_adder_15),
    .io_o_adder_16(FDPE_io_o_adder_16),
    .io_o_adder_17(FDPE_io_o_adder_17),
    .io_o_adder_18(FDPE_io_o_adder_18),
    .io_o_adder_19(FDPE_io_o_adder_19),
    .io_o_adder_20(FDPE_io_o_adder_20),
    .io_o_adder_21(FDPE_io_o_adder_21),
    .io_o_adder_22(FDPE_io_o_adder_22),
    .io_o_adder_23(FDPE_io_o_adder_23),
    .io_o_adder_24(FDPE_io_o_adder_24),
    .io_o_adder_25(FDPE_io_o_adder_25),
    .io_o_adder_26(FDPE_io_o_adder_26),
    .io_o_adder_27(FDPE_io_o_adder_27),
    .io_o_adder_28(FDPE_io_o_adder_28),
    .io_o_adder_29(FDPE_io_o_adder_29),
    .io_o_adder_30(FDPE_io_o_adder_30)
  );
  assign io_o_valid_0 = FDPE_io_o_valid_0; // @[FDPEWrapper.scala 45:16]
  assign io_o_valid_1 = FDPE_io_o_valid_1; // @[FDPEWrapper.scala 45:16]
  assign io_o_valid_2 = FDPE_io_o_valid_2; // @[FDPEWrapper.scala 45:16]
  assign io_o_valid_3 = FDPE_io_o_valid_3; // @[FDPEWrapper.scala 45:16]
  assign io_o_valid_4 = FDPE_io_o_valid_4; // @[FDPEWrapper.scala 45:16]
  assign io_o_valid_5 = FDPE_io_o_valid_5; // @[FDPEWrapper.scala 45:16]
  assign io_o_valid_6 = FDPE_io_o_valid_6; // @[FDPEWrapper.scala 45:16]
  assign io_o_valid_7 = FDPE_io_o_valid_7; // @[FDPEWrapper.scala 45:16]
  assign io_o_valid_8 = FDPE_io_o_valid_8; // @[FDPEWrapper.scala 45:16]
  assign io_o_valid_9 = FDPE_io_o_valid_9; // @[FDPEWrapper.scala 45:16]
  assign io_o_valid_10 = FDPE_io_o_valid_10; // @[FDPEWrapper.scala 45:16]
  assign io_o_valid_11 = FDPE_io_o_valid_11; // @[FDPEWrapper.scala 45:16]
  assign io_o_valid_12 = FDPE_io_o_valid_12; // @[FDPEWrapper.scala 45:16]
  assign io_o_valid_13 = FDPE_io_o_valid_13; // @[FDPEWrapper.scala 45:16]
  assign io_o_valid_14 = FDPE_io_o_valid_14; // @[FDPEWrapper.scala 45:16]
  assign io_o_valid_15 = FDPE_io_o_valid_15; // @[FDPEWrapper.scala 45:16]
  assign io_o_valid_16 = FDPE_io_o_valid_16; // @[FDPEWrapper.scala 45:16]
  assign io_o_valid_17 = FDPE_io_o_valid_17; // @[FDPEWrapper.scala 45:16]
  assign io_o_valid_18 = FDPE_io_o_valid_18; // @[FDPEWrapper.scala 45:16]
  assign io_o_valid_19 = FDPE_io_o_valid_19; // @[FDPEWrapper.scala 45:16]
  assign io_o_valid_20 = FDPE_io_o_valid_20; // @[FDPEWrapper.scala 45:16]
  assign io_o_valid_21 = FDPE_io_o_valid_21; // @[FDPEWrapper.scala 45:16]
  assign io_o_valid_22 = FDPE_io_o_valid_22; // @[FDPEWrapper.scala 45:16]
  assign io_o_valid_23 = FDPE_io_o_valid_23; // @[FDPEWrapper.scala 45:16]
  assign io_o_valid_24 = FDPE_io_o_valid_24; // @[FDPEWrapper.scala 45:16]
  assign io_o_valid_25 = FDPE_io_o_valid_25; // @[FDPEWrapper.scala 45:16]
  assign io_o_valid_26 = FDPE_io_o_valid_26; // @[FDPEWrapper.scala 45:16]
  assign io_o_valid_27 = FDPE_io_o_valid_27; // @[FDPEWrapper.scala 45:16]
  assign io_o_valid_28 = FDPE_io_o_valid_28; // @[FDPEWrapper.scala 45:16]
  assign io_o_valid_29 = FDPE_io_o_valid_29; // @[FDPEWrapper.scala 45:16]
  assign io_o_valid_30 = FDPE_io_o_valid_30; // @[FDPEWrapper.scala 45:16]
  assign io_o_valid_31 = FDPE_io_o_valid_31; // @[FDPEWrapper.scala 45:16]
  assign io_o_data_bus_0 = FDPE_io_o_data_bus_0[15:0]; // @[FDPEWrapper.scala 46:19]
  assign io_o_data_bus_1 = FDPE_io_o_data_bus_1[15:0]; // @[FDPEWrapper.scala 46:19]
  assign io_o_data_bus_2 = FDPE_io_o_data_bus_2[15:0]; // @[FDPEWrapper.scala 46:19]
  assign io_o_data_bus_3 = FDPE_io_o_data_bus_3[15:0]; // @[FDPEWrapper.scala 46:19]
  assign io_o_data_bus_4 = FDPE_io_o_data_bus_4[15:0]; // @[FDPEWrapper.scala 46:19]
  assign io_o_data_bus_5 = FDPE_io_o_data_bus_5[15:0]; // @[FDPEWrapper.scala 46:19]
  assign io_o_data_bus_6 = FDPE_io_o_data_bus_6[15:0]; // @[FDPEWrapper.scala 46:19]
  assign io_o_data_bus_7 = FDPE_io_o_data_bus_7[15:0]; // @[FDPEWrapper.scala 46:19]
  assign io_o_data_bus_8 = FDPE_io_o_data_bus_8[15:0]; // @[FDPEWrapper.scala 46:19]
  assign io_o_data_bus_9 = FDPE_io_o_data_bus_9[15:0]; // @[FDPEWrapper.scala 46:19]
  assign io_o_data_bus_10 = FDPE_io_o_data_bus_10[15:0]; // @[FDPEWrapper.scala 46:19]
  assign io_o_data_bus_11 = FDPE_io_o_data_bus_11[15:0]; // @[FDPEWrapper.scala 46:19]
  assign io_o_data_bus_12 = FDPE_io_o_data_bus_12[15:0]; // @[FDPEWrapper.scala 46:19]
  assign io_o_data_bus_13 = FDPE_io_o_data_bus_13[15:0]; // @[FDPEWrapper.scala 46:19]
  assign io_o_data_bus_14 = FDPE_io_o_data_bus_14[15:0]; // @[FDPEWrapper.scala 46:19]
  assign io_o_data_bus_15 = FDPE_io_o_data_bus_15[15:0]; // @[FDPEWrapper.scala 46:19]
  assign io_o_data_bus_16 = FDPE_io_o_data_bus_16[15:0]; // @[FDPEWrapper.scala 46:19]
  assign io_o_data_bus_17 = FDPE_io_o_data_bus_17[15:0]; // @[FDPEWrapper.scala 46:19]
  assign io_o_data_bus_18 = FDPE_io_o_data_bus_18[15:0]; // @[FDPEWrapper.scala 46:19]
  assign io_o_data_bus_19 = FDPE_io_o_data_bus_19[15:0]; // @[FDPEWrapper.scala 46:19]
  assign io_o_data_bus_20 = FDPE_io_o_data_bus_20[15:0]; // @[FDPEWrapper.scala 46:19]
  assign io_o_data_bus_21 = FDPE_io_o_data_bus_21[15:0]; // @[FDPEWrapper.scala 46:19]
  assign io_o_data_bus_22 = FDPE_io_o_data_bus_22[15:0]; // @[FDPEWrapper.scala 46:19]
  assign io_o_data_bus_23 = FDPE_io_o_data_bus_23[15:0]; // @[FDPEWrapper.scala 46:19]
  assign io_o_data_bus_24 = FDPE_io_o_data_bus_24[15:0]; // @[FDPEWrapper.scala 46:19]
  assign io_o_data_bus_25 = FDPE_io_o_data_bus_25[15:0]; // @[FDPEWrapper.scala 46:19]
  assign io_o_data_bus_26 = FDPE_io_o_data_bus_26[15:0]; // @[FDPEWrapper.scala 46:19]
  assign io_o_data_bus_27 = FDPE_io_o_data_bus_27[15:0]; // @[FDPEWrapper.scala 46:19]
  assign io_o_data_bus_28 = FDPE_io_o_data_bus_28[15:0]; // @[FDPEWrapper.scala 46:19]
  assign io_o_data_bus_29 = FDPE_io_o_data_bus_29[15:0]; // @[FDPEWrapper.scala 46:19]
  assign io_o_data_bus_30 = FDPE_io_o_data_bus_30[15:0]; // @[FDPEWrapper.scala 46:19]
  assign io_o_data_bus_31 = FDPE_io_o_data_bus_31[15:0]; // @[FDPEWrapper.scala 46:19]
  assign io_o_adder_0 = FDPE_io_o_adder_0[15:0]; // @[FDPEWrapper.scala 47:16]
  assign io_o_adder_1 = FDPE_io_o_adder_1[15:0]; // @[FDPEWrapper.scala 47:16]
  assign io_o_adder_2 = FDPE_io_o_adder_2[15:0]; // @[FDPEWrapper.scala 47:16]
  assign io_o_adder_3 = FDPE_io_o_adder_3[15:0]; // @[FDPEWrapper.scala 47:16]
  assign io_o_adder_4 = FDPE_io_o_adder_4[15:0]; // @[FDPEWrapper.scala 47:16]
  assign io_o_adder_5 = FDPE_io_o_adder_5[15:0]; // @[FDPEWrapper.scala 47:16]
  assign io_o_adder_6 = FDPE_io_o_adder_6[15:0]; // @[FDPEWrapper.scala 47:16]
  assign io_o_adder_7 = FDPE_io_o_adder_7[15:0]; // @[FDPEWrapper.scala 47:16]
  assign io_o_adder_8 = FDPE_io_o_adder_8[15:0]; // @[FDPEWrapper.scala 47:16]
  assign io_o_adder_9 = FDPE_io_o_adder_9[15:0]; // @[FDPEWrapper.scala 47:16]
  assign io_o_adder_10 = FDPE_io_o_adder_10[15:0]; // @[FDPEWrapper.scala 47:16]
  assign io_o_adder_11 = FDPE_io_o_adder_11[15:0]; // @[FDPEWrapper.scala 47:16]
  assign io_o_adder_12 = FDPE_io_o_adder_12[15:0]; // @[FDPEWrapper.scala 47:16]
  assign io_o_adder_13 = FDPE_io_o_adder_13[15:0]; // @[FDPEWrapper.scala 47:16]
  assign io_o_adder_14 = FDPE_io_o_adder_14[15:0]; // @[FDPEWrapper.scala 47:16]
  assign io_o_adder_15 = FDPE_io_o_adder_15[15:0]; // @[FDPEWrapper.scala 47:16]
  assign io_o_adder_16 = FDPE_io_o_adder_16[15:0]; // @[FDPEWrapper.scala 47:16]
  assign io_o_adder_17 = FDPE_io_o_adder_17[15:0]; // @[FDPEWrapper.scala 47:16]
  assign io_o_adder_18 = FDPE_io_o_adder_18[15:0]; // @[FDPEWrapper.scala 47:16]
  assign io_o_adder_19 = FDPE_io_o_adder_19[15:0]; // @[FDPEWrapper.scala 47:16]
  assign io_o_adder_20 = FDPE_io_o_adder_20[15:0]; // @[FDPEWrapper.scala 47:16]
  assign io_o_adder_21 = FDPE_io_o_adder_21[15:0]; // @[FDPEWrapper.scala 47:16]
  assign io_o_adder_22 = FDPE_io_o_adder_22[15:0]; // @[FDPEWrapper.scala 47:16]
  assign io_o_adder_23 = FDPE_io_o_adder_23[15:0]; // @[FDPEWrapper.scala 47:16]
  assign io_o_adder_24 = FDPE_io_o_adder_24[15:0]; // @[FDPEWrapper.scala 47:16]
  assign io_o_adder_25 = FDPE_io_o_adder_25[15:0]; // @[FDPEWrapper.scala 47:16]
  assign io_o_adder_26 = FDPE_io_o_adder_26[15:0]; // @[FDPEWrapper.scala 47:16]
  assign io_o_adder_27 = FDPE_io_o_adder_27[15:0]; // @[FDPEWrapper.scala 47:16]
  assign io_o_adder_28 = FDPE_io_o_adder_28[15:0]; // @[FDPEWrapper.scala 47:16]
  assign io_o_adder_29 = FDPE_io_o_adder_29[15:0]; // @[FDPEWrapper.scala 47:16]
  assign io_o_adder_30 = FDPE_io_o_adder_30[15:0]; // @[FDPEWrapper.scala 47:16]
  assign io_o_adder_31 = 16'h0; // @[FDPEWrapper.scala 47:16]
  assign FDPE_clock = clock;
  assign FDPE_reset = reset;
endmodule
