module stationary(
  input         clock,
  input         reset,
  input  [15:0] io_Stationary_matrix_0_0,
  input  [15:0] io_Stationary_matrix_0_1,
  input  [15:0] io_Stationary_matrix_0_2,
  input  [15:0] io_Stationary_matrix_0_3,
  input  [15:0] io_Stationary_matrix_0_4,
  input  [15:0] io_Stationary_matrix_0_5,
  input  [15:0] io_Stationary_matrix_0_6,
  input  [15:0] io_Stationary_matrix_0_7,
  input  [15:0] io_Stationary_matrix_1_0,
  input  [15:0] io_Stationary_matrix_1_1,
  input  [15:0] io_Stationary_matrix_1_2,
  input  [15:0] io_Stationary_matrix_1_3,
  input  [15:0] io_Stationary_matrix_1_4,
  input  [15:0] io_Stationary_matrix_1_5,
  input  [15:0] io_Stationary_matrix_1_6,
  input  [15:0] io_Stationary_matrix_1_7,
  input  [15:0] io_Stationary_matrix_2_0,
  input  [15:0] io_Stationary_matrix_2_1,
  input  [15:0] io_Stationary_matrix_2_2,
  input  [15:0] io_Stationary_matrix_2_3,
  input  [15:0] io_Stationary_matrix_2_4,
  input  [15:0] io_Stationary_matrix_2_5,
  input  [15:0] io_Stationary_matrix_2_6,
  input  [15:0] io_Stationary_matrix_2_7,
  input  [15:0] io_Stationary_matrix_3_0,
  input  [15:0] io_Stationary_matrix_3_1,
  input  [15:0] io_Stationary_matrix_3_2,
  input  [15:0] io_Stationary_matrix_3_3,
  input  [15:0] io_Stationary_matrix_3_4,
  input  [15:0] io_Stationary_matrix_3_5,
  input  [15:0] io_Stationary_matrix_3_6,
  input  [15:0] io_Stationary_matrix_3_7,
  input  [15:0] io_Stationary_matrix_4_0,
  input  [15:0] io_Stationary_matrix_4_1,
  input  [15:0] io_Stationary_matrix_4_2,
  input  [15:0] io_Stationary_matrix_4_3,
  input  [15:0] io_Stationary_matrix_4_4,
  input  [15:0] io_Stationary_matrix_4_5,
  input  [15:0] io_Stationary_matrix_4_6,
  input  [15:0] io_Stationary_matrix_4_7,
  input  [15:0] io_Stationary_matrix_5_0,
  input  [15:0] io_Stationary_matrix_5_1,
  input  [15:0] io_Stationary_matrix_5_2,
  input  [15:0] io_Stationary_matrix_5_3,
  input  [15:0] io_Stationary_matrix_5_4,
  input  [15:0] io_Stationary_matrix_5_5,
  input  [15:0] io_Stationary_matrix_5_6,
  input  [15:0] io_Stationary_matrix_5_7,
  input  [15:0] io_Stationary_matrix_6_0,
  input  [15:0] io_Stationary_matrix_6_1,
  input  [15:0] io_Stationary_matrix_6_2,
  input  [15:0] io_Stationary_matrix_6_3,
  input  [15:0] io_Stationary_matrix_6_4,
  input  [15:0] io_Stationary_matrix_6_5,
  input  [15:0] io_Stationary_matrix_6_6,
  input  [15:0] io_Stationary_matrix_6_7,
  input  [15:0] io_Stationary_matrix_7_0,
  input  [15:0] io_Stationary_matrix_7_1,
  input  [15:0] io_Stationary_matrix_7_2,
  input  [15:0] io_Stationary_matrix_7_3,
  input  [15:0] io_Stationary_matrix_7_4,
  input  [15:0] io_Stationary_matrix_7_5,
  input  [15:0] io_Stationary_matrix_7_6,
  input  [15:0] io_Stationary_matrix_7_7,
  output [15:0] io_o_Stationary_matrix1_0_0,
  output [15:0] io_o_Stationary_matrix1_0_1,
  output [15:0] io_o_Stationary_matrix1_0_2,
  output [15:0] io_o_Stationary_matrix1_0_3,
  output [15:0] io_o_Stationary_matrix1_0_4,
  output [15:0] io_o_Stationary_matrix1_0_5,
  output [15:0] io_o_Stationary_matrix1_0_6,
  output [15:0] io_o_Stationary_matrix1_0_7,
  output [15:0] io_o_Stationary_matrix1_1_0,
  output [15:0] io_o_Stationary_matrix1_1_1,
  output [15:0] io_o_Stationary_matrix1_1_2,
  output [15:0] io_o_Stationary_matrix1_1_3,
  output [15:0] io_o_Stationary_matrix1_1_4,
  output [15:0] io_o_Stationary_matrix1_1_5,
  output [15:0] io_o_Stationary_matrix1_1_6,
  output [15:0] io_o_Stationary_matrix1_1_7,
  output [15:0] io_o_Stationary_matrix1_2_0,
  output [15:0] io_o_Stationary_matrix1_2_1,
  output [15:0] io_o_Stationary_matrix1_2_2,
  output [15:0] io_o_Stationary_matrix1_2_3,
  output [15:0] io_o_Stationary_matrix1_2_4,
  output [15:0] io_o_Stationary_matrix1_2_5,
  output [15:0] io_o_Stationary_matrix1_2_6,
  output [15:0] io_o_Stationary_matrix1_2_7,
  output [15:0] io_o_Stationary_matrix1_3_0,
  output [15:0] io_o_Stationary_matrix1_3_1,
  output [15:0] io_o_Stationary_matrix1_3_2,
  output [15:0] io_o_Stationary_matrix1_3_3,
  output [15:0] io_o_Stationary_matrix1_3_4,
  output [15:0] io_o_Stationary_matrix1_3_5,
  output [15:0] io_o_Stationary_matrix1_3_6,
  output [15:0] io_o_Stationary_matrix1_3_7,
  output [15:0] io_o_Stationary_matrix1_4_0,
  output [15:0] io_o_Stationary_matrix1_4_1,
  output [15:0] io_o_Stationary_matrix1_4_2,
  output [15:0] io_o_Stationary_matrix1_4_3,
  output [15:0] io_o_Stationary_matrix1_4_4,
  output [15:0] io_o_Stationary_matrix1_4_5,
  output [15:0] io_o_Stationary_matrix1_4_6,
  output [15:0] io_o_Stationary_matrix1_4_7,
  output [15:0] io_o_Stationary_matrix1_5_0,
  output [15:0] io_o_Stationary_matrix1_5_1,
  output [15:0] io_o_Stationary_matrix1_5_2,
  output [15:0] io_o_Stationary_matrix1_5_3,
  output [15:0] io_o_Stationary_matrix1_5_4,
  output [15:0] io_o_Stationary_matrix1_5_5,
  output [15:0] io_o_Stationary_matrix1_5_6,
  output [15:0] io_o_Stationary_matrix1_5_7,
  output [15:0] io_o_Stationary_matrix1_6_0,
  output [15:0] io_o_Stationary_matrix1_6_1,
  output [15:0] io_o_Stationary_matrix1_6_2,
  output [15:0] io_o_Stationary_matrix1_6_3,
  output [15:0] io_o_Stationary_matrix1_6_4,
  output [15:0] io_o_Stationary_matrix1_6_5,
  output [15:0] io_o_Stationary_matrix1_6_6,
  output [15:0] io_o_Stationary_matrix1_6_7,
  output [15:0] io_o_Stationary_matrix1_7_0,
  output [15:0] io_o_Stationary_matrix1_7_1,
  output [15:0] io_o_Stationary_matrix1_7_2,
  output [15:0] io_o_Stationary_matrix1_7_3,
  output [15:0] io_o_Stationary_matrix1_7_4,
  output [15:0] io_o_Stationary_matrix1_7_5,
  output [15:0] io_o_Stationary_matrix1_7_6,
  output [15:0] io_o_Stationary_matrix1_7_7,
  output [15:0] io_o_Stationary_matrix2_0_0,
  output [15:0] io_o_Stationary_matrix2_0_1,
  output [15:0] io_o_Stationary_matrix2_0_2,
  output [15:0] io_o_Stationary_matrix2_0_3,
  output [15:0] io_o_Stationary_matrix2_0_4,
  output [15:0] io_o_Stationary_matrix2_0_5,
  output [15:0] io_o_Stationary_matrix2_0_6,
  output [15:0] io_o_Stationary_matrix2_0_7,
  output [15:0] io_o_Stationary_matrix2_1_0,
  output [15:0] io_o_Stationary_matrix2_1_1,
  output [15:0] io_o_Stationary_matrix2_1_2,
  output [15:0] io_o_Stationary_matrix2_1_3,
  output [15:0] io_o_Stationary_matrix2_1_4,
  output [15:0] io_o_Stationary_matrix2_1_5,
  output [15:0] io_o_Stationary_matrix2_1_6,
  output [15:0] io_o_Stationary_matrix2_1_7,
  output [15:0] io_o_Stationary_matrix2_2_0,
  output [15:0] io_o_Stationary_matrix2_2_1,
  output [15:0] io_o_Stationary_matrix2_2_2,
  output [15:0] io_o_Stationary_matrix2_2_3,
  output [15:0] io_o_Stationary_matrix2_2_4,
  output [15:0] io_o_Stationary_matrix2_2_5,
  output [15:0] io_o_Stationary_matrix2_2_6,
  output [15:0] io_o_Stationary_matrix2_2_7,
  output [15:0] io_o_Stationary_matrix2_3_0,
  output [15:0] io_o_Stationary_matrix2_3_1,
  output [15:0] io_o_Stationary_matrix2_3_2,
  output [15:0] io_o_Stationary_matrix2_3_3,
  output [15:0] io_o_Stationary_matrix2_3_4,
  output [15:0] io_o_Stationary_matrix2_3_5,
  output [15:0] io_o_Stationary_matrix2_3_6,
  output [15:0] io_o_Stationary_matrix2_3_7,
  output [15:0] io_o_Stationary_matrix2_4_0,
  output [15:0] io_o_Stationary_matrix2_4_1,
  output [15:0] io_o_Stationary_matrix2_4_2,
  output [15:0] io_o_Stationary_matrix2_4_3,
  output [15:0] io_o_Stationary_matrix2_4_4,
  output [15:0] io_o_Stationary_matrix2_4_5,
  output [15:0] io_o_Stationary_matrix2_4_6,
  output [15:0] io_o_Stationary_matrix2_4_7,
  output [15:0] io_o_Stationary_matrix2_5_0,
  output [15:0] io_o_Stationary_matrix2_5_1,
  output [15:0] io_o_Stationary_matrix2_5_2,
  output [15:0] io_o_Stationary_matrix2_5_3,
  output [15:0] io_o_Stationary_matrix2_5_4,
  output [15:0] io_o_Stationary_matrix2_5_5,
  output [15:0] io_o_Stationary_matrix2_5_6,
  output [15:0] io_o_Stationary_matrix2_5_7,
  output [15:0] io_o_Stationary_matrix2_6_0,
  output [15:0] io_o_Stationary_matrix2_6_1,
  output [15:0] io_o_Stationary_matrix2_6_2,
  output [15:0] io_o_Stationary_matrix2_6_3,
  output [15:0] io_o_Stationary_matrix2_6_4,
  output [15:0] io_o_Stationary_matrix2_6_5,
  output [15:0] io_o_Stationary_matrix2_6_6,
  output [15:0] io_o_Stationary_matrix2_6_7,
  output [15:0] io_o_Stationary_matrix2_7_0,
  output [15:0] io_o_Stationary_matrix2_7_1,
  output [15:0] io_o_Stationary_matrix2_7_2,
  output [15:0] io_o_Stationary_matrix2_7_3,
  output [15:0] io_o_Stationary_matrix2_7_4,
  output [15:0] io_o_Stationary_matrix2_7_5,
  output [15:0] io_o_Stationary_matrix2_7_6,
  output [15:0] io_o_Stationary_matrix2_7_7,
  output [15:0] io_o_Stationary_matrix3_0_0,
  output [15:0] io_o_Stationary_matrix3_0_1,
  output [15:0] io_o_Stationary_matrix3_0_2,
  output [15:0] io_o_Stationary_matrix3_0_3,
  output [15:0] io_o_Stationary_matrix3_0_4,
  output [15:0] io_o_Stationary_matrix3_0_5,
  output [15:0] io_o_Stationary_matrix3_0_6,
  output [15:0] io_o_Stationary_matrix3_0_7,
  output [15:0] io_o_Stationary_matrix3_1_0,
  output [15:0] io_o_Stationary_matrix3_1_1,
  output [15:0] io_o_Stationary_matrix3_1_2,
  output [15:0] io_o_Stationary_matrix3_1_3,
  output [15:0] io_o_Stationary_matrix3_1_4,
  output [15:0] io_o_Stationary_matrix3_1_5,
  output [15:0] io_o_Stationary_matrix3_1_6,
  output [15:0] io_o_Stationary_matrix3_1_7,
  output [15:0] io_o_Stationary_matrix3_2_0,
  output [15:0] io_o_Stationary_matrix3_2_1,
  output [15:0] io_o_Stationary_matrix3_2_2,
  output [15:0] io_o_Stationary_matrix3_2_3,
  output [15:0] io_o_Stationary_matrix3_2_4,
  output [15:0] io_o_Stationary_matrix3_2_5,
  output [15:0] io_o_Stationary_matrix3_2_6,
  output [15:0] io_o_Stationary_matrix3_2_7,
  output [15:0] io_o_Stationary_matrix3_3_0,
  output [15:0] io_o_Stationary_matrix3_3_1,
  output [15:0] io_o_Stationary_matrix3_3_2,
  output [15:0] io_o_Stationary_matrix3_3_3,
  output [15:0] io_o_Stationary_matrix3_3_4,
  output [15:0] io_o_Stationary_matrix3_3_5,
  output [15:0] io_o_Stationary_matrix3_3_6,
  output [15:0] io_o_Stationary_matrix3_3_7,
  output [15:0] io_o_Stationary_matrix3_4_0,
  output [15:0] io_o_Stationary_matrix3_4_1,
  output [15:0] io_o_Stationary_matrix3_4_2,
  output [15:0] io_o_Stationary_matrix3_4_3,
  output [15:0] io_o_Stationary_matrix3_4_4,
  output [15:0] io_o_Stationary_matrix3_4_5,
  output [15:0] io_o_Stationary_matrix3_4_6,
  output [15:0] io_o_Stationary_matrix3_4_7,
  output [15:0] io_o_Stationary_matrix3_5_0,
  output [15:0] io_o_Stationary_matrix3_5_1,
  output [15:0] io_o_Stationary_matrix3_5_2,
  output [15:0] io_o_Stationary_matrix3_5_3,
  output [15:0] io_o_Stationary_matrix3_5_4,
  output [15:0] io_o_Stationary_matrix3_5_5,
  output [15:0] io_o_Stationary_matrix3_5_6,
  output [15:0] io_o_Stationary_matrix3_5_7,
  output [15:0] io_o_Stationary_matrix3_6_0,
  output [15:0] io_o_Stationary_matrix3_6_1,
  output [15:0] io_o_Stationary_matrix3_6_2,
  output [15:0] io_o_Stationary_matrix3_6_3,
  output [15:0] io_o_Stationary_matrix3_6_4,
  output [15:0] io_o_Stationary_matrix3_6_5,
  output [15:0] io_o_Stationary_matrix3_6_6,
  output [15:0] io_o_Stationary_matrix3_6_7,
  output [15:0] io_o_Stationary_matrix3_7_0,
  output [15:0] io_o_Stationary_matrix3_7_1,
  output [15:0] io_o_Stationary_matrix3_7_2,
  output [15:0] io_o_Stationary_matrix3_7_3,
  output [15:0] io_o_Stationary_matrix3_7_4,
  output [15:0] io_o_Stationary_matrix3_7_5,
  output [15:0] io_o_Stationary_matrix3_7_6,
  output [15:0] io_o_Stationary_matrix3_7_7,
  output [15:0] io_o_Stationary_matrix4_0_0,
  output [15:0] io_o_Stationary_matrix4_0_1,
  output [15:0] io_o_Stationary_matrix4_0_2,
  output [15:0] io_o_Stationary_matrix4_0_3,
  output [15:0] io_o_Stationary_matrix4_0_4,
  output [15:0] io_o_Stationary_matrix4_0_5,
  output [15:0] io_o_Stationary_matrix4_0_6,
  output [15:0] io_o_Stationary_matrix4_0_7,
  output [15:0] io_o_Stationary_matrix4_1_0,
  output [15:0] io_o_Stationary_matrix4_1_1,
  output [15:0] io_o_Stationary_matrix4_1_2,
  output [15:0] io_o_Stationary_matrix4_1_3,
  output [15:0] io_o_Stationary_matrix4_1_4,
  output [15:0] io_o_Stationary_matrix4_1_5,
  output [15:0] io_o_Stationary_matrix4_1_6,
  output [15:0] io_o_Stationary_matrix4_1_7,
  output [15:0] io_o_Stationary_matrix4_2_0,
  output [15:0] io_o_Stationary_matrix4_2_1,
  output [15:0] io_o_Stationary_matrix4_2_2,
  output [15:0] io_o_Stationary_matrix4_2_3,
  output [15:0] io_o_Stationary_matrix4_2_4,
  output [15:0] io_o_Stationary_matrix4_2_5,
  output [15:0] io_o_Stationary_matrix4_2_6,
  output [15:0] io_o_Stationary_matrix4_2_7,
  output [15:0] io_o_Stationary_matrix4_3_0,
  output [15:0] io_o_Stationary_matrix4_3_1,
  output [15:0] io_o_Stationary_matrix4_3_2,
  output [15:0] io_o_Stationary_matrix4_3_3,
  output [15:0] io_o_Stationary_matrix4_3_4,
  output [15:0] io_o_Stationary_matrix4_3_5,
  output [15:0] io_o_Stationary_matrix4_3_6,
  output [15:0] io_o_Stationary_matrix4_3_7,
  output [15:0] io_o_Stationary_matrix4_4_0,
  output [15:0] io_o_Stationary_matrix4_4_1,
  output [15:0] io_o_Stationary_matrix4_4_2,
  output [15:0] io_o_Stationary_matrix4_4_3,
  output [15:0] io_o_Stationary_matrix4_4_4,
  output [15:0] io_o_Stationary_matrix4_4_5,
  output [15:0] io_o_Stationary_matrix4_4_6,
  output [15:0] io_o_Stationary_matrix4_4_7,
  output [15:0] io_o_Stationary_matrix4_5_0,
  output [15:0] io_o_Stationary_matrix4_5_1,
  output [15:0] io_o_Stationary_matrix4_5_2,
  output [15:0] io_o_Stationary_matrix4_5_3,
  output [15:0] io_o_Stationary_matrix4_5_4,
  output [15:0] io_o_Stationary_matrix4_5_5,
  output [15:0] io_o_Stationary_matrix4_5_6,
  output [15:0] io_o_Stationary_matrix4_5_7,
  output [15:0] io_o_Stationary_matrix4_6_0,
  output [15:0] io_o_Stationary_matrix4_6_1,
  output [15:0] io_o_Stationary_matrix4_6_2,
  output [15:0] io_o_Stationary_matrix4_6_3,
  output [15:0] io_o_Stationary_matrix4_6_4,
  output [15:0] io_o_Stationary_matrix4_6_5,
  output [15:0] io_o_Stationary_matrix4_6_6,
  output [15:0] io_o_Stationary_matrix4_6_7,
  output [15:0] io_o_Stationary_matrix4_7_0,
  output [15:0] io_o_Stationary_matrix4_7_1,
  output [15:0] io_o_Stationary_matrix4_7_2,
  output [15:0] io_o_Stationary_matrix4_7_3,
  output [15:0] io_o_Stationary_matrix4_7_4,
  output [15:0] io_o_Stationary_matrix4_7_5,
  output [15:0] io_o_Stationary_matrix4_7_6,
  output [15:0] io_o_Stationary_matrix4_7_7,
  output [15:0] io_o_Stationary_matrix5_0_0,
  output [15:0] io_o_Stationary_matrix5_0_1,
  output [15:0] io_o_Stationary_matrix5_0_2,
  output [15:0] io_o_Stationary_matrix5_0_3,
  output [15:0] io_o_Stationary_matrix5_0_4,
  output [15:0] io_o_Stationary_matrix5_0_5,
  output [15:0] io_o_Stationary_matrix5_0_6,
  output [15:0] io_o_Stationary_matrix5_0_7,
  output [15:0] io_o_Stationary_matrix5_1_0,
  output [15:0] io_o_Stationary_matrix5_1_1,
  output [15:0] io_o_Stationary_matrix5_1_2,
  output [15:0] io_o_Stationary_matrix5_1_3,
  output [15:0] io_o_Stationary_matrix5_1_4,
  output [15:0] io_o_Stationary_matrix5_1_5,
  output [15:0] io_o_Stationary_matrix5_1_6,
  output [15:0] io_o_Stationary_matrix5_1_7,
  output [15:0] io_o_Stationary_matrix5_2_0,
  output [15:0] io_o_Stationary_matrix5_2_1,
  output [15:0] io_o_Stationary_matrix5_2_2,
  output [15:0] io_o_Stationary_matrix5_2_3,
  output [15:0] io_o_Stationary_matrix5_2_4,
  output [15:0] io_o_Stationary_matrix5_2_5,
  output [15:0] io_o_Stationary_matrix5_2_6,
  output [15:0] io_o_Stationary_matrix5_2_7,
  output [15:0] io_o_Stationary_matrix5_3_0,
  output [15:0] io_o_Stationary_matrix5_3_1,
  output [15:0] io_o_Stationary_matrix5_3_2,
  output [15:0] io_o_Stationary_matrix5_3_3,
  output [15:0] io_o_Stationary_matrix5_3_4,
  output [15:0] io_o_Stationary_matrix5_3_5,
  output [15:0] io_o_Stationary_matrix5_3_6,
  output [15:0] io_o_Stationary_matrix5_3_7,
  output [15:0] io_o_Stationary_matrix5_4_0,
  output [15:0] io_o_Stationary_matrix5_4_1,
  output [15:0] io_o_Stationary_matrix5_4_2,
  output [15:0] io_o_Stationary_matrix5_4_3,
  output [15:0] io_o_Stationary_matrix5_4_4,
  output [15:0] io_o_Stationary_matrix5_4_5,
  output [15:0] io_o_Stationary_matrix5_4_6,
  output [15:0] io_o_Stationary_matrix5_4_7,
  output [15:0] io_o_Stationary_matrix5_5_0,
  output [15:0] io_o_Stationary_matrix5_5_1,
  output [15:0] io_o_Stationary_matrix5_5_2,
  output [15:0] io_o_Stationary_matrix5_5_3,
  output [15:0] io_o_Stationary_matrix5_5_4,
  output [15:0] io_o_Stationary_matrix5_5_5,
  output [15:0] io_o_Stationary_matrix5_5_6,
  output [15:0] io_o_Stationary_matrix5_5_7,
  output [15:0] io_o_Stationary_matrix5_6_0,
  output [15:0] io_o_Stationary_matrix5_6_1,
  output [15:0] io_o_Stationary_matrix5_6_2,
  output [15:0] io_o_Stationary_matrix5_6_3,
  output [15:0] io_o_Stationary_matrix5_6_4,
  output [15:0] io_o_Stationary_matrix5_6_5,
  output [15:0] io_o_Stationary_matrix5_6_6,
  output [15:0] io_o_Stationary_matrix5_6_7,
  output [15:0] io_o_Stationary_matrix5_7_0,
  output [15:0] io_o_Stationary_matrix5_7_1,
  output [15:0] io_o_Stationary_matrix5_7_2,
  output [15:0] io_o_Stationary_matrix5_7_3,
  output [15:0] io_o_Stationary_matrix5_7_4,
  output [15:0] io_o_Stationary_matrix5_7_5,
  output [15:0] io_o_Stationary_matrix5_7_6,
  output [15:0] io_o_Stationary_matrix5_7_7,
  output [15:0] io_o_Stationary_matrix6_0_0,
  output [15:0] io_o_Stationary_matrix6_0_1,
  output [15:0] io_o_Stationary_matrix6_0_2,
  output [15:0] io_o_Stationary_matrix6_0_3,
  output [15:0] io_o_Stationary_matrix6_0_4,
  output [15:0] io_o_Stationary_matrix6_0_5,
  output [15:0] io_o_Stationary_matrix6_0_6,
  output [15:0] io_o_Stationary_matrix6_0_7,
  output [15:0] io_o_Stationary_matrix6_1_0,
  output [15:0] io_o_Stationary_matrix6_1_1,
  output [15:0] io_o_Stationary_matrix6_1_2,
  output [15:0] io_o_Stationary_matrix6_1_3,
  output [15:0] io_o_Stationary_matrix6_1_4,
  output [15:0] io_o_Stationary_matrix6_1_5,
  output [15:0] io_o_Stationary_matrix6_1_6,
  output [15:0] io_o_Stationary_matrix6_1_7,
  output [15:0] io_o_Stationary_matrix6_2_0,
  output [15:0] io_o_Stationary_matrix6_2_1,
  output [15:0] io_o_Stationary_matrix6_2_2,
  output [15:0] io_o_Stationary_matrix6_2_3,
  output [15:0] io_o_Stationary_matrix6_2_4,
  output [15:0] io_o_Stationary_matrix6_2_5,
  output [15:0] io_o_Stationary_matrix6_2_6,
  output [15:0] io_o_Stationary_matrix6_2_7,
  output [15:0] io_o_Stationary_matrix6_3_0,
  output [15:0] io_o_Stationary_matrix6_3_1,
  output [15:0] io_o_Stationary_matrix6_3_2,
  output [15:0] io_o_Stationary_matrix6_3_3,
  output [15:0] io_o_Stationary_matrix6_3_4,
  output [15:0] io_o_Stationary_matrix6_3_5,
  output [15:0] io_o_Stationary_matrix6_3_6,
  output [15:0] io_o_Stationary_matrix6_3_7,
  output [15:0] io_o_Stationary_matrix6_4_0,
  output [15:0] io_o_Stationary_matrix6_4_1,
  output [15:0] io_o_Stationary_matrix6_4_2,
  output [15:0] io_o_Stationary_matrix6_4_3,
  output [15:0] io_o_Stationary_matrix6_4_4,
  output [15:0] io_o_Stationary_matrix6_4_5,
  output [15:0] io_o_Stationary_matrix6_4_6,
  output [15:0] io_o_Stationary_matrix6_4_7,
  output [15:0] io_o_Stationary_matrix6_5_0,
  output [15:0] io_o_Stationary_matrix6_5_1,
  output [15:0] io_o_Stationary_matrix6_5_2,
  output [15:0] io_o_Stationary_matrix6_5_3,
  output [15:0] io_o_Stationary_matrix6_5_4,
  output [15:0] io_o_Stationary_matrix6_5_5,
  output [15:0] io_o_Stationary_matrix6_5_6,
  output [15:0] io_o_Stationary_matrix6_5_7,
  output [15:0] io_o_Stationary_matrix6_6_0,
  output [15:0] io_o_Stationary_matrix6_6_1,
  output [15:0] io_o_Stationary_matrix6_6_2,
  output [15:0] io_o_Stationary_matrix6_6_3,
  output [15:0] io_o_Stationary_matrix6_6_4,
  output [15:0] io_o_Stationary_matrix6_6_5,
  output [15:0] io_o_Stationary_matrix6_6_6,
  output [15:0] io_o_Stationary_matrix6_6_7,
  output [15:0] io_o_Stationary_matrix6_7_0,
  output [15:0] io_o_Stationary_matrix6_7_1,
  output [15:0] io_o_Stationary_matrix6_7_2,
  output [15:0] io_o_Stationary_matrix6_7_3,
  output [15:0] io_o_Stationary_matrix6_7_4,
  output [15:0] io_o_Stationary_matrix6_7_5,
  output [15:0] io_o_Stationary_matrix6_7_6,
  output [15:0] io_o_Stationary_matrix6_7_7,
  output [15:0] io_o_Stationary_matrix7_0_0,
  output [15:0] io_o_Stationary_matrix7_0_1,
  output [15:0] io_o_Stationary_matrix7_0_2,
  output [15:0] io_o_Stationary_matrix7_0_3,
  output [15:0] io_o_Stationary_matrix7_0_4,
  output [15:0] io_o_Stationary_matrix7_0_5,
  output [15:0] io_o_Stationary_matrix7_0_6,
  output [15:0] io_o_Stationary_matrix7_0_7,
  output [15:0] io_o_Stationary_matrix7_1_0,
  output [15:0] io_o_Stationary_matrix7_1_1,
  output [15:0] io_o_Stationary_matrix7_1_2,
  output [15:0] io_o_Stationary_matrix7_1_3,
  output [15:0] io_o_Stationary_matrix7_1_4,
  output [15:0] io_o_Stationary_matrix7_1_5,
  output [15:0] io_o_Stationary_matrix7_1_6,
  output [15:0] io_o_Stationary_matrix7_1_7,
  output [15:0] io_o_Stationary_matrix7_2_0,
  output [15:0] io_o_Stationary_matrix7_2_1,
  output [15:0] io_o_Stationary_matrix7_2_2,
  output [15:0] io_o_Stationary_matrix7_2_3,
  output [15:0] io_o_Stationary_matrix7_2_4,
  output [15:0] io_o_Stationary_matrix7_2_5,
  output [15:0] io_o_Stationary_matrix7_2_6,
  output [15:0] io_o_Stationary_matrix7_2_7,
  output [15:0] io_o_Stationary_matrix7_3_0,
  output [15:0] io_o_Stationary_matrix7_3_1,
  output [15:0] io_o_Stationary_matrix7_3_2,
  output [15:0] io_o_Stationary_matrix7_3_3,
  output [15:0] io_o_Stationary_matrix7_3_4,
  output [15:0] io_o_Stationary_matrix7_3_5,
  output [15:0] io_o_Stationary_matrix7_3_6,
  output [15:0] io_o_Stationary_matrix7_3_7,
  output [15:0] io_o_Stationary_matrix7_4_0,
  output [15:0] io_o_Stationary_matrix7_4_1,
  output [15:0] io_o_Stationary_matrix7_4_2,
  output [15:0] io_o_Stationary_matrix7_4_3,
  output [15:0] io_o_Stationary_matrix7_4_4,
  output [15:0] io_o_Stationary_matrix7_4_5,
  output [15:0] io_o_Stationary_matrix7_4_6,
  output [15:0] io_o_Stationary_matrix7_4_7,
  output [15:0] io_o_Stationary_matrix7_5_0,
  output [15:0] io_o_Stationary_matrix7_5_1,
  output [15:0] io_o_Stationary_matrix7_5_2,
  output [15:0] io_o_Stationary_matrix7_5_3,
  output [15:0] io_o_Stationary_matrix7_5_4,
  output [15:0] io_o_Stationary_matrix7_5_5,
  output [15:0] io_o_Stationary_matrix7_5_6,
  output [15:0] io_o_Stationary_matrix7_5_7,
  output [15:0] io_o_Stationary_matrix7_6_0,
  output [15:0] io_o_Stationary_matrix7_6_1,
  output [15:0] io_o_Stationary_matrix7_6_2,
  output [15:0] io_o_Stationary_matrix7_6_3,
  output [15:0] io_o_Stationary_matrix7_6_4,
  output [15:0] io_o_Stationary_matrix7_6_5,
  output [15:0] io_o_Stationary_matrix7_6_6,
  output [15:0] io_o_Stationary_matrix7_6_7,
  output [15:0] io_o_Stationary_matrix7_7_0,
  output [15:0] io_o_Stationary_matrix7_7_1,
  output [15:0] io_o_Stationary_matrix7_7_2,
  output [15:0] io_o_Stationary_matrix7_7_3,
  output [15:0] io_o_Stationary_matrix7_7_4,
  output [15:0] io_o_Stationary_matrix7_7_5,
  output [15:0] io_o_Stationary_matrix7_7_6,
  output [15:0] io_o_Stationary_matrix7_7_7,
  output [15:0] io_o_Stationary_matrix8_0_0,
  output [15:0] io_o_Stationary_matrix8_0_1,
  output [15:0] io_o_Stationary_matrix8_0_2,
  output [15:0] io_o_Stationary_matrix8_0_3,
  output [15:0] io_o_Stationary_matrix8_0_4,
  output [15:0] io_o_Stationary_matrix8_0_5,
  output [15:0] io_o_Stationary_matrix8_0_6,
  output [15:0] io_o_Stationary_matrix8_0_7,
  output [15:0] io_o_Stationary_matrix8_1_0,
  output [15:0] io_o_Stationary_matrix8_1_1,
  output [15:0] io_o_Stationary_matrix8_1_2,
  output [15:0] io_o_Stationary_matrix8_1_3,
  output [15:0] io_o_Stationary_matrix8_1_4,
  output [15:0] io_o_Stationary_matrix8_1_5,
  output [15:0] io_o_Stationary_matrix8_1_6,
  output [15:0] io_o_Stationary_matrix8_1_7,
  output [15:0] io_o_Stationary_matrix8_2_0,
  output [15:0] io_o_Stationary_matrix8_2_1,
  output [15:0] io_o_Stationary_matrix8_2_2,
  output [15:0] io_o_Stationary_matrix8_2_3,
  output [15:0] io_o_Stationary_matrix8_2_4,
  output [15:0] io_o_Stationary_matrix8_2_5,
  output [15:0] io_o_Stationary_matrix8_2_6,
  output [15:0] io_o_Stationary_matrix8_2_7,
  output [15:0] io_o_Stationary_matrix8_3_0,
  output [15:0] io_o_Stationary_matrix8_3_1,
  output [15:0] io_o_Stationary_matrix8_3_2,
  output [15:0] io_o_Stationary_matrix8_3_3,
  output [15:0] io_o_Stationary_matrix8_3_4,
  output [15:0] io_o_Stationary_matrix8_3_5,
  output [15:0] io_o_Stationary_matrix8_3_6,
  output [15:0] io_o_Stationary_matrix8_3_7,
  output [15:0] io_o_Stationary_matrix8_4_0,
  output [15:0] io_o_Stationary_matrix8_4_1,
  output [15:0] io_o_Stationary_matrix8_4_2,
  output [15:0] io_o_Stationary_matrix8_4_3,
  output [15:0] io_o_Stationary_matrix8_4_4,
  output [15:0] io_o_Stationary_matrix8_4_5,
  output [15:0] io_o_Stationary_matrix8_4_6,
  output [15:0] io_o_Stationary_matrix8_4_7,
  output [15:0] io_o_Stationary_matrix8_5_0,
  output [15:0] io_o_Stationary_matrix8_5_1,
  output [15:0] io_o_Stationary_matrix8_5_2,
  output [15:0] io_o_Stationary_matrix8_5_3,
  output [15:0] io_o_Stationary_matrix8_5_4,
  output [15:0] io_o_Stationary_matrix8_5_5,
  output [15:0] io_o_Stationary_matrix8_5_6,
  output [15:0] io_o_Stationary_matrix8_5_7,
  output [15:0] io_o_Stationary_matrix8_6_0,
  output [15:0] io_o_Stationary_matrix8_6_1,
  output [15:0] io_o_Stationary_matrix8_6_2,
  output [15:0] io_o_Stationary_matrix8_6_3,
  output [15:0] io_o_Stationary_matrix8_6_4,
  output [15:0] io_o_Stationary_matrix8_6_5,
  output [15:0] io_o_Stationary_matrix8_6_6,
  output [15:0] io_o_Stationary_matrix8_6_7,
  output [15:0] io_o_Stationary_matrix8_7_0,
  output [15:0] io_o_Stationary_matrix8_7_1,
  output [15:0] io_o_Stationary_matrix8_7_2,
  output [15:0] io_o_Stationary_matrix8_7_3,
  output [15:0] io_o_Stationary_matrix8_7_4,
  output [15:0] io_o_Stationary_matrix8_7_5,
  output [15:0] io_o_Stationary_matrix8_7_6,
  output [15:0] io_o_Stationary_matrix8_7_7
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] count; // @[stationary_dpe.scala 23:27]
  reg [15:0] Station2_0_0; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_0_1; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_0_2; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_0_3; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_0_4; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_0_5; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_0_6; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_0_7; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_1_0; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_1_1; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_1_2; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_1_3; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_1_4; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_1_5; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_1_6; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_1_7; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_2_0; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_2_1; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_2_2; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_2_3; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_2_4; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_2_5; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_2_6; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_2_7; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_3_0; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_3_1; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_3_2; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_3_3; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_3_4; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_3_5; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_3_6; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_3_7; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_4_0; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_4_1; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_4_2; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_4_3; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_4_4; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_4_5; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_4_6; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_4_7; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_5_0; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_5_1; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_5_2; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_5_3; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_5_4; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_5_5; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_5_6; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_5_7; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_6_0; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_6_1; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_6_2; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_6_3; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_6_4; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_6_5; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_6_6; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_6_7; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_7_0; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_7_1; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_7_2; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_7_3; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_7_4; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_7_5; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_7_6; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_7_7; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station3_0_0; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_0_1; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_0_2; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_0_3; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_0_4; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_0_5; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_0_6; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_0_7; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_1_0; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_1_1; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_1_2; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_1_3; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_1_4; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_1_5; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_1_6; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_1_7; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_2_0; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_2_1; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_2_2; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_2_3; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_2_4; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_2_5; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_2_6; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_2_7; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_3_0; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_3_1; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_3_2; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_3_3; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_3_4; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_3_5; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_3_6; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_3_7; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_4_0; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_4_1; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_4_2; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_4_3; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_4_4; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_4_5; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_4_6; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_4_7; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_5_0; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_5_1; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_5_2; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_5_3; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_5_4; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_5_5; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_5_6; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_5_7; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_6_0; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_6_1; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_6_2; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_6_3; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_6_4; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_6_5; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_6_6; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_6_7; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_7_0; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_7_1; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_7_2; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_7_3; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_7_4; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_7_5; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_7_6; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_7_7; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station4_0_0; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_0_1; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_0_2; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_0_3; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_0_4; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_0_5; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_0_6; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_0_7; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_1_0; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_1_1; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_1_2; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_1_3; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_1_4; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_1_5; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_1_6; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_1_7; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_2_0; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_2_1; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_2_2; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_2_3; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_2_4; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_2_5; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_2_6; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_2_7; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_3_0; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_3_1; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_3_2; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_3_3; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_3_4; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_3_5; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_3_6; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_3_7; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_4_0; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_4_1; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_4_2; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_4_3; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_4_4; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_4_5; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_4_6; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_4_7; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_5_0; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_5_1; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_5_2; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_5_3; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_5_4; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_5_5; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_5_6; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_5_7; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_6_0; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_6_1; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_6_2; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_6_3; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_6_4; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_6_5; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_6_6; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_6_7; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_7_0; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_7_1; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_7_2; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_7_3; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_7_4; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_7_5; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_7_6; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_7_7; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station5_0_0; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_0_1; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_0_2; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_0_3; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_0_4; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_0_5; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_0_6; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_0_7; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_1_0; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_1_1; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_1_2; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_1_3; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_1_4; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_1_5; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_1_6; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_1_7; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_2_0; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_2_1; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_2_2; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_2_3; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_2_4; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_2_5; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_2_6; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_2_7; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_3_0; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_3_1; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_3_2; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_3_3; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_3_4; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_3_5; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_3_6; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_3_7; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_4_0; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_4_1; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_4_2; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_4_3; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_4_4; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_4_5; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_4_6; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_4_7; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_5_0; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_5_1; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_5_2; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_5_3; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_5_4; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_5_5; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_5_6; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_5_7; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_6_0; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_6_1; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_6_2; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_6_3; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_6_4; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_6_5; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_6_6; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_6_7; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_7_0; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_7_1; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_7_2; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_7_3; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_7_4; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_7_5; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_7_6; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_7_7; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station6_0_0; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_0_1; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_0_2; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_0_3; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_0_4; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_0_5; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_0_6; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_0_7; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_1_0; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_1_1; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_1_2; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_1_3; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_1_4; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_1_5; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_1_6; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_1_7; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_2_0; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_2_1; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_2_2; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_2_3; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_2_4; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_2_5; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_2_6; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_2_7; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_3_0; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_3_1; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_3_2; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_3_3; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_3_4; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_3_5; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_3_6; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_3_7; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_4_0; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_4_1; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_4_2; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_4_3; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_4_4; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_4_5; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_4_6; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_4_7; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_5_0; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_5_1; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_5_2; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_5_3; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_5_4; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_5_5; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_5_6; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_5_7; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_6_0; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_6_1; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_6_2; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_6_3; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_6_4; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_6_5; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_6_6; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_6_7; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_7_0; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_7_1; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_7_2; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_7_3; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_7_4; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_7_5; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_7_6; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_7_7; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station7_0_0; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_0_1; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_0_2; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_0_3; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_0_4; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_0_5; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_0_6; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_0_7; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_1_0; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_1_1; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_1_2; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_1_3; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_1_4; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_1_5; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_1_6; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_1_7; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_2_0; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_2_1; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_2_2; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_2_3; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_2_4; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_2_5; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_2_6; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_2_7; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_3_0; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_3_1; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_3_2; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_3_3; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_3_4; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_3_5; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_3_6; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_3_7; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_4_0; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_4_1; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_4_2; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_4_3; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_4_4; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_4_5; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_4_6; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_4_7; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_5_0; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_5_1; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_5_2; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_5_3; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_5_4; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_5_5; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_5_6; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_5_7; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_6_0; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_6_1; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_6_2; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_6_3; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_6_4; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_6_5; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_6_6; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_6_7; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_7_0; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_7_1; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_7_2; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_7_3; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_7_4; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_7_5; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_7_6; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_7_7; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station8_0_0; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_0_1; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_0_2; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_0_3; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_0_4; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_0_5; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_0_6; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_0_7; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_1_0; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_1_1; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_1_2; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_1_3; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_1_4; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_1_5; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_1_6; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_1_7; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_2_0; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_2_1; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_2_2; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_2_3; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_2_4; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_2_5; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_2_6; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_2_7; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_3_0; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_3_1; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_3_2; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_3_3; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_3_4; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_3_5; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_3_6; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_3_7; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_4_0; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_4_1; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_4_2; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_4_3; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_4_4; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_4_5; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_4_6; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_4_7; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_5_0; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_5_1; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_5_2; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_5_3; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_5_4; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_5_5; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_5_6; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_5_7; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_6_0; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_6_1; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_6_2; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_6_3; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_6_4; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_6_5; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_6_6; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_6_7; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_7_0; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_7_1; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_7_2; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_7_3; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_7_4; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_7_5; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_7_6; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_7_7; // @[stationary_dpe.scala 32:31]
  wire [15:0] _GEN_0 = count == 32'h0 ? io_Stationary_matrix_0_0 : Station2_0_0; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_1 = count == 32'h0 ? io_Stationary_matrix_0_1 : Station2_0_1; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_2 = count == 32'h0 ? io_Stationary_matrix_0_2 : Station2_0_2; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_3 = count == 32'h0 ? io_Stationary_matrix_0_3 : Station2_0_3; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_4 = count == 32'h0 ? io_Stationary_matrix_0_4 : Station2_0_4; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_5 = count == 32'h0 ? io_Stationary_matrix_0_5 : Station2_0_5; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_6 = count == 32'h0 ? io_Stationary_matrix_0_6 : Station2_0_6; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_7 = count == 32'h0 ? io_Stationary_matrix_0_7 : Station2_0_7; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_8 = count == 32'h0 ? io_Stationary_matrix_1_0 : Station2_1_0; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_9 = count == 32'h0 ? io_Stationary_matrix_1_1 : Station2_1_1; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_10 = count == 32'h0 ? io_Stationary_matrix_1_2 : Station2_1_2; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_11 = count == 32'h0 ? io_Stationary_matrix_1_3 : Station2_1_3; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_12 = count == 32'h0 ? io_Stationary_matrix_1_4 : Station2_1_4; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_13 = count == 32'h0 ? io_Stationary_matrix_1_5 : Station2_1_5; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_14 = count == 32'h0 ? io_Stationary_matrix_1_6 : Station2_1_6; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_15 = count == 32'h0 ? io_Stationary_matrix_1_7 : Station2_1_7; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_16 = count == 32'h0 ? io_Stationary_matrix_2_0 : Station2_2_0; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_17 = count == 32'h0 ? io_Stationary_matrix_2_1 : Station2_2_1; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_18 = count == 32'h0 ? io_Stationary_matrix_2_2 : Station2_2_2; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_19 = count == 32'h0 ? io_Stationary_matrix_2_3 : Station2_2_3; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_20 = count == 32'h0 ? io_Stationary_matrix_2_4 : Station2_2_4; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_21 = count == 32'h0 ? io_Stationary_matrix_2_5 : Station2_2_5; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_22 = count == 32'h0 ? io_Stationary_matrix_2_6 : Station2_2_6; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_23 = count == 32'h0 ? io_Stationary_matrix_2_7 : Station2_2_7; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_24 = count == 32'h0 ? io_Stationary_matrix_3_0 : Station2_3_0; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_25 = count == 32'h0 ? io_Stationary_matrix_3_1 : Station2_3_1; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_26 = count == 32'h0 ? io_Stationary_matrix_3_2 : Station2_3_2; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_27 = count == 32'h0 ? io_Stationary_matrix_3_3 : Station2_3_3; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_28 = count == 32'h0 ? io_Stationary_matrix_3_4 : Station2_3_4; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_29 = count == 32'h0 ? io_Stationary_matrix_3_5 : Station2_3_5; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_30 = count == 32'h0 ? io_Stationary_matrix_3_6 : Station2_3_6; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_31 = count == 32'h0 ? io_Stationary_matrix_3_7 : Station2_3_7; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_32 = count == 32'h0 ? io_Stationary_matrix_4_0 : Station2_4_0; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_33 = count == 32'h0 ? io_Stationary_matrix_4_1 : Station2_4_1; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_34 = count == 32'h0 ? io_Stationary_matrix_4_2 : Station2_4_2; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_35 = count == 32'h0 ? io_Stationary_matrix_4_3 : Station2_4_3; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_36 = count == 32'h0 ? io_Stationary_matrix_4_4 : Station2_4_4; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_37 = count == 32'h0 ? io_Stationary_matrix_4_5 : Station2_4_5; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_38 = count == 32'h0 ? io_Stationary_matrix_4_6 : Station2_4_6; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_39 = count == 32'h0 ? io_Stationary_matrix_4_7 : Station2_4_7; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_40 = count == 32'h0 ? io_Stationary_matrix_5_0 : Station2_5_0; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_41 = count == 32'h0 ? io_Stationary_matrix_5_1 : Station2_5_1; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_42 = count == 32'h0 ? io_Stationary_matrix_5_2 : Station2_5_2; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_43 = count == 32'h0 ? io_Stationary_matrix_5_3 : Station2_5_3; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_44 = count == 32'h0 ? io_Stationary_matrix_5_4 : Station2_5_4; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_45 = count == 32'h0 ? io_Stationary_matrix_5_5 : Station2_5_5; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_46 = count == 32'h0 ? io_Stationary_matrix_5_6 : Station2_5_6; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_47 = count == 32'h0 ? io_Stationary_matrix_5_7 : Station2_5_7; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_48 = count == 32'h0 ? io_Stationary_matrix_6_0 : Station2_6_0; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_49 = count == 32'h0 ? io_Stationary_matrix_6_1 : Station2_6_1; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_50 = count == 32'h0 ? io_Stationary_matrix_6_2 : Station2_6_2; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_51 = count == 32'h0 ? io_Stationary_matrix_6_3 : Station2_6_3; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_52 = count == 32'h0 ? io_Stationary_matrix_6_4 : Station2_6_4; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_53 = count == 32'h0 ? io_Stationary_matrix_6_5 : Station2_6_5; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_54 = count == 32'h0 ? io_Stationary_matrix_6_6 : Station2_6_6; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_55 = count == 32'h0 ? io_Stationary_matrix_6_7 : Station2_6_7; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_56 = count == 32'h0 ? io_Stationary_matrix_7_0 : Station2_7_0; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_57 = count == 32'h0 ? io_Stationary_matrix_7_1 : Station2_7_1; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_58 = count == 32'h0 ? io_Stationary_matrix_7_2 : Station2_7_2; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_59 = count == 32'h0 ? io_Stationary_matrix_7_3 : Station2_7_3; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_60 = count == 32'h0 ? io_Stationary_matrix_7_4 : Station2_7_4; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_61 = count == 32'h0 ? io_Stationary_matrix_7_5 : Station2_7_5; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_62 = count == 32'h0 ? io_Stationary_matrix_7_6 : Station2_7_6; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_63 = count == 32'h0 ? io_Stationary_matrix_7_7 : Station2_7_7; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_64 = count == 32'h8 ? Station2_0_0 : Station3_0_0; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_65 = count == 32'h8 ? Station2_0_1 : Station3_0_1; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_66 = count == 32'h8 ? Station2_0_2 : Station3_0_2; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_67 = count == 32'h8 ? Station2_0_3 : Station3_0_3; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_68 = count == 32'h8 ? Station2_0_4 : Station3_0_4; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_69 = count == 32'h8 ? Station2_0_5 : Station3_0_5; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_70 = count == 32'h8 ? Station2_0_6 : Station3_0_6; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_71 = count == 32'h8 ? Station2_0_7 : Station3_0_7; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_72 = count == 32'h8 ? Station2_1_0 : Station3_1_0; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_73 = count == 32'h8 ? Station2_1_1 : Station3_1_1; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_74 = count == 32'h8 ? Station2_1_2 : Station3_1_2; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_75 = count == 32'h8 ? Station2_1_3 : Station3_1_3; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_76 = count == 32'h8 ? Station2_1_4 : Station3_1_4; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_77 = count == 32'h8 ? Station2_1_5 : Station3_1_5; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_78 = count == 32'h8 ? Station2_1_6 : Station3_1_6; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_79 = count == 32'h8 ? Station2_1_7 : Station3_1_7; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_80 = count == 32'h8 ? Station2_2_0 : Station3_2_0; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_81 = count == 32'h8 ? Station2_2_1 : Station3_2_1; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_82 = count == 32'h8 ? Station2_2_2 : Station3_2_2; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_83 = count == 32'h8 ? Station2_2_3 : Station3_2_3; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_84 = count == 32'h8 ? Station2_2_4 : Station3_2_4; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_85 = count == 32'h8 ? Station2_2_5 : Station3_2_5; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_86 = count == 32'h8 ? Station2_2_6 : Station3_2_6; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_87 = count == 32'h8 ? Station2_2_7 : Station3_2_7; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_88 = count == 32'h8 ? Station2_3_0 : Station3_3_0; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_89 = count == 32'h8 ? Station2_3_1 : Station3_3_1; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_90 = count == 32'h8 ? Station2_3_2 : Station3_3_2; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_91 = count == 32'h8 ? Station2_3_3 : Station3_3_3; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_92 = count == 32'h8 ? Station2_3_4 : Station3_3_4; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_93 = count == 32'h8 ? Station2_3_5 : Station3_3_5; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_94 = count == 32'h8 ? Station2_3_6 : Station3_3_6; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_95 = count == 32'h8 ? Station2_3_7 : Station3_3_7; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_96 = count == 32'h8 ? Station2_4_0 : Station3_4_0; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_97 = count == 32'h8 ? Station2_4_1 : Station3_4_1; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_98 = count == 32'h8 ? Station2_4_2 : Station3_4_2; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_99 = count == 32'h8 ? Station2_4_3 : Station3_4_3; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_100 = count == 32'h8 ? Station2_4_4 : Station3_4_4; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_101 = count == 32'h8 ? Station2_4_5 : Station3_4_5; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_102 = count == 32'h8 ? Station2_4_6 : Station3_4_6; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_103 = count == 32'h8 ? Station2_4_7 : Station3_4_7; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_104 = count == 32'h8 ? Station2_5_0 : Station3_5_0; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_105 = count == 32'h8 ? Station2_5_1 : Station3_5_1; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_106 = count == 32'h8 ? Station2_5_2 : Station3_5_2; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_107 = count == 32'h8 ? Station2_5_3 : Station3_5_3; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_108 = count == 32'h8 ? Station2_5_4 : Station3_5_4; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_109 = count == 32'h8 ? Station2_5_5 : Station3_5_5; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_110 = count == 32'h8 ? Station2_5_6 : Station3_5_6; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_111 = count == 32'h8 ? Station2_5_7 : Station3_5_7; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_112 = count == 32'h8 ? Station2_6_0 : Station3_6_0; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_113 = count == 32'h8 ? Station2_6_1 : Station3_6_1; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_114 = count == 32'h8 ? Station2_6_2 : Station3_6_2; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_115 = count == 32'h8 ? Station2_6_3 : Station3_6_3; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_116 = count == 32'h8 ? Station2_6_4 : Station3_6_4; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_117 = count == 32'h8 ? Station2_6_5 : Station3_6_5; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_118 = count == 32'h8 ? Station2_6_6 : Station3_6_6; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_119 = count == 32'h8 ? Station2_6_7 : Station3_6_7; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_120 = count == 32'h8 ? Station2_7_0 : Station3_7_0; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_121 = count == 32'h8 ? Station2_7_1 : Station3_7_1; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_122 = count == 32'h8 ? Station2_7_2 : Station3_7_2; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_123 = count == 32'h8 ? Station2_7_3 : Station3_7_3; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_124 = count == 32'h8 ? Station2_7_4 : Station3_7_4; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_125 = count == 32'h8 ? Station2_7_5 : Station3_7_5; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_126 = count == 32'h8 ? Station2_7_6 : Station3_7_6; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_127 = count == 32'h8 ? Station2_7_7 : Station3_7_7; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_128 = count == 32'h10 ? Station3_0_0 : Station4_0_0; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_129 = count == 32'h10 ? Station3_0_1 : Station4_0_1; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_130 = count == 32'h10 ? Station3_0_2 : Station4_0_2; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_131 = count == 32'h10 ? Station3_0_3 : Station4_0_3; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_132 = count == 32'h10 ? Station3_0_4 : Station4_0_4; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_133 = count == 32'h10 ? Station3_0_5 : Station4_0_5; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_134 = count == 32'h10 ? Station3_0_6 : Station4_0_6; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_135 = count == 32'h10 ? Station3_0_7 : Station4_0_7; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_136 = count == 32'h10 ? Station3_1_0 : Station4_1_0; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_137 = count == 32'h10 ? Station3_1_1 : Station4_1_1; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_138 = count == 32'h10 ? Station3_1_2 : Station4_1_2; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_139 = count == 32'h10 ? Station3_1_3 : Station4_1_3; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_140 = count == 32'h10 ? Station3_1_4 : Station4_1_4; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_141 = count == 32'h10 ? Station3_1_5 : Station4_1_5; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_142 = count == 32'h10 ? Station3_1_6 : Station4_1_6; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_143 = count == 32'h10 ? Station3_1_7 : Station4_1_7; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_144 = count == 32'h10 ? Station3_2_0 : Station4_2_0; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_145 = count == 32'h10 ? Station3_2_1 : Station4_2_1; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_146 = count == 32'h10 ? Station3_2_2 : Station4_2_2; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_147 = count == 32'h10 ? Station3_2_3 : Station4_2_3; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_148 = count == 32'h10 ? Station3_2_4 : Station4_2_4; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_149 = count == 32'h10 ? Station3_2_5 : Station4_2_5; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_150 = count == 32'h10 ? Station3_2_6 : Station4_2_6; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_151 = count == 32'h10 ? Station3_2_7 : Station4_2_7; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_152 = count == 32'h10 ? Station3_3_0 : Station4_3_0; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_153 = count == 32'h10 ? Station3_3_1 : Station4_3_1; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_154 = count == 32'h10 ? Station3_3_2 : Station4_3_2; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_155 = count == 32'h10 ? Station3_3_3 : Station4_3_3; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_156 = count == 32'h10 ? Station3_3_4 : Station4_3_4; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_157 = count == 32'h10 ? Station3_3_5 : Station4_3_5; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_158 = count == 32'h10 ? Station3_3_6 : Station4_3_6; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_159 = count == 32'h10 ? Station3_3_7 : Station4_3_7; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_160 = count == 32'h10 ? Station3_4_0 : Station4_4_0; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_161 = count == 32'h10 ? Station3_4_1 : Station4_4_1; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_162 = count == 32'h10 ? Station3_4_2 : Station4_4_2; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_163 = count == 32'h10 ? Station3_4_3 : Station4_4_3; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_164 = count == 32'h10 ? Station3_4_4 : Station4_4_4; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_165 = count == 32'h10 ? Station3_4_5 : Station4_4_5; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_166 = count == 32'h10 ? Station3_4_6 : Station4_4_6; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_167 = count == 32'h10 ? Station3_4_7 : Station4_4_7; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_168 = count == 32'h10 ? Station3_5_0 : Station4_5_0; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_169 = count == 32'h10 ? Station3_5_1 : Station4_5_1; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_170 = count == 32'h10 ? Station3_5_2 : Station4_5_2; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_171 = count == 32'h10 ? Station3_5_3 : Station4_5_3; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_172 = count == 32'h10 ? Station3_5_4 : Station4_5_4; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_173 = count == 32'h10 ? Station3_5_5 : Station4_5_5; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_174 = count == 32'h10 ? Station3_5_6 : Station4_5_6; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_175 = count == 32'h10 ? Station3_5_7 : Station4_5_7; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_176 = count == 32'h10 ? Station3_6_0 : Station4_6_0; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_177 = count == 32'h10 ? Station3_6_1 : Station4_6_1; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_178 = count == 32'h10 ? Station3_6_2 : Station4_6_2; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_179 = count == 32'h10 ? Station3_6_3 : Station4_6_3; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_180 = count == 32'h10 ? Station3_6_4 : Station4_6_4; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_181 = count == 32'h10 ? Station3_6_5 : Station4_6_5; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_182 = count == 32'h10 ? Station3_6_6 : Station4_6_6; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_183 = count == 32'h10 ? Station3_6_7 : Station4_6_7; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_184 = count == 32'h10 ? Station3_7_0 : Station4_7_0; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_185 = count == 32'h10 ? Station3_7_1 : Station4_7_1; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_186 = count == 32'h10 ? Station3_7_2 : Station4_7_2; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_187 = count == 32'h10 ? Station3_7_3 : Station4_7_3; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_188 = count == 32'h10 ? Station3_7_4 : Station4_7_4; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_189 = count == 32'h10 ? Station3_7_5 : Station4_7_5; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_190 = count == 32'h10 ? Station3_7_6 : Station4_7_6; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_191 = count == 32'h10 ? Station3_7_7 : Station4_7_7; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_192 = count == 32'h18 ? Station4_0_0 : Station5_0_0; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_193 = count == 32'h18 ? Station4_0_1 : Station5_0_1; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_194 = count == 32'h18 ? Station4_0_2 : Station5_0_2; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_195 = count == 32'h18 ? Station4_0_3 : Station5_0_3; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_196 = count == 32'h18 ? Station4_0_4 : Station5_0_4; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_197 = count == 32'h18 ? Station4_0_5 : Station5_0_5; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_198 = count == 32'h18 ? Station4_0_6 : Station5_0_6; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_199 = count == 32'h18 ? Station4_0_7 : Station5_0_7; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_200 = count == 32'h18 ? Station4_1_0 : Station5_1_0; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_201 = count == 32'h18 ? Station4_1_1 : Station5_1_1; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_202 = count == 32'h18 ? Station4_1_2 : Station5_1_2; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_203 = count == 32'h18 ? Station4_1_3 : Station5_1_3; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_204 = count == 32'h18 ? Station4_1_4 : Station5_1_4; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_205 = count == 32'h18 ? Station4_1_5 : Station5_1_5; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_206 = count == 32'h18 ? Station4_1_6 : Station5_1_6; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_207 = count == 32'h18 ? Station4_1_7 : Station5_1_7; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_208 = count == 32'h18 ? Station4_2_0 : Station5_2_0; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_209 = count == 32'h18 ? Station4_2_1 : Station5_2_1; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_210 = count == 32'h18 ? Station4_2_2 : Station5_2_2; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_211 = count == 32'h18 ? Station4_2_3 : Station5_2_3; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_212 = count == 32'h18 ? Station4_2_4 : Station5_2_4; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_213 = count == 32'h18 ? Station4_2_5 : Station5_2_5; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_214 = count == 32'h18 ? Station4_2_6 : Station5_2_6; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_215 = count == 32'h18 ? Station4_2_7 : Station5_2_7; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_216 = count == 32'h18 ? Station4_3_0 : Station5_3_0; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_217 = count == 32'h18 ? Station4_3_1 : Station5_3_1; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_218 = count == 32'h18 ? Station4_3_2 : Station5_3_2; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_219 = count == 32'h18 ? Station4_3_3 : Station5_3_3; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_220 = count == 32'h18 ? Station4_3_4 : Station5_3_4; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_221 = count == 32'h18 ? Station4_3_5 : Station5_3_5; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_222 = count == 32'h18 ? Station4_3_6 : Station5_3_6; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_223 = count == 32'h18 ? Station4_3_7 : Station5_3_7; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_224 = count == 32'h18 ? Station4_4_0 : Station5_4_0; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_225 = count == 32'h18 ? Station4_4_1 : Station5_4_1; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_226 = count == 32'h18 ? Station4_4_2 : Station5_4_2; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_227 = count == 32'h18 ? Station4_4_3 : Station5_4_3; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_228 = count == 32'h18 ? Station4_4_4 : Station5_4_4; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_229 = count == 32'h18 ? Station4_4_5 : Station5_4_5; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_230 = count == 32'h18 ? Station4_4_6 : Station5_4_6; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_231 = count == 32'h18 ? Station4_4_7 : Station5_4_7; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_232 = count == 32'h18 ? Station4_5_0 : Station5_5_0; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_233 = count == 32'h18 ? Station4_5_1 : Station5_5_1; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_234 = count == 32'h18 ? Station4_5_2 : Station5_5_2; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_235 = count == 32'h18 ? Station4_5_3 : Station5_5_3; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_236 = count == 32'h18 ? Station4_5_4 : Station5_5_4; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_237 = count == 32'h18 ? Station4_5_5 : Station5_5_5; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_238 = count == 32'h18 ? Station4_5_6 : Station5_5_6; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_239 = count == 32'h18 ? Station4_5_7 : Station5_5_7; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_240 = count == 32'h18 ? Station4_6_0 : Station5_6_0; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_241 = count == 32'h18 ? Station4_6_1 : Station5_6_1; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_242 = count == 32'h18 ? Station4_6_2 : Station5_6_2; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_243 = count == 32'h18 ? Station4_6_3 : Station5_6_3; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_244 = count == 32'h18 ? Station4_6_4 : Station5_6_4; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_245 = count == 32'h18 ? Station4_6_5 : Station5_6_5; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_246 = count == 32'h18 ? Station4_6_6 : Station5_6_6; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_247 = count == 32'h18 ? Station4_6_7 : Station5_6_7; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_248 = count == 32'h18 ? Station4_7_0 : Station5_7_0; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_249 = count == 32'h18 ? Station4_7_1 : Station5_7_1; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_250 = count == 32'h18 ? Station4_7_2 : Station5_7_2; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_251 = count == 32'h18 ? Station4_7_3 : Station5_7_3; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_252 = count == 32'h18 ? Station4_7_4 : Station5_7_4; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_253 = count == 32'h18 ? Station4_7_5 : Station5_7_5; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_254 = count == 32'h18 ? Station4_7_6 : Station5_7_6; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_255 = count == 32'h18 ? Station4_7_7 : Station5_7_7; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_256 = count == 32'h20 ? Station5_0_0 : Station6_0_0; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_257 = count == 32'h20 ? Station5_0_1 : Station6_0_1; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_258 = count == 32'h20 ? Station5_0_2 : Station6_0_2; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_259 = count == 32'h20 ? Station5_0_3 : Station6_0_3; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_260 = count == 32'h20 ? Station5_0_4 : Station6_0_4; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_261 = count == 32'h20 ? Station5_0_5 : Station6_0_5; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_262 = count == 32'h20 ? Station5_0_6 : Station6_0_6; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_263 = count == 32'h20 ? Station5_0_7 : Station6_0_7; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_264 = count == 32'h20 ? Station5_1_0 : Station6_1_0; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_265 = count == 32'h20 ? Station5_1_1 : Station6_1_1; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_266 = count == 32'h20 ? Station5_1_2 : Station6_1_2; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_267 = count == 32'h20 ? Station5_1_3 : Station6_1_3; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_268 = count == 32'h20 ? Station5_1_4 : Station6_1_4; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_269 = count == 32'h20 ? Station5_1_5 : Station6_1_5; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_270 = count == 32'h20 ? Station5_1_6 : Station6_1_6; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_271 = count == 32'h20 ? Station5_1_7 : Station6_1_7; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_272 = count == 32'h20 ? Station5_2_0 : Station6_2_0; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_273 = count == 32'h20 ? Station5_2_1 : Station6_2_1; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_274 = count == 32'h20 ? Station5_2_2 : Station6_2_2; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_275 = count == 32'h20 ? Station5_2_3 : Station6_2_3; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_276 = count == 32'h20 ? Station5_2_4 : Station6_2_4; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_277 = count == 32'h20 ? Station5_2_5 : Station6_2_5; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_278 = count == 32'h20 ? Station5_2_6 : Station6_2_6; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_279 = count == 32'h20 ? Station5_2_7 : Station6_2_7; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_280 = count == 32'h20 ? Station5_3_0 : Station6_3_0; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_281 = count == 32'h20 ? Station5_3_1 : Station6_3_1; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_282 = count == 32'h20 ? Station5_3_2 : Station6_3_2; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_283 = count == 32'h20 ? Station5_3_3 : Station6_3_3; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_284 = count == 32'h20 ? Station5_3_4 : Station6_3_4; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_285 = count == 32'h20 ? Station5_3_5 : Station6_3_5; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_286 = count == 32'h20 ? Station5_3_6 : Station6_3_6; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_287 = count == 32'h20 ? Station5_3_7 : Station6_3_7; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_288 = count == 32'h20 ? Station5_4_0 : Station6_4_0; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_289 = count == 32'h20 ? Station5_4_1 : Station6_4_1; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_290 = count == 32'h20 ? Station5_4_2 : Station6_4_2; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_291 = count == 32'h20 ? Station5_4_3 : Station6_4_3; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_292 = count == 32'h20 ? Station5_4_4 : Station6_4_4; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_293 = count == 32'h20 ? Station5_4_5 : Station6_4_5; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_294 = count == 32'h20 ? Station5_4_6 : Station6_4_6; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_295 = count == 32'h20 ? Station5_4_7 : Station6_4_7; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_296 = count == 32'h20 ? Station5_5_0 : Station6_5_0; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_297 = count == 32'h20 ? Station5_5_1 : Station6_5_1; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_298 = count == 32'h20 ? Station5_5_2 : Station6_5_2; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_299 = count == 32'h20 ? Station5_5_3 : Station6_5_3; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_300 = count == 32'h20 ? Station5_5_4 : Station6_5_4; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_301 = count == 32'h20 ? Station5_5_5 : Station6_5_5; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_302 = count == 32'h20 ? Station5_5_6 : Station6_5_6; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_303 = count == 32'h20 ? Station5_5_7 : Station6_5_7; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_304 = count == 32'h20 ? Station5_6_0 : Station6_6_0; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_305 = count == 32'h20 ? Station5_6_1 : Station6_6_1; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_306 = count == 32'h20 ? Station5_6_2 : Station6_6_2; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_307 = count == 32'h20 ? Station5_6_3 : Station6_6_3; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_308 = count == 32'h20 ? Station5_6_4 : Station6_6_4; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_309 = count == 32'h20 ? Station5_6_5 : Station6_6_5; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_310 = count == 32'h20 ? Station5_6_6 : Station6_6_6; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_311 = count == 32'h20 ? Station5_6_7 : Station6_6_7; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_312 = count == 32'h20 ? Station5_7_0 : Station6_7_0; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_313 = count == 32'h20 ? Station5_7_1 : Station6_7_1; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_314 = count == 32'h20 ? Station5_7_2 : Station6_7_2; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_315 = count == 32'h20 ? Station5_7_3 : Station6_7_3; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_316 = count == 32'h20 ? Station5_7_4 : Station6_7_4; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_317 = count == 32'h20 ? Station5_7_5 : Station6_7_5; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_318 = count == 32'h20 ? Station5_7_6 : Station6_7_6; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_319 = count == 32'h20 ? Station5_7_7 : Station6_7_7; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_320 = count == 32'h28 ? Station6_0_0 : Station7_0_0; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_321 = count == 32'h28 ? Station6_0_1 : Station7_0_1; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_322 = count == 32'h28 ? Station6_0_2 : Station7_0_2; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_323 = count == 32'h28 ? Station6_0_3 : Station7_0_3; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_324 = count == 32'h28 ? Station6_0_4 : Station7_0_4; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_325 = count == 32'h28 ? Station6_0_5 : Station7_0_5; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_326 = count == 32'h28 ? Station6_0_6 : Station7_0_6; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_327 = count == 32'h28 ? Station6_0_7 : Station7_0_7; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_328 = count == 32'h28 ? Station6_1_0 : Station7_1_0; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_329 = count == 32'h28 ? Station6_1_1 : Station7_1_1; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_330 = count == 32'h28 ? Station6_1_2 : Station7_1_2; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_331 = count == 32'h28 ? Station6_1_3 : Station7_1_3; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_332 = count == 32'h28 ? Station6_1_4 : Station7_1_4; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_333 = count == 32'h28 ? Station6_1_5 : Station7_1_5; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_334 = count == 32'h28 ? Station6_1_6 : Station7_1_6; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_335 = count == 32'h28 ? Station6_1_7 : Station7_1_7; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_336 = count == 32'h28 ? Station6_2_0 : Station7_2_0; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_337 = count == 32'h28 ? Station6_2_1 : Station7_2_1; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_338 = count == 32'h28 ? Station6_2_2 : Station7_2_2; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_339 = count == 32'h28 ? Station6_2_3 : Station7_2_3; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_340 = count == 32'h28 ? Station6_2_4 : Station7_2_4; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_341 = count == 32'h28 ? Station6_2_5 : Station7_2_5; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_342 = count == 32'h28 ? Station6_2_6 : Station7_2_6; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_343 = count == 32'h28 ? Station6_2_7 : Station7_2_7; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_344 = count == 32'h28 ? Station6_3_0 : Station7_3_0; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_345 = count == 32'h28 ? Station6_3_1 : Station7_3_1; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_346 = count == 32'h28 ? Station6_3_2 : Station7_3_2; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_347 = count == 32'h28 ? Station6_3_3 : Station7_3_3; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_348 = count == 32'h28 ? Station6_3_4 : Station7_3_4; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_349 = count == 32'h28 ? Station6_3_5 : Station7_3_5; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_350 = count == 32'h28 ? Station6_3_6 : Station7_3_6; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_351 = count == 32'h28 ? Station6_3_7 : Station7_3_7; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_352 = count == 32'h28 ? Station6_4_0 : Station7_4_0; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_353 = count == 32'h28 ? Station6_4_1 : Station7_4_1; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_354 = count == 32'h28 ? Station6_4_2 : Station7_4_2; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_355 = count == 32'h28 ? Station6_4_3 : Station7_4_3; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_356 = count == 32'h28 ? Station6_4_4 : Station7_4_4; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_357 = count == 32'h28 ? Station6_4_5 : Station7_4_5; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_358 = count == 32'h28 ? Station6_4_6 : Station7_4_6; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_359 = count == 32'h28 ? Station6_4_7 : Station7_4_7; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_360 = count == 32'h28 ? Station6_5_0 : Station7_5_0; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_361 = count == 32'h28 ? Station6_5_1 : Station7_5_1; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_362 = count == 32'h28 ? Station6_5_2 : Station7_5_2; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_363 = count == 32'h28 ? Station6_5_3 : Station7_5_3; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_364 = count == 32'h28 ? Station6_5_4 : Station7_5_4; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_365 = count == 32'h28 ? Station6_5_5 : Station7_5_5; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_366 = count == 32'h28 ? Station6_5_6 : Station7_5_6; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_367 = count == 32'h28 ? Station6_5_7 : Station7_5_7; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_368 = count == 32'h28 ? Station6_6_0 : Station7_6_0; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_369 = count == 32'h28 ? Station6_6_1 : Station7_6_1; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_370 = count == 32'h28 ? Station6_6_2 : Station7_6_2; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_371 = count == 32'h28 ? Station6_6_3 : Station7_6_3; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_372 = count == 32'h28 ? Station6_6_4 : Station7_6_4; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_373 = count == 32'h28 ? Station6_6_5 : Station7_6_5; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_374 = count == 32'h28 ? Station6_6_6 : Station7_6_6; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_375 = count == 32'h28 ? Station6_6_7 : Station7_6_7; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_376 = count == 32'h28 ? Station6_7_0 : Station7_7_0; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_377 = count == 32'h28 ? Station6_7_1 : Station7_7_1; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_378 = count == 32'h28 ? Station6_7_2 : Station7_7_2; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_379 = count == 32'h28 ? Station6_7_3 : Station7_7_3; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_380 = count == 32'h28 ? Station6_7_4 : Station7_7_4; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_381 = count == 32'h28 ? Station6_7_5 : Station7_7_5; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_382 = count == 32'h28 ? Station6_7_6 : Station7_7_6; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_383 = count == 32'h28 ? Station6_7_7 : Station7_7_7; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_384 = count == 32'h30 ? Station7_0_0 : Station8_0_0; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_385 = count == 32'h30 ? Station7_0_1 : Station8_0_1; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_386 = count == 32'h30 ? Station7_0_2 : Station8_0_2; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_387 = count == 32'h30 ? Station7_0_3 : Station8_0_3; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_388 = count == 32'h30 ? Station7_0_4 : Station8_0_4; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_389 = count == 32'h30 ? Station7_0_5 : Station8_0_5; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_390 = count == 32'h30 ? Station7_0_6 : Station8_0_6; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_391 = count == 32'h30 ? Station7_0_7 : Station8_0_7; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_392 = count == 32'h30 ? Station7_1_0 : Station8_1_0; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_393 = count == 32'h30 ? Station7_1_1 : Station8_1_1; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_394 = count == 32'h30 ? Station7_1_2 : Station8_1_2; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_395 = count == 32'h30 ? Station7_1_3 : Station8_1_3; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_396 = count == 32'h30 ? Station7_1_4 : Station8_1_4; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_397 = count == 32'h30 ? Station7_1_5 : Station8_1_5; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_398 = count == 32'h30 ? Station7_1_6 : Station8_1_6; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_399 = count == 32'h30 ? Station7_1_7 : Station8_1_7; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_400 = count == 32'h30 ? Station7_2_0 : Station8_2_0; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_401 = count == 32'h30 ? Station7_2_1 : Station8_2_1; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_402 = count == 32'h30 ? Station7_2_2 : Station8_2_2; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_403 = count == 32'h30 ? Station7_2_3 : Station8_2_3; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_404 = count == 32'h30 ? Station7_2_4 : Station8_2_4; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_405 = count == 32'h30 ? Station7_2_5 : Station8_2_5; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_406 = count == 32'h30 ? Station7_2_6 : Station8_2_6; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_407 = count == 32'h30 ? Station7_2_7 : Station8_2_7; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_408 = count == 32'h30 ? Station7_3_0 : Station8_3_0; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_409 = count == 32'h30 ? Station7_3_1 : Station8_3_1; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_410 = count == 32'h30 ? Station7_3_2 : Station8_3_2; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_411 = count == 32'h30 ? Station7_3_3 : Station8_3_3; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_412 = count == 32'h30 ? Station7_3_4 : Station8_3_4; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_413 = count == 32'h30 ? Station7_3_5 : Station8_3_5; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_414 = count == 32'h30 ? Station7_3_6 : Station8_3_6; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_415 = count == 32'h30 ? Station7_3_7 : Station8_3_7; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_416 = count == 32'h30 ? Station7_4_0 : Station8_4_0; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_417 = count == 32'h30 ? Station7_4_1 : Station8_4_1; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_418 = count == 32'h30 ? Station7_4_2 : Station8_4_2; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_419 = count == 32'h30 ? Station7_4_3 : Station8_4_3; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_420 = count == 32'h30 ? Station7_4_4 : Station8_4_4; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_421 = count == 32'h30 ? Station7_4_5 : Station8_4_5; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_422 = count == 32'h30 ? Station7_4_6 : Station8_4_6; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_423 = count == 32'h30 ? Station7_4_7 : Station8_4_7; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_424 = count == 32'h30 ? Station7_5_0 : Station8_5_0; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_425 = count == 32'h30 ? Station7_5_1 : Station8_5_1; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_426 = count == 32'h30 ? Station7_5_2 : Station8_5_2; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_427 = count == 32'h30 ? Station7_5_3 : Station8_5_3; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_428 = count == 32'h30 ? Station7_5_4 : Station8_5_4; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_429 = count == 32'h30 ? Station7_5_5 : Station8_5_5; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_430 = count == 32'h30 ? Station7_5_6 : Station8_5_6; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_431 = count == 32'h30 ? Station7_5_7 : Station8_5_7; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_432 = count == 32'h30 ? Station7_6_0 : Station8_6_0; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_433 = count == 32'h30 ? Station7_6_1 : Station8_6_1; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_434 = count == 32'h30 ? Station7_6_2 : Station8_6_2; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_435 = count == 32'h30 ? Station7_6_3 : Station8_6_3; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_436 = count == 32'h30 ? Station7_6_4 : Station8_6_4; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_437 = count == 32'h30 ? Station7_6_5 : Station8_6_5; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_438 = count == 32'h30 ? Station7_6_6 : Station8_6_6; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_439 = count == 32'h30 ? Station7_6_7 : Station8_6_7; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_440 = count == 32'h30 ? Station7_7_0 : Station8_7_0; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_441 = count == 32'h30 ? Station7_7_1 : Station8_7_1; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_442 = count == 32'h30 ? Station7_7_2 : Station8_7_2; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_443 = count == 32'h30 ? Station7_7_3 : Station8_7_3; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_444 = count == 32'h30 ? Station7_7_4 : Station8_7_4; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_445 = count == 32'h30 ? Station7_7_5 : Station8_7_5; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_446 = count == 32'h30 ? Station7_7_6 : Station8_7_6; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_447 = count == 32'h30 ? Station7_7_7 : Station8_7_7; // @[stationary_dpe.scala 70:27 71:15 32:31]
  reg [31:0] i; // @[stationary_dpe.scala 79:20]
  reg [31:0] j; // @[stationary_dpe.scala 80:20]
  wire  valid = count >= 32'h8; // @[stationary_dpe.scala 190:17]
  wire  _GEN_2264 = 3'h0 == i[2:0]; // @[stationary_dpe.scala 94:{43,43}]
  wire  _GEN_2265 = 3'h1 == j[2:0]; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_449 = 3'h0 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_0_1 : io_Stationary_matrix_0_0; // @[stationary_dpe.scala 94:{43,43}]
  wire  _GEN_2267 = 3'h2 == j[2:0]; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_450 = 3'h0 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_0_2 : _GEN_449; // @[stationary_dpe.scala 94:{43,43}]
  wire  _GEN_2269 = 3'h3 == j[2:0]; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_451 = 3'h0 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_0_3 : _GEN_450; // @[stationary_dpe.scala 94:{43,43}]
  wire  _GEN_2271 = 3'h4 == j[2:0]; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_452 = 3'h0 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_0_4 : _GEN_451; // @[stationary_dpe.scala 94:{43,43}]
  wire  _GEN_2273 = 3'h5 == j[2:0]; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_453 = 3'h0 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_0_5 : _GEN_452; // @[stationary_dpe.scala 94:{43,43}]
  wire  _GEN_2275 = 3'h6 == j[2:0]; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_454 = 3'h0 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_0_6 : _GEN_453; // @[stationary_dpe.scala 94:{43,43}]
  wire  _GEN_2277 = 3'h7 == j[2:0]; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_455 = 3'h0 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_0_7 : _GEN_454; // @[stationary_dpe.scala 94:{43,43}]
  wire  _GEN_2278 = 3'h1 == i[2:0]; // @[stationary_dpe.scala 94:{43,43}]
  wire  _GEN_2279 = 3'h0 == j[2:0]; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_456 = 3'h1 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_1_0 : _GEN_455; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_457 = 3'h1 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_1_1 : _GEN_456; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_458 = 3'h1 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_1_2 : _GEN_457; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_459 = 3'h1 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_1_3 : _GEN_458; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_460 = 3'h1 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_1_4 : _GEN_459; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_461 = 3'h1 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_1_5 : _GEN_460; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_462 = 3'h1 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_1_6 : _GEN_461; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_463 = 3'h1 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_1_7 : _GEN_462; // @[stationary_dpe.scala 94:{43,43}]
  wire  _GEN_2294 = 3'h2 == i[2:0]; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_464 = 3'h2 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_2_0 : _GEN_463; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_465 = 3'h2 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_2_1 : _GEN_464; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_466 = 3'h2 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_2_2 : _GEN_465; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_467 = 3'h2 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_2_3 : _GEN_466; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_468 = 3'h2 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_2_4 : _GEN_467; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_469 = 3'h2 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_2_5 : _GEN_468; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_470 = 3'h2 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_2_6 : _GEN_469; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_471 = 3'h2 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_2_7 : _GEN_470; // @[stationary_dpe.scala 94:{43,43}]
  wire  _GEN_2310 = 3'h3 == i[2:0]; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_472 = 3'h3 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_3_0 : _GEN_471; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_473 = 3'h3 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_3_1 : _GEN_472; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_474 = 3'h3 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_3_2 : _GEN_473; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_475 = 3'h3 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_3_3 : _GEN_474; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_476 = 3'h3 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_3_4 : _GEN_475; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_477 = 3'h3 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_3_5 : _GEN_476; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_478 = 3'h3 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_3_6 : _GEN_477; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_479 = 3'h3 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_3_7 : _GEN_478; // @[stationary_dpe.scala 94:{43,43}]
  wire  _GEN_2326 = 3'h4 == i[2:0]; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_480 = 3'h4 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_4_0 : _GEN_479; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_481 = 3'h4 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_4_1 : _GEN_480; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_482 = 3'h4 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_4_2 : _GEN_481; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_483 = 3'h4 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_4_3 : _GEN_482; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_484 = 3'h4 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_4_4 : _GEN_483; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_485 = 3'h4 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_4_5 : _GEN_484; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_486 = 3'h4 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_4_6 : _GEN_485; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_487 = 3'h4 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_4_7 : _GEN_486; // @[stationary_dpe.scala 94:{43,43}]
  wire  _GEN_2342 = 3'h5 == i[2:0]; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_488 = 3'h5 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_5_0 : _GEN_487; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_489 = 3'h5 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_5_1 : _GEN_488; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_490 = 3'h5 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_5_2 : _GEN_489; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_491 = 3'h5 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_5_3 : _GEN_490; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_492 = 3'h5 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_5_4 : _GEN_491; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_493 = 3'h5 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_5_5 : _GEN_492; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_494 = 3'h5 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_5_6 : _GEN_493; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_495 = 3'h5 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_5_7 : _GEN_494; // @[stationary_dpe.scala 94:{43,43}]
  wire  _GEN_2358 = 3'h6 == i[2:0]; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_496 = 3'h6 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_6_0 : _GEN_495; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_497 = 3'h6 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_6_1 : _GEN_496; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_498 = 3'h6 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_6_2 : _GEN_497; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_499 = 3'h6 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_6_3 : _GEN_498; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_500 = 3'h6 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_6_4 : _GEN_499; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_501 = 3'h6 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_6_5 : _GEN_500; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_502 = 3'h6 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_6_6 : _GEN_501; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_503 = 3'h6 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_6_7 : _GEN_502; // @[stationary_dpe.scala 94:{43,43}]
  wire  _GEN_2374 = 3'h7 == i[2:0]; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_504 = 3'h7 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_7_0 : _GEN_503; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_505 = 3'h7 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_7_1 : _GEN_504; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_506 = 3'h7 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_7_2 : _GEN_505; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_507 = 3'h7 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_7_3 : _GEN_506; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_508 = 3'h7 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_7_4 : _GEN_507; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_509 = 3'h7 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_7_5 : _GEN_508; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_510 = 3'h7 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_7_6 : _GEN_509; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_511 = 3'h7 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_7_7 : _GEN_510; // @[stationary_dpe.scala 94:{43,43}]
  wire [31:0] _count_T_1 = count + 32'h1; // @[stationary_dpe.scala 97:27]
  wire [31:0] _GEN_640 = _GEN_511 != 16'h0 ? _count_T_1 : count; // @[stationary_dpe.scala 94:51 97:18 23:27]
  wire [31:0] _GEN_705 = ~valid ? _GEN_640 : count; // @[stationary_dpe.scala 23:27 93:27]
  wire  valid1 = count >= 32'h10; // @[stationary_dpe.scala 194:18]
  wire [15:0] _GEN_707 = _GEN_2264 & _GEN_2265 ? Station2_0_1 : Station2_0_0; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_708 = _GEN_2264 & _GEN_2267 ? Station2_0_2 : _GEN_707; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_709 = _GEN_2264 & _GEN_2269 ? Station2_0_3 : _GEN_708; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_710 = _GEN_2264 & _GEN_2271 ? Station2_0_4 : _GEN_709; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_711 = _GEN_2264 & _GEN_2273 ? Station2_0_5 : _GEN_710; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_712 = _GEN_2264 & _GEN_2275 ? Station2_0_6 : _GEN_711; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_713 = _GEN_2264 & _GEN_2277 ? Station2_0_7 : _GEN_712; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_714 = _GEN_2278 & _GEN_2279 ? Station2_1_0 : _GEN_713; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_715 = _GEN_2278 & _GEN_2265 ? Station2_1_1 : _GEN_714; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_716 = _GEN_2278 & _GEN_2267 ? Station2_1_2 : _GEN_715; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_717 = _GEN_2278 & _GEN_2269 ? Station2_1_3 : _GEN_716; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_718 = _GEN_2278 & _GEN_2271 ? Station2_1_4 : _GEN_717; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_719 = _GEN_2278 & _GEN_2273 ? Station2_1_5 : _GEN_718; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_720 = _GEN_2278 & _GEN_2275 ? Station2_1_6 : _GEN_719; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_721 = _GEN_2278 & _GEN_2277 ? Station2_1_7 : _GEN_720; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_722 = _GEN_2294 & _GEN_2279 ? Station2_2_0 : _GEN_721; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_723 = _GEN_2294 & _GEN_2265 ? Station2_2_1 : _GEN_722; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_724 = _GEN_2294 & _GEN_2267 ? Station2_2_2 : _GEN_723; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_725 = _GEN_2294 & _GEN_2269 ? Station2_2_3 : _GEN_724; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_726 = _GEN_2294 & _GEN_2271 ? Station2_2_4 : _GEN_725; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_727 = _GEN_2294 & _GEN_2273 ? Station2_2_5 : _GEN_726; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_728 = _GEN_2294 & _GEN_2275 ? Station2_2_6 : _GEN_727; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_729 = _GEN_2294 & _GEN_2277 ? Station2_2_7 : _GEN_728; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_730 = _GEN_2310 & _GEN_2279 ? Station2_3_0 : _GEN_729; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_731 = _GEN_2310 & _GEN_2265 ? Station2_3_1 : _GEN_730; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_732 = _GEN_2310 & _GEN_2267 ? Station2_3_2 : _GEN_731; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_733 = _GEN_2310 & _GEN_2269 ? Station2_3_3 : _GEN_732; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_734 = _GEN_2310 & _GEN_2271 ? Station2_3_4 : _GEN_733; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_735 = _GEN_2310 & _GEN_2273 ? Station2_3_5 : _GEN_734; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_736 = _GEN_2310 & _GEN_2275 ? Station2_3_6 : _GEN_735; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_737 = _GEN_2310 & _GEN_2277 ? Station2_3_7 : _GEN_736; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_738 = _GEN_2326 & _GEN_2279 ? Station2_4_0 : _GEN_737; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_739 = _GEN_2326 & _GEN_2265 ? Station2_4_1 : _GEN_738; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_740 = _GEN_2326 & _GEN_2267 ? Station2_4_2 : _GEN_739; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_741 = _GEN_2326 & _GEN_2269 ? Station2_4_3 : _GEN_740; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_742 = _GEN_2326 & _GEN_2271 ? Station2_4_4 : _GEN_741; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_743 = _GEN_2326 & _GEN_2273 ? Station2_4_5 : _GEN_742; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_744 = _GEN_2326 & _GEN_2275 ? Station2_4_6 : _GEN_743; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_745 = _GEN_2326 & _GEN_2277 ? Station2_4_7 : _GEN_744; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_746 = _GEN_2342 & _GEN_2279 ? Station2_5_0 : _GEN_745; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_747 = _GEN_2342 & _GEN_2265 ? Station2_5_1 : _GEN_746; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_748 = _GEN_2342 & _GEN_2267 ? Station2_5_2 : _GEN_747; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_749 = _GEN_2342 & _GEN_2269 ? Station2_5_3 : _GEN_748; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_750 = _GEN_2342 & _GEN_2271 ? Station2_5_4 : _GEN_749; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_751 = _GEN_2342 & _GEN_2273 ? Station2_5_5 : _GEN_750; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_752 = _GEN_2342 & _GEN_2275 ? Station2_5_6 : _GEN_751; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_753 = _GEN_2342 & _GEN_2277 ? Station2_5_7 : _GEN_752; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_754 = _GEN_2358 & _GEN_2279 ? Station2_6_0 : _GEN_753; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_755 = _GEN_2358 & _GEN_2265 ? Station2_6_1 : _GEN_754; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_756 = _GEN_2358 & _GEN_2267 ? Station2_6_2 : _GEN_755; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_757 = _GEN_2358 & _GEN_2269 ? Station2_6_3 : _GEN_756; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_758 = _GEN_2358 & _GEN_2271 ? Station2_6_4 : _GEN_757; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_759 = _GEN_2358 & _GEN_2273 ? Station2_6_5 : _GEN_758; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_760 = _GEN_2358 & _GEN_2275 ? Station2_6_6 : _GEN_759; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_761 = _GEN_2358 & _GEN_2277 ? Station2_6_7 : _GEN_760; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_762 = _GEN_2374 & _GEN_2279 ? Station2_7_0 : _GEN_761; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_763 = _GEN_2374 & _GEN_2265 ? Station2_7_1 : _GEN_762; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_764 = _GEN_2374 & _GEN_2267 ? Station2_7_2 : _GEN_763; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_765 = _GEN_2374 & _GEN_2269 ? Station2_7_3 : _GEN_764; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_766 = _GEN_2374 & _GEN_2271 ? Station2_7_4 : _GEN_765; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_767 = _GEN_2374 & _GEN_2273 ? Station2_7_5 : _GEN_766; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_768 = _GEN_2374 & _GEN_2275 ? Station2_7_6 : _GEN_767; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_769 = _GEN_2374 & _GEN_2277 ? Station2_7_7 : _GEN_768; // @[stationary_dpe.scala 115:{31,31}]
  wire [31:0] _GEN_898 = _GEN_769 != 16'h0 ? _count_T_1 : _GEN_705; // @[stationary_dpe.scala 115:39 118:18]
  wire [31:0] _GEN_963 = ~valid1 ? _GEN_898 : _GEN_705; // @[stationary_dpe.scala 114:29]
  wire  valid2 = count >= 32'h18; // @[stationary_dpe.scala 198:17]
  wire [15:0] _GEN_965 = _GEN_2264 & _GEN_2265 ? Station3_0_1 : Station3_0_0; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_966 = _GEN_2264 & _GEN_2267 ? Station3_0_2 : _GEN_965; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_967 = _GEN_2264 & _GEN_2269 ? Station3_0_3 : _GEN_966; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_968 = _GEN_2264 & _GEN_2271 ? Station3_0_4 : _GEN_967; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_969 = _GEN_2264 & _GEN_2273 ? Station3_0_5 : _GEN_968; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_970 = _GEN_2264 & _GEN_2275 ? Station3_0_6 : _GEN_969; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_971 = _GEN_2264 & _GEN_2277 ? Station3_0_7 : _GEN_970; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_972 = _GEN_2278 & _GEN_2279 ? Station3_1_0 : _GEN_971; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_973 = _GEN_2278 & _GEN_2265 ? Station3_1_1 : _GEN_972; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_974 = _GEN_2278 & _GEN_2267 ? Station3_1_2 : _GEN_973; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_975 = _GEN_2278 & _GEN_2269 ? Station3_1_3 : _GEN_974; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_976 = _GEN_2278 & _GEN_2271 ? Station3_1_4 : _GEN_975; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_977 = _GEN_2278 & _GEN_2273 ? Station3_1_5 : _GEN_976; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_978 = _GEN_2278 & _GEN_2275 ? Station3_1_6 : _GEN_977; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_979 = _GEN_2278 & _GEN_2277 ? Station3_1_7 : _GEN_978; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_980 = _GEN_2294 & _GEN_2279 ? Station3_2_0 : _GEN_979; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_981 = _GEN_2294 & _GEN_2265 ? Station3_2_1 : _GEN_980; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_982 = _GEN_2294 & _GEN_2267 ? Station3_2_2 : _GEN_981; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_983 = _GEN_2294 & _GEN_2269 ? Station3_2_3 : _GEN_982; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_984 = _GEN_2294 & _GEN_2271 ? Station3_2_4 : _GEN_983; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_985 = _GEN_2294 & _GEN_2273 ? Station3_2_5 : _GEN_984; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_986 = _GEN_2294 & _GEN_2275 ? Station3_2_6 : _GEN_985; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_987 = _GEN_2294 & _GEN_2277 ? Station3_2_7 : _GEN_986; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_988 = _GEN_2310 & _GEN_2279 ? Station3_3_0 : _GEN_987; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_989 = _GEN_2310 & _GEN_2265 ? Station3_3_1 : _GEN_988; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_990 = _GEN_2310 & _GEN_2267 ? Station3_3_2 : _GEN_989; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_991 = _GEN_2310 & _GEN_2269 ? Station3_3_3 : _GEN_990; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_992 = _GEN_2310 & _GEN_2271 ? Station3_3_4 : _GEN_991; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_993 = _GEN_2310 & _GEN_2273 ? Station3_3_5 : _GEN_992; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_994 = _GEN_2310 & _GEN_2275 ? Station3_3_6 : _GEN_993; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_995 = _GEN_2310 & _GEN_2277 ? Station3_3_7 : _GEN_994; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_996 = _GEN_2326 & _GEN_2279 ? Station3_4_0 : _GEN_995; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_997 = _GEN_2326 & _GEN_2265 ? Station3_4_1 : _GEN_996; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_998 = _GEN_2326 & _GEN_2267 ? Station3_4_2 : _GEN_997; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_999 = _GEN_2326 & _GEN_2269 ? Station3_4_3 : _GEN_998; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_1000 = _GEN_2326 & _GEN_2271 ? Station3_4_4 : _GEN_999; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_1001 = _GEN_2326 & _GEN_2273 ? Station3_4_5 : _GEN_1000; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_1002 = _GEN_2326 & _GEN_2275 ? Station3_4_6 : _GEN_1001; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_1003 = _GEN_2326 & _GEN_2277 ? Station3_4_7 : _GEN_1002; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_1004 = _GEN_2342 & _GEN_2279 ? Station3_5_0 : _GEN_1003; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_1005 = _GEN_2342 & _GEN_2265 ? Station3_5_1 : _GEN_1004; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_1006 = _GEN_2342 & _GEN_2267 ? Station3_5_2 : _GEN_1005; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_1007 = _GEN_2342 & _GEN_2269 ? Station3_5_3 : _GEN_1006; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_1008 = _GEN_2342 & _GEN_2271 ? Station3_5_4 : _GEN_1007; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_1009 = _GEN_2342 & _GEN_2273 ? Station3_5_5 : _GEN_1008; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_1010 = _GEN_2342 & _GEN_2275 ? Station3_5_6 : _GEN_1009; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_1011 = _GEN_2342 & _GEN_2277 ? Station3_5_7 : _GEN_1010; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_1012 = _GEN_2358 & _GEN_2279 ? Station3_6_0 : _GEN_1011; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_1013 = _GEN_2358 & _GEN_2265 ? Station3_6_1 : _GEN_1012; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_1014 = _GEN_2358 & _GEN_2267 ? Station3_6_2 : _GEN_1013; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_1015 = _GEN_2358 & _GEN_2269 ? Station3_6_3 : _GEN_1014; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_1016 = _GEN_2358 & _GEN_2271 ? Station3_6_4 : _GEN_1015; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_1017 = _GEN_2358 & _GEN_2273 ? Station3_6_5 : _GEN_1016; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_1018 = _GEN_2358 & _GEN_2275 ? Station3_6_6 : _GEN_1017; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_1019 = _GEN_2358 & _GEN_2277 ? Station3_6_7 : _GEN_1018; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_1020 = _GEN_2374 & _GEN_2279 ? Station3_7_0 : _GEN_1019; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_1021 = _GEN_2374 & _GEN_2265 ? Station3_7_1 : _GEN_1020; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_1022 = _GEN_2374 & _GEN_2267 ? Station3_7_2 : _GEN_1021; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_1023 = _GEN_2374 & _GEN_2269 ? Station3_7_3 : _GEN_1022; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_1024 = _GEN_2374 & _GEN_2271 ? Station3_7_4 : _GEN_1023; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_1025 = _GEN_2374 & _GEN_2273 ? Station3_7_5 : _GEN_1024; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_1026 = _GEN_2374 & _GEN_2275 ? Station3_7_6 : _GEN_1025; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_1027 = _GEN_2374 & _GEN_2277 ? Station3_7_7 : _GEN_1026; // @[stationary_dpe.scala 127:{31,31}]
  wire [31:0] _GEN_1156 = _GEN_1027 != 16'h0 ? _count_T_1 : _GEN_963; // @[stationary_dpe.scala 127:39 130:18]
  wire [31:0] _GEN_1221 = ~valid2 ? _GEN_1156 : _GEN_963; // @[stationary_dpe.scala 126:29]
  wire  valid3 = count >= 32'h20; // @[stationary_dpe.scala 202:17]
  wire [15:0] _GEN_1223 = _GEN_2264 & _GEN_2265 ? Station4_0_1 : Station4_0_0; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1224 = _GEN_2264 & _GEN_2267 ? Station4_0_2 : _GEN_1223; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1225 = _GEN_2264 & _GEN_2269 ? Station4_0_3 : _GEN_1224; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1226 = _GEN_2264 & _GEN_2271 ? Station4_0_4 : _GEN_1225; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1227 = _GEN_2264 & _GEN_2273 ? Station4_0_5 : _GEN_1226; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1228 = _GEN_2264 & _GEN_2275 ? Station4_0_6 : _GEN_1227; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1229 = _GEN_2264 & _GEN_2277 ? Station4_0_7 : _GEN_1228; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1230 = _GEN_2278 & _GEN_2279 ? Station4_1_0 : _GEN_1229; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1231 = _GEN_2278 & _GEN_2265 ? Station4_1_1 : _GEN_1230; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1232 = _GEN_2278 & _GEN_2267 ? Station4_1_2 : _GEN_1231; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1233 = _GEN_2278 & _GEN_2269 ? Station4_1_3 : _GEN_1232; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1234 = _GEN_2278 & _GEN_2271 ? Station4_1_4 : _GEN_1233; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1235 = _GEN_2278 & _GEN_2273 ? Station4_1_5 : _GEN_1234; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1236 = _GEN_2278 & _GEN_2275 ? Station4_1_6 : _GEN_1235; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1237 = _GEN_2278 & _GEN_2277 ? Station4_1_7 : _GEN_1236; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1238 = _GEN_2294 & _GEN_2279 ? Station4_2_0 : _GEN_1237; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1239 = _GEN_2294 & _GEN_2265 ? Station4_2_1 : _GEN_1238; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1240 = _GEN_2294 & _GEN_2267 ? Station4_2_2 : _GEN_1239; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1241 = _GEN_2294 & _GEN_2269 ? Station4_2_3 : _GEN_1240; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1242 = _GEN_2294 & _GEN_2271 ? Station4_2_4 : _GEN_1241; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1243 = _GEN_2294 & _GEN_2273 ? Station4_2_5 : _GEN_1242; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1244 = _GEN_2294 & _GEN_2275 ? Station4_2_6 : _GEN_1243; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1245 = _GEN_2294 & _GEN_2277 ? Station4_2_7 : _GEN_1244; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1246 = _GEN_2310 & _GEN_2279 ? Station4_3_0 : _GEN_1245; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1247 = _GEN_2310 & _GEN_2265 ? Station4_3_1 : _GEN_1246; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1248 = _GEN_2310 & _GEN_2267 ? Station4_3_2 : _GEN_1247; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1249 = _GEN_2310 & _GEN_2269 ? Station4_3_3 : _GEN_1248; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1250 = _GEN_2310 & _GEN_2271 ? Station4_3_4 : _GEN_1249; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1251 = _GEN_2310 & _GEN_2273 ? Station4_3_5 : _GEN_1250; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1252 = _GEN_2310 & _GEN_2275 ? Station4_3_6 : _GEN_1251; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1253 = _GEN_2310 & _GEN_2277 ? Station4_3_7 : _GEN_1252; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1254 = _GEN_2326 & _GEN_2279 ? Station4_4_0 : _GEN_1253; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1255 = _GEN_2326 & _GEN_2265 ? Station4_4_1 : _GEN_1254; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1256 = _GEN_2326 & _GEN_2267 ? Station4_4_2 : _GEN_1255; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1257 = _GEN_2326 & _GEN_2269 ? Station4_4_3 : _GEN_1256; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1258 = _GEN_2326 & _GEN_2271 ? Station4_4_4 : _GEN_1257; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1259 = _GEN_2326 & _GEN_2273 ? Station4_4_5 : _GEN_1258; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1260 = _GEN_2326 & _GEN_2275 ? Station4_4_6 : _GEN_1259; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1261 = _GEN_2326 & _GEN_2277 ? Station4_4_7 : _GEN_1260; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1262 = _GEN_2342 & _GEN_2279 ? Station4_5_0 : _GEN_1261; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1263 = _GEN_2342 & _GEN_2265 ? Station4_5_1 : _GEN_1262; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1264 = _GEN_2342 & _GEN_2267 ? Station4_5_2 : _GEN_1263; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1265 = _GEN_2342 & _GEN_2269 ? Station4_5_3 : _GEN_1264; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1266 = _GEN_2342 & _GEN_2271 ? Station4_5_4 : _GEN_1265; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1267 = _GEN_2342 & _GEN_2273 ? Station4_5_5 : _GEN_1266; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1268 = _GEN_2342 & _GEN_2275 ? Station4_5_6 : _GEN_1267; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1269 = _GEN_2342 & _GEN_2277 ? Station4_5_7 : _GEN_1268; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1270 = _GEN_2358 & _GEN_2279 ? Station4_6_0 : _GEN_1269; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1271 = _GEN_2358 & _GEN_2265 ? Station4_6_1 : _GEN_1270; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1272 = _GEN_2358 & _GEN_2267 ? Station4_6_2 : _GEN_1271; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1273 = _GEN_2358 & _GEN_2269 ? Station4_6_3 : _GEN_1272; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1274 = _GEN_2358 & _GEN_2271 ? Station4_6_4 : _GEN_1273; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1275 = _GEN_2358 & _GEN_2273 ? Station4_6_5 : _GEN_1274; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1276 = _GEN_2358 & _GEN_2275 ? Station4_6_6 : _GEN_1275; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1277 = _GEN_2358 & _GEN_2277 ? Station4_6_7 : _GEN_1276; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1278 = _GEN_2374 & _GEN_2279 ? Station4_7_0 : _GEN_1277; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1279 = _GEN_2374 & _GEN_2265 ? Station4_7_1 : _GEN_1278; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1280 = _GEN_2374 & _GEN_2267 ? Station4_7_2 : _GEN_1279; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1281 = _GEN_2374 & _GEN_2269 ? Station4_7_3 : _GEN_1280; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1282 = _GEN_2374 & _GEN_2271 ? Station4_7_4 : _GEN_1281; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1283 = _GEN_2374 & _GEN_2273 ? Station4_7_5 : _GEN_1282; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1284 = _GEN_2374 & _GEN_2275 ? Station4_7_6 : _GEN_1283; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1285 = _GEN_2374 & _GEN_2277 ? Station4_7_7 : _GEN_1284; // @[stationary_dpe.scala 139:{31,31}]
  wire [31:0] _GEN_1414 = _GEN_1285 != 16'h0 ? _count_T_1 : _GEN_1221; // @[stationary_dpe.scala 139:39 142:18]
  wire [31:0] _GEN_1479 = ~valid3 ? _GEN_1414 : _GEN_1221; // @[stationary_dpe.scala 138:28]
  wire  valid4 = count >= 32'h28; // @[stationary_dpe.scala 206:17]
  wire [15:0] _GEN_1481 = _GEN_2264 & _GEN_2265 ? Station5_0_1 : Station5_0_0; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1482 = _GEN_2264 & _GEN_2267 ? Station5_0_2 : _GEN_1481; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1483 = _GEN_2264 & _GEN_2269 ? Station5_0_3 : _GEN_1482; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1484 = _GEN_2264 & _GEN_2271 ? Station5_0_4 : _GEN_1483; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1485 = _GEN_2264 & _GEN_2273 ? Station5_0_5 : _GEN_1484; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1486 = _GEN_2264 & _GEN_2275 ? Station5_0_6 : _GEN_1485; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1487 = _GEN_2264 & _GEN_2277 ? Station5_0_7 : _GEN_1486; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1488 = _GEN_2278 & _GEN_2279 ? Station5_1_0 : _GEN_1487; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1489 = _GEN_2278 & _GEN_2265 ? Station5_1_1 : _GEN_1488; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1490 = _GEN_2278 & _GEN_2267 ? Station5_1_2 : _GEN_1489; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1491 = _GEN_2278 & _GEN_2269 ? Station5_1_3 : _GEN_1490; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1492 = _GEN_2278 & _GEN_2271 ? Station5_1_4 : _GEN_1491; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1493 = _GEN_2278 & _GEN_2273 ? Station5_1_5 : _GEN_1492; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1494 = _GEN_2278 & _GEN_2275 ? Station5_1_6 : _GEN_1493; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1495 = _GEN_2278 & _GEN_2277 ? Station5_1_7 : _GEN_1494; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1496 = _GEN_2294 & _GEN_2279 ? Station5_2_0 : _GEN_1495; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1497 = _GEN_2294 & _GEN_2265 ? Station5_2_1 : _GEN_1496; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1498 = _GEN_2294 & _GEN_2267 ? Station5_2_2 : _GEN_1497; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1499 = _GEN_2294 & _GEN_2269 ? Station5_2_3 : _GEN_1498; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1500 = _GEN_2294 & _GEN_2271 ? Station5_2_4 : _GEN_1499; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1501 = _GEN_2294 & _GEN_2273 ? Station5_2_5 : _GEN_1500; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1502 = _GEN_2294 & _GEN_2275 ? Station5_2_6 : _GEN_1501; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1503 = _GEN_2294 & _GEN_2277 ? Station5_2_7 : _GEN_1502; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1504 = _GEN_2310 & _GEN_2279 ? Station5_3_0 : _GEN_1503; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1505 = _GEN_2310 & _GEN_2265 ? Station5_3_1 : _GEN_1504; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1506 = _GEN_2310 & _GEN_2267 ? Station5_3_2 : _GEN_1505; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1507 = _GEN_2310 & _GEN_2269 ? Station5_3_3 : _GEN_1506; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1508 = _GEN_2310 & _GEN_2271 ? Station5_3_4 : _GEN_1507; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1509 = _GEN_2310 & _GEN_2273 ? Station5_3_5 : _GEN_1508; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1510 = _GEN_2310 & _GEN_2275 ? Station5_3_6 : _GEN_1509; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1511 = _GEN_2310 & _GEN_2277 ? Station5_3_7 : _GEN_1510; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1512 = _GEN_2326 & _GEN_2279 ? Station5_4_0 : _GEN_1511; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1513 = _GEN_2326 & _GEN_2265 ? Station5_4_1 : _GEN_1512; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1514 = _GEN_2326 & _GEN_2267 ? Station5_4_2 : _GEN_1513; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1515 = _GEN_2326 & _GEN_2269 ? Station5_4_3 : _GEN_1514; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1516 = _GEN_2326 & _GEN_2271 ? Station5_4_4 : _GEN_1515; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1517 = _GEN_2326 & _GEN_2273 ? Station5_4_5 : _GEN_1516; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1518 = _GEN_2326 & _GEN_2275 ? Station5_4_6 : _GEN_1517; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1519 = _GEN_2326 & _GEN_2277 ? Station5_4_7 : _GEN_1518; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1520 = _GEN_2342 & _GEN_2279 ? Station5_5_0 : _GEN_1519; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1521 = _GEN_2342 & _GEN_2265 ? Station5_5_1 : _GEN_1520; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1522 = _GEN_2342 & _GEN_2267 ? Station5_5_2 : _GEN_1521; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1523 = _GEN_2342 & _GEN_2269 ? Station5_5_3 : _GEN_1522; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1524 = _GEN_2342 & _GEN_2271 ? Station5_5_4 : _GEN_1523; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1525 = _GEN_2342 & _GEN_2273 ? Station5_5_5 : _GEN_1524; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1526 = _GEN_2342 & _GEN_2275 ? Station5_5_6 : _GEN_1525; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1527 = _GEN_2342 & _GEN_2277 ? Station5_5_7 : _GEN_1526; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1528 = _GEN_2358 & _GEN_2279 ? Station5_6_0 : _GEN_1527; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1529 = _GEN_2358 & _GEN_2265 ? Station5_6_1 : _GEN_1528; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1530 = _GEN_2358 & _GEN_2267 ? Station5_6_2 : _GEN_1529; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1531 = _GEN_2358 & _GEN_2269 ? Station5_6_3 : _GEN_1530; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1532 = _GEN_2358 & _GEN_2271 ? Station5_6_4 : _GEN_1531; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1533 = _GEN_2358 & _GEN_2273 ? Station5_6_5 : _GEN_1532; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1534 = _GEN_2358 & _GEN_2275 ? Station5_6_6 : _GEN_1533; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1535 = _GEN_2358 & _GEN_2277 ? Station5_6_7 : _GEN_1534; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1536 = _GEN_2374 & _GEN_2279 ? Station5_7_0 : _GEN_1535; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1537 = _GEN_2374 & _GEN_2265 ? Station5_7_1 : _GEN_1536; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1538 = _GEN_2374 & _GEN_2267 ? Station5_7_2 : _GEN_1537; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1539 = _GEN_2374 & _GEN_2269 ? Station5_7_3 : _GEN_1538; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1540 = _GEN_2374 & _GEN_2271 ? Station5_7_4 : _GEN_1539; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1541 = _GEN_2374 & _GEN_2273 ? Station5_7_5 : _GEN_1540; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1542 = _GEN_2374 & _GEN_2275 ? Station5_7_6 : _GEN_1541; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1543 = _GEN_2374 & _GEN_2277 ? Station5_7_7 : _GEN_1542; // @[stationary_dpe.scala 151:{31,31}]
  wire [31:0] _GEN_1672 = _GEN_1543 != 16'h0 ? _count_T_1 : _GEN_1479; // @[stationary_dpe.scala 151:39 154:18]
  wire [31:0] _GEN_1737 = ~valid4 ? _GEN_1672 : _GEN_1479; // @[stationary_dpe.scala 150:28]
  wire  valid5 = count >= 32'h30; // @[stationary_dpe.scala 210:17]
  wire [15:0] _GEN_1739 = _GEN_2264 & _GEN_2265 ? Station6_0_1 : Station6_0_0; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1740 = _GEN_2264 & _GEN_2267 ? Station6_0_2 : _GEN_1739; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1741 = _GEN_2264 & _GEN_2269 ? Station6_0_3 : _GEN_1740; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1742 = _GEN_2264 & _GEN_2271 ? Station6_0_4 : _GEN_1741; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1743 = _GEN_2264 & _GEN_2273 ? Station6_0_5 : _GEN_1742; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1744 = _GEN_2264 & _GEN_2275 ? Station6_0_6 : _GEN_1743; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1745 = _GEN_2264 & _GEN_2277 ? Station6_0_7 : _GEN_1744; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1746 = _GEN_2278 & _GEN_2279 ? Station6_1_0 : _GEN_1745; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1747 = _GEN_2278 & _GEN_2265 ? Station6_1_1 : _GEN_1746; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1748 = _GEN_2278 & _GEN_2267 ? Station6_1_2 : _GEN_1747; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1749 = _GEN_2278 & _GEN_2269 ? Station6_1_3 : _GEN_1748; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1750 = _GEN_2278 & _GEN_2271 ? Station6_1_4 : _GEN_1749; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1751 = _GEN_2278 & _GEN_2273 ? Station6_1_5 : _GEN_1750; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1752 = _GEN_2278 & _GEN_2275 ? Station6_1_6 : _GEN_1751; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1753 = _GEN_2278 & _GEN_2277 ? Station6_1_7 : _GEN_1752; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1754 = _GEN_2294 & _GEN_2279 ? Station6_2_0 : _GEN_1753; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1755 = _GEN_2294 & _GEN_2265 ? Station6_2_1 : _GEN_1754; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1756 = _GEN_2294 & _GEN_2267 ? Station6_2_2 : _GEN_1755; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1757 = _GEN_2294 & _GEN_2269 ? Station6_2_3 : _GEN_1756; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1758 = _GEN_2294 & _GEN_2271 ? Station6_2_4 : _GEN_1757; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1759 = _GEN_2294 & _GEN_2273 ? Station6_2_5 : _GEN_1758; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1760 = _GEN_2294 & _GEN_2275 ? Station6_2_6 : _GEN_1759; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1761 = _GEN_2294 & _GEN_2277 ? Station6_2_7 : _GEN_1760; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1762 = _GEN_2310 & _GEN_2279 ? Station6_3_0 : _GEN_1761; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1763 = _GEN_2310 & _GEN_2265 ? Station6_3_1 : _GEN_1762; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1764 = _GEN_2310 & _GEN_2267 ? Station6_3_2 : _GEN_1763; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1765 = _GEN_2310 & _GEN_2269 ? Station6_3_3 : _GEN_1764; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1766 = _GEN_2310 & _GEN_2271 ? Station6_3_4 : _GEN_1765; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1767 = _GEN_2310 & _GEN_2273 ? Station6_3_5 : _GEN_1766; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1768 = _GEN_2310 & _GEN_2275 ? Station6_3_6 : _GEN_1767; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1769 = _GEN_2310 & _GEN_2277 ? Station6_3_7 : _GEN_1768; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1770 = _GEN_2326 & _GEN_2279 ? Station6_4_0 : _GEN_1769; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1771 = _GEN_2326 & _GEN_2265 ? Station6_4_1 : _GEN_1770; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1772 = _GEN_2326 & _GEN_2267 ? Station6_4_2 : _GEN_1771; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1773 = _GEN_2326 & _GEN_2269 ? Station6_4_3 : _GEN_1772; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1774 = _GEN_2326 & _GEN_2271 ? Station6_4_4 : _GEN_1773; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1775 = _GEN_2326 & _GEN_2273 ? Station6_4_5 : _GEN_1774; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1776 = _GEN_2326 & _GEN_2275 ? Station6_4_6 : _GEN_1775; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1777 = _GEN_2326 & _GEN_2277 ? Station6_4_7 : _GEN_1776; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1778 = _GEN_2342 & _GEN_2279 ? Station6_5_0 : _GEN_1777; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1779 = _GEN_2342 & _GEN_2265 ? Station6_5_1 : _GEN_1778; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1780 = _GEN_2342 & _GEN_2267 ? Station6_5_2 : _GEN_1779; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1781 = _GEN_2342 & _GEN_2269 ? Station6_5_3 : _GEN_1780; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1782 = _GEN_2342 & _GEN_2271 ? Station6_5_4 : _GEN_1781; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1783 = _GEN_2342 & _GEN_2273 ? Station6_5_5 : _GEN_1782; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1784 = _GEN_2342 & _GEN_2275 ? Station6_5_6 : _GEN_1783; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1785 = _GEN_2342 & _GEN_2277 ? Station6_5_7 : _GEN_1784; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1786 = _GEN_2358 & _GEN_2279 ? Station6_6_0 : _GEN_1785; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1787 = _GEN_2358 & _GEN_2265 ? Station6_6_1 : _GEN_1786; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1788 = _GEN_2358 & _GEN_2267 ? Station6_6_2 : _GEN_1787; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1789 = _GEN_2358 & _GEN_2269 ? Station6_6_3 : _GEN_1788; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1790 = _GEN_2358 & _GEN_2271 ? Station6_6_4 : _GEN_1789; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1791 = _GEN_2358 & _GEN_2273 ? Station6_6_5 : _GEN_1790; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1792 = _GEN_2358 & _GEN_2275 ? Station6_6_6 : _GEN_1791; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1793 = _GEN_2358 & _GEN_2277 ? Station6_6_7 : _GEN_1792; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1794 = _GEN_2374 & _GEN_2279 ? Station6_7_0 : _GEN_1793; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1795 = _GEN_2374 & _GEN_2265 ? Station6_7_1 : _GEN_1794; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1796 = _GEN_2374 & _GEN_2267 ? Station6_7_2 : _GEN_1795; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1797 = _GEN_2374 & _GEN_2269 ? Station6_7_3 : _GEN_1796; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1798 = _GEN_2374 & _GEN_2271 ? Station6_7_4 : _GEN_1797; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1799 = _GEN_2374 & _GEN_2273 ? Station6_7_5 : _GEN_1798; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1800 = _GEN_2374 & _GEN_2275 ? Station6_7_6 : _GEN_1799; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1801 = _GEN_2374 & _GEN_2277 ? Station6_7_7 : _GEN_1800; // @[stationary_dpe.scala 163:{31,31}]
  wire [31:0] _GEN_1930 = _GEN_1801 != 16'h0 ? _count_T_1 : _GEN_1737; // @[stationary_dpe.scala 163:39 166:18]
  wire [31:0] _GEN_1995 = ~valid5 ? _GEN_1930 : _GEN_1737; // @[stationary_dpe.scala 162:28]
  wire  valid6 = count >= 32'h38; // @[stationary_dpe.scala 215:17]
  wire [15:0] _GEN_1997 = _GEN_2264 & _GEN_2265 ? Station7_0_1 : Station7_0_0; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_1998 = _GEN_2264 & _GEN_2267 ? Station7_0_2 : _GEN_1997; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_1999 = _GEN_2264 & _GEN_2269 ? Station7_0_3 : _GEN_1998; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2000 = _GEN_2264 & _GEN_2271 ? Station7_0_4 : _GEN_1999; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2001 = _GEN_2264 & _GEN_2273 ? Station7_0_5 : _GEN_2000; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2002 = _GEN_2264 & _GEN_2275 ? Station7_0_6 : _GEN_2001; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2003 = _GEN_2264 & _GEN_2277 ? Station7_0_7 : _GEN_2002; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2004 = _GEN_2278 & _GEN_2279 ? Station7_1_0 : _GEN_2003; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2005 = _GEN_2278 & _GEN_2265 ? Station7_1_1 : _GEN_2004; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2006 = _GEN_2278 & _GEN_2267 ? Station7_1_2 : _GEN_2005; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2007 = _GEN_2278 & _GEN_2269 ? Station7_1_3 : _GEN_2006; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2008 = _GEN_2278 & _GEN_2271 ? Station7_1_4 : _GEN_2007; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2009 = _GEN_2278 & _GEN_2273 ? Station7_1_5 : _GEN_2008; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2010 = _GEN_2278 & _GEN_2275 ? Station7_1_6 : _GEN_2009; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2011 = _GEN_2278 & _GEN_2277 ? Station7_1_7 : _GEN_2010; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2012 = _GEN_2294 & _GEN_2279 ? Station7_2_0 : _GEN_2011; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2013 = _GEN_2294 & _GEN_2265 ? Station7_2_1 : _GEN_2012; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2014 = _GEN_2294 & _GEN_2267 ? Station7_2_2 : _GEN_2013; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2015 = _GEN_2294 & _GEN_2269 ? Station7_2_3 : _GEN_2014; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2016 = _GEN_2294 & _GEN_2271 ? Station7_2_4 : _GEN_2015; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2017 = _GEN_2294 & _GEN_2273 ? Station7_2_5 : _GEN_2016; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2018 = _GEN_2294 & _GEN_2275 ? Station7_2_6 : _GEN_2017; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2019 = _GEN_2294 & _GEN_2277 ? Station7_2_7 : _GEN_2018; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2020 = _GEN_2310 & _GEN_2279 ? Station7_3_0 : _GEN_2019; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2021 = _GEN_2310 & _GEN_2265 ? Station7_3_1 : _GEN_2020; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2022 = _GEN_2310 & _GEN_2267 ? Station7_3_2 : _GEN_2021; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2023 = _GEN_2310 & _GEN_2269 ? Station7_3_3 : _GEN_2022; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2024 = _GEN_2310 & _GEN_2271 ? Station7_3_4 : _GEN_2023; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2025 = _GEN_2310 & _GEN_2273 ? Station7_3_5 : _GEN_2024; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2026 = _GEN_2310 & _GEN_2275 ? Station7_3_6 : _GEN_2025; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2027 = _GEN_2310 & _GEN_2277 ? Station7_3_7 : _GEN_2026; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2028 = _GEN_2326 & _GEN_2279 ? Station7_4_0 : _GEN_2027; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2029 = _GEN_2326 & _GEN_2265 ? Station7_4_1 : _GEN_2028; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2030 = _GEN_2326 & _GEN_2267 ? Station7_4_2 : _GEN_2029; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2031 = _GEN_2326 & _GEN_2269 ? Station7_4_3 : _GEN_2030; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2032 = _GEN_2326 & _GEN_2271 ? Station7_4_4 : _GEN_2031; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2033 = _GEN_2326 & _GEN_2273 ? Station7_4_5 : _GEN_2032; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2034 = _GEN_2326 & _GEN_2275 ? Station7_4_6 : _GEN_2033; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2035 = _GEN_2326 & _GEN_2277 ? Station7_4_7 : _GEN_2034; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2036 = _GEN_2342 & _GEN_2279 ? Station7_5_0 : _GEN_2035; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2037 = _GEN_2342 & _GEN_2265 ? Station7_5_1 : _GEN_2036; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2038 = _GEN_2342 & _GEN_2267 ? Station7_5_2 : _GEN_2037; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2039 = _GEN_2342 & _GEN_2269 ? Station7_5_3 : _GEN_2038; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2040 = _GEN_2342 & _GEN_2271 ? Station7_5_4 : _GEN_2039; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2041 = _GEN_2342 & _GEN_2273 ? Station7_5_5 : _GEN_2040; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2042 = _GEN_2342 & _GEN_2275 ? Station7_5_6 : _GEN_2041; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2043 = _GEN_2342 & _GEN_2277 ? Station7_5_7 : _GEN_2042; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2044 = _GEN_2358 & _GEN_2279 ? Station7_6_0 : _GEN_2043; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2045 = _GEN_2358 & _GEN_2265 ? Station7_6_1 : _GEN_2044; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2046 = _GEN_2358 & _GEN_2267 ? Station7_6_2 : _GEN_2045; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2047 = _GEN_2358 & _GEN_2269 ? Station7_6_3 : _GEN_2046; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2048 = _GEN_2358 & _GEN_2271 ? Station7_6_4 : _GEN_2047; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2049 = _GEN_2358 & _GEN_2273 ? Station7_6_5 : _GEN_2048; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2050 = _GEN_2358 & _GEN_2275 ? Station7_6_6 : _GEN_2049; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2051 = _GEN_2358 & _GEN_2277 ? Station7_6_7 : _GEN_2050; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2052 = _GEN_2374 & _GEN_2279 ? Station7_7_0 : _GEN_2051; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2053 = _GEN_2374 & _GEN_2265 ? Station7_7_1 : _GEN_2052; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2054 = _GEN_2374 & _GEN_2267 ? Station7_7_2 : _GEN_2053; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2055 = _GEN_2374 & _GEN_2269 ? Station7_7_3 : _GEN_2054; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2056 = _GEN_2374 & _GEN_2271 ? Station7_7_4 : _GEN_2055; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2057 = _GEN_2374 & _GEN_2273 ? Station7_7_5 : _GEN_2056; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2058 = _GEN_2374 & _GEN_2275 ? Station7_7_6 : _GEN_2057; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2059 = _GEN_2374 & _GEN_2277 ? Station7_7_7 : _GEN_2058; // @[stationary_dpe.scala 175:{31,31}]
  wire  _T_57 = j == 32'h7; // @[stationary_dpe.scala 222:46]
  wire [31:0] _i_T_1 = i + 32'h1; // @[stationary_dpe.scala 223:16]
  wire [31:0] _j_T_1 = j + 32'h1; // @[stationary_dpe.scala 227:16]
  assign io_o_Stationary_matrix1_0_0 = io_Stationary_matrix_0_0; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_0_1 = io_Stationary_matrix_0_1; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_0_2 = io_Stationary_matrix_0_2; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_0_3 = io_Stationary_matrix_0_3; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_0_4 = io_Stationary_matrix_0_4; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_0_5 = io_Stationary_matrix_0_5; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_0_6 = io_Stationary_matrix_0_6; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_0_7 = io_Stationary_matrix_0_7; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_1_0 = io_Stationary_matrix_1_0; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_1_1 = io_Stationary_matrix_1_1; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_1_2 = io_Stationary_matrix_1_2; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_1_3 = io_Stationary_matrix_1_3; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_1_4 = io_Stationary_matrix_1_4; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_1_5 = io_Stationary_matrix_1_5; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_1_6 = io_Stationary_matrix_1_6; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_1_7 = io_Stationary_matrix_1_7; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_2_0 = io_Stationary_matrix_2_0; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_2_1 = io_Stationary_matrix_2_1; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_2_2 = io_Stationary_matrix_2_2; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_2_3 = io_Stationary_matrix_2_3; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_2_4 = io_Stationary_matrix_2_4; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_2_5 = io_Stationary_matrix_2_5; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_2_6 = io_Stationary_matrix_2_6; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_2_7 = io_Stationary_matrix_2_7; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_3_0 = io_Stationary_matrix_3_0; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_3_1 = io_Stationary_matrix_3_1; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_3_2 = io_Stationary_matrix_3_2; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_3_3 = io_Stationary_matrix_3_3; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_3_4 = io_Stationary_matrix_3_4; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_3_5 = io_Stationary_matrix_3_5; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_3_6 = io_Stationary_matrix_3_6; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_3_7 = io_Stationary_matrix_3_7; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_4_0 = io_Stationary_matrix_4_0; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_4_1 = io_Stationary_matrix_4_1; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_4_2 = io_Stationary_matrix_4_2; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_4_3 = io_Stationary_matrix_4_3; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_4_4 = io_Stationary_matrix_4_4; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_4_5 = io_Stationary_matrix_4_5; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_4_6 = io_Stationary_matrix_4_6; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_4_7 = io_Stationary_matrix_4_7; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_5_0 = io_Stationary_matrix_5_0; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_5_1 = io_Stationary_matrix_5_1; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_5_2 = io_Stationary_matrix_5_2; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_5_3 = io_Stationary_matrix_5_3; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_5_4 = io_Stationary_matrix_5_4; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_5_5 = io_Stationary_matrix_5_5; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_5_6 = io_Stationary_matrix_5_6; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_5_7 = io_Stationary_matrix_5_7; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_6_0 = io_Stationary_matrix_6_0; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_6_1 = io_Stationary_matrix_6_1; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_6_2 = io_Stationary_matrix_6_2; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_6_3 = io_Stationary_matrix_6_3; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_6_4 = io_Stationary_matrix_6_4; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_6_5 = io_Stationary_matrix_6_5; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_6_6 = io_Stationary_matrix_6_6; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_6_7 = io_Stationary_matrix_6_7; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_7_0 = io_Stationary_matrix_7_0; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_7_1 = io_Stationary_matrix_7_1; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_7_2 = io_Stationary_matrix_7_2; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_7_3 = io_Stationary_matrix_7_3; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_7_4 = io_Stationary_matrix_7_4; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_7_5 = io_Stationary_matrix_7_5; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_7_6 = io_Stationary_matrix_7_6; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_7_7 = io_Stationary_matrix_7_7; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix2_0_0 = Station2_0_0; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_0_1 = Station2_0_1; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_0_2 = Station2_0_2; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_0_3 = Station2_0_3; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_0_4 = Station2_0_4; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_0_5 = Station2_0_5; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_0_6 = Station2_0_6; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_0_7 = Station2_0_7; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_1_0 = Station2_1_0; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_1_1 = Station2_1_1; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_1_2 = Station2_1_2; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_1_3 = Station2_1_3; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_1_4 = Station2_1_4; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_1_5 = Station2_1_5; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_1_6 = Station2_1_6; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_1_7 = Station2_1_7; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_2_0 = Station2_2_0; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_2_1 = Station2_2_1; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_2_2 = Station2_2_2; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_2_3 = Station2_2_3; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_2_4 = Station2_2_4; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_2_5 = Station2_2_5; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_2_6 = Station2_2_6; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_2_7 = Station2_2_7; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_3_0 = Station2_3_0; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_3_1 = Station2_3_1; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_3_2 = Station2_3_2; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_3_3 = Station2_3_3; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_3_4 = Station2_3_4; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_3_5 = Station2_3_5; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_3_6 = Station2_3_6; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_3_7 = Station2_3_7; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_4_0 = Station2_4_0; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_4_1 = Station2_4_1; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_4_2 = Station2_4_2; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_4_3 = Station2_4_3; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_4_4 = Station2_4_4; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_4_5 = Station2_4_5; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_4_6 = Station2_4_6; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_4_7 = Station2_4_7; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_5_0 = Station2_5_0; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_5_1 = Station2_5_1; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_5_2 = Station2_5_2; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_5_3 = Station2_5_3; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_5_4 = Station2_5_4; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_5_5 = Station2_5_5; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_5_6 = Station2_5_6; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_5_7 = Station2_5_7; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_6_0 = Station2_6_0; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_6_1 = Station2_6_1; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_6_2 = Station2_6_2; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_6_3 = Station2_6_3; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_6_4 = Station2_6_4; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_6_5 = Station2_6_5; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_6_6 = Station2_6_6; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_6_7 = Station2_6_7; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_7_0 = Station2_7_0; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_7_1 = Station2_7_1; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_7_2 = Station2_7_2; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_7_3 = Station2_7_3; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_7_4 = Station2_7_4; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_7_5 = Station2_7_5; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_7_6 = Station2_7_6; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_7_7 = Station2_7_7; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix3_0_0 = Station3_0_0; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_0_1 = Station3_0_1; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_0_2 = Station3_0_2; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_0_3 = Station3_0_3; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_0_4 = Station3_0_4; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_0_5 = Station3_0_5; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_0_6 = Station3_0_6; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_0_7 = Station3_0_7; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_1_0 = Station3_1_0; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_1_1 = Station3_1_1; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_1_2 = Station3_1_2; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_1_3 = Station3_1_3; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_1_4 = Station3_1_4; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_1_5 = Station3_1_5; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_1_6 = Station3_1_6; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_1_7 = Station3_1_7; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_2_0 = Station3_2_0; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_2_1 = Station3_2_1; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_2_2 = Station3_2_2; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_2_3 = Station3_2_3; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_2_4 = Station3_2_4; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_2_5 = Station3_2_5; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_2_6 = Station3_2_6; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_2_7 = Station3_2_7; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_3_0 = Station3_3_0; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_3_1 = Station3_3_1; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_3_2 = Station3_3_2; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_3_3 = Station3_3_3; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_3_4 = Station3_3_4; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_3_5 = Station3_3_5; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_3_6 = Station3_3_6; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_3_7 = Station3_3_7; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_4_0 = Station3_4_0; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_4_1 = Station3_4_1; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_4_2 = Station3_4_2; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_4_3 = Station3_4_3; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_4_4 = Station3_4_4; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_4_5 = Station3_4_5; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_4_6 = Station3_4_6; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_4_7 = Station3_4_7; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_5_0 = Station3_5_0; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_5_1 = Station3_5_1; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_5_2 = Station3_5_2; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_5_3 = Station3_5_3; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_5_4 = Station3_5_4; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_5_5 = Station3_5_5; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_5_6 = Station3_5_6; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_5_7 = Station3_5_7; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_6_0 = Station3_6_0; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_6_1 = Station3_6_1; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_6_2 = Station3_6_2; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_6_3 = Station3_6_3; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_6_4 = Station3_6_4; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_6_5 = Station3_6_5; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_6_6 = Station3_6_6; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_6_7 = Station3_6_7; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_7_0 = Station3_7_0; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_7_1 = Station3_7_1; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_7_2 = Station3_7_2; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_7_3 = Station3_7_3; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_7_4 = Station3_7_4; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_7_5 = Station3_7_5; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_7_6 = Station3_7_6; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_7_7 = Station3_7_7; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix4_0_0 = Station4_0_0; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_0_1 = Station4_0_1; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_0_2 = Station4_0_2; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_0_3 = Station4_0_3; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_0_4 = Station4_0_4; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_0_5 = Station4_0_5; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_0_6 = Station4_0_6; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_0_7 = Station4_0_7; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_1_0 = Station4_1_0; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_1_1 = Station4_1_1; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_1_2 = Station4_1_2; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_1_3 = Station4_1_3; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_1_4 = Station4_1_4; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_1_5 = Station4_1_5; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_1_6 = Station4_1_6; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_1_7 = Station4_1_7; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_2_0 = Station4_2_0; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_2_1 = Station4_2_1; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_2_2 = Station4_2_2; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_2_3 = Station4_2_3; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_2_4 = Station4_2_4; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_2_5 = Station4_2_5; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_2_6 = Station4_2_6; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_2_7 = Station4_2_7; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_3_0 = Station4_3_0; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_3_1 = Station4_3_1; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_3_2 = Station4_3_2; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_3_3 = Station4_3_3; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_3_4 = Station4_3_4; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_3_5 = Station4_3_5; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_3_6 = Station4_3_6; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_3_7 = Station4_3_7; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_4_0 = Station4_4_0; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_4_1 = Station4_4_1; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_4_2 = Station4_4_2; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_4_3 = Station4_4_3; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_4_4 = Station4_4_4; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_4_5 = Station4_4_5; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_4_6 = Station4_4_6; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_4_7 = Station4_4_7; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_5_0 = Station4_5_0; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_5_1 = Station4_5_1; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_5_2 = Station4_5_2; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_5_3 = Station4_5_3; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_5_4 = Station4_5_4; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_5_5 = Station4_5_5; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_5_6 = Station4_5_6; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_5_7 = Station4_5_7; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_6_0 = Station4_6_0; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_6_1 = Station4_6_1; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_6_2 = Station4_6_2; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_6_3 = Station4_6_3; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_6_4 = Station4_6_4; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_6_5 = Station4_6_5; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_6_6 = Station4_6_6; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_6_7 = Station4_6_7; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_7_0 = Station4_7_0; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_7_1 = Station4_7_1; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_7_2 = Station4_7_2; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_7_3 = Station4_7_3; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_7_4 = Station4_7_4; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_7_5 = Station4_7_5; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_7_6 = Station4_7_6; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_7_7 = Station4_7_7; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix5_0_0 = Station5_0_0; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_0_1 = Station5_0_1; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_0_2 = Station5_0_2; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_0_3 = Station5_0_3; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_0_4 = Station5_0_4; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_0_5 = Station5_0_5; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_0_6 = Station5_0_6; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_0_7 = Station5_0_7; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_1_0 = Station5_1_0; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_1_1 = Station5_1_1; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_1_2 = Station5_1_2; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_1_3 = Station5_1_3; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_1_4 = Station5_1_4; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_1_5 = Station5_1_5; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_1_6 = Station5_1_6; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_1_7 = Station5_1_7; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_2_0 = Station5_2_0; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_2_1 = Station5_2_1; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_2_2 = Station5_2_2; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_2_3 = Station5_2_3; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_2_4 = Station5_2_4; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_2_5 = Station5_2_5; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_2_6 = Station5_2_6; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_2_7 = Station5_2_7; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_3_0 = Station5_3_0; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_3_1 = Station5_3_1; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_3_2 = Station5_3_2; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_3_3 = Station5_3_3; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_3_4 = Station5_3_4; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_3_5 = Station5_3_5; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_3_6 = Station5_3_6; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_3_7 = Station5_3_7; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_4_0 = Station5_4_0; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_4_1 = Station5_4_1; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_4_2 = Station5_4_2; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_4_3 = Station5_4_3; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_4_4 = Station5_4_4; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_4_5 = Station5_4_5; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_4_6 = Station5_4_6; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_4_7 = Station5_4_7; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_5_0 = Station5_5_0; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_5_1 = Station5_5_1; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_5_2 = Station5_5_2; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_5_3 = Station5_5_3; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_5_4 = Station5_5_4; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_5_5 = Station5_5_5; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_5_6 = Station5_5_6; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_5_7 = Station5_5_7; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_6_0 = Station5_6_0; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_6_1 = Station5_6_1; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_6_2 = Station5_6_2; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_6_3 = Station5_6_3; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_6_4 = Station5_6_4; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_6_5 = Station5_6_5; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_6_6 = Station5_6_6; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_6_7 = Station5_6_7; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_7_0 = Station5_7_0; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_7_1 = Station5_7_1; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_7_2 = Station5_7_2; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_7_3 = Station5_7_3; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_7_4 = Station5_7_4; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_7_5 = Station5_7_5; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_7_6 = Station5_7_6; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_7_7 = Station5_7_7; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix6_0_0 = Station6_0_0; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_0_1 = Station6_0_1; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_0_2 = Station6_0_2; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_0_3 = Station6_0_3; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_0_4 = Station6_0_4; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_0_5 = Station6_0_5; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_0_6 = Station6_0_6; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_0_7 = Station6_0_7; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_1_0 = Station6_1_0; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_1_1 = Station6_1_1; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_1_2 = Station6_1_2; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_1_3 = Station6_1_3; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_1_4 = Station6_1_4; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_1_5 = Station6_1_5; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_1_6 = Station6_1_6; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_1_7 = Station6_1_7; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_2_0 = Station6_2_0; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_2_1 = Station6_2_1; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_2_2 = Station6_2_2; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_2_3 = Station6_2_3; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_2_4 = Station6_2_4; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_2_5 = Station6_2_5; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_2_6 = Station6_2_6; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_2_7 = Station6_2_7; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_3_0 = Station6_3_0; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_3_1 = Station6_3_1; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_3_2 = Station6_3_2; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_3_3 = Station6_3_3; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_3_4 = Station6_3_4; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_3_5 = Station6_3_5; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_3_6 = Station6_3_6; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_3_7 = Station6_3_7; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_4_0 = Station6_4_0; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_4_1 = Station6_4_1; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_4_2 = Station6_4_2; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_4_3 = Station6_4_3; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_4_4 = Station6_4_4; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_4_5 = Station6_4_5; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_4_6 = Station6_4_6; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_4_7 = Station6_4_7; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_5_0 = Station6_5_0; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_5_1 = Station6_5_1; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_5_2 = Station6_5_2; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_5_3 = Station6_5_3; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_5_4 = Station6_5_4; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_5_5 = Station6_5_5; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_5_6 = Station6_5_6; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_5_7 = Station6_5_7; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_6_0 = Station6_6_0; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_6_1 = Station6_6_1; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_6_2 = Station6_6_2; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_6_3 = Station6_6_3; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_6_4 = Station6_6_4; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_6_5 = Station6_6_5; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_6_6 = Station6_6_6; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_6_7 = Station6_6_7; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_7_0 = Station6_7_0; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_7_1 = Station6_7_1; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_7_2 = Station6_7_2; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_7_3 = Station6_7_3; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_7_4 = Station6_7_4; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_7_5 = Station6_7_5; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_7_6 = Station6_7_6; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_7_7 = Station6_7_7; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix7_0_0 = Station7_0_0; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_0_1 = Station7_0_1; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_0_2 = Station7_0_2; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_0_3 = Station7_0_3; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_0_4 = Station7_0_4; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_0_5 = Station7_0_5; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_0_6 = Station7_0_6; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_0_7 = Station7_0_7; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_1_0 = Station7_1_0; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_1_1 = Station7_1_1; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_1_2 = Station7_1_2; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_1_3 = Station7_1_3; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_1_4 = Station7_1_4; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_1_5 = Station7_1_5; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_1_6 = Station7_1_6; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_1_7 = Station7_1_7; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_2_0 = Station7_2_0; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_2_1 = Station7_2_1; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_2_2 = Station7_2_2; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_2_3 = Station7_2_3; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_2_4 = Station7_2_4; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_2_5 = Station7_2_5; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_2_6 = Station7_2_6; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_2_7 = Station7_2_7; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_3_0 = Station7_3_0; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_3_1 = Station7_3_1; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_3_2 = Station7_3_2; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_3_3 = Station7_3_3; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_3_4 = Station7_3_4; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_3_5 = Station7_3_5; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_3_6 = Station7_3_6; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_3_7 = Station7_3_7; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_4_0 = Station7_4_0; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_4_1 = Station7_4_1; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_4_2 = Station7_4_2; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_4_3 = Station7_4_3; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_4_4 = Station7_4_4; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_4_5 = Station7_4_5; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_4_6 = Station7_4_6; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_4_7 = Station7_4_7; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_5_0 = Station7_5_0; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_5_1 = Station7_5_1; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_5_2 = Station7_5_2; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_5_3 = Station7_5_3; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_5_4 = Station7_5_4; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_5_5 = Station7_5_5; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_5_6 = Station7_5_6; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_5_7 = Station7_5_7; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_6_0 = Station7_6_0; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_6_1 = Station7_6_1; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_6_2 = Station7_6_2; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_6_3 = Station7_6_3; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_6_4 = Station7_6_4; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_6_5 = Station7_6_5; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_6_6 = Station7_6_6; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_6_7 = Station7_6_7; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_7_0 = Station7_7_0; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_7_1 = Station7_7_1; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_7_2 = Station7_7_2; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_7_3 = Station7_7_3; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_7_4 = Station7_7_4; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_7_5 = Station7_7_5; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_7_6 = Station7_7_6; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_7_7 = Station7_7_7; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix8_0_0 = Station8_0_0; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_0_1 = Station8_0_1; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_0_2 = Station8_0_2; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_0_3 = Station8_0_3; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_0_4 = Station8_0_4; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_0_5 = Station8_0_5; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_0_6 = Station8_0_6; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_0_7 = Station8_0_7; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_1_0 = Station8_1_0; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_1_1 = Station8_1_1; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_1_2 = Station8_1_2; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_1_3 = Station8_1_3; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_1_4 = Station8_1_4; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_1_5 = Station8_1_5; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_1_6 = Station8_1_6; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_1_7 = Station8_1_7; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_2_0 = Station8_2_0; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_2_1 = Station8_2_1; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_2_2 = Station8_2_2; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_2_3 = Station8_2_3; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_2_4 = Station8_2_4; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_2_5 = Station8_2_5; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_2_6 = Station8_2_6; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_2_7 = Station8_2_7; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_3_0 = Station8_3_0; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_3_1 = Station8_3_1; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_3_2 = Station8_3_2; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_3_3 = Station8_3_3; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_3_4 = Station8_3_4; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_3_5 = Station8_3_5; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_3_6 = Station8_3_6; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_3_7 = Station8_3_7; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_4_0 = Station8_4_0; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_4_1 = Station8_4_1; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_4_2 = Station8_4_2; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_4_3 = Station8_4_3; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_4_4 = Station8_4_4; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_4_5 = Station8_4_5; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_4_6 = Station8_4_6; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_4_7 = Station8_4_7; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_5_0 = Station8_5_0; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_5_1 = Station8_5_1; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_5_2 = Station8_5_2; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_5_3 = Station8_5_3; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_5_4 = Station8_5_4; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_5_5 = Station8_5_5; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_5_6 = Station8_5_6; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_5_7 = Station8_5_7; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_6_0 = Station8_6_0; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_6_1 = Station8_6_1; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_6_2 = Station8_6_2; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_6_3 = Station8_6_3; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_6_4 = Station8_6_4; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_6_5 = Station8_6_5; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_6_6 = Station8_6_6; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_6_7 = Station8_6_7; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_7_0 = Station8_7_0; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_7_1 = Station8_7_1; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_7_2 = Station8_7_2; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_7_3 = Station8_7_3; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_7_4 = Station8_7_4; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_7_5 = Station8_7_5; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_7_6 = Station8_7_6; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_7_7 = Station8_7_7; // @[stationary_dpe.scala 184:29]
  always @(posedge clock) begin
    if (reset) begin // @[stationary_dpe.scala 23:27]
      count <= 32'h0; // @[stationary_dpe.scala 23:27]
    end else if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        count <= _count_T_1; // @[stationary_dpe.scala 178:18]
      end else begin
        count <= _GEN_1995;
      end
    end else begin
      count <= _GEN_1995;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2264 & _GEN_2279) begin // @[stationary_dpe.scala 95:32]
          Station2_0_0 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_0_0 <= _GEN_0;
        end
      end else begin
        Station2_0_0 <= _GEN_0;
      end
    end else begin
      Station2_0_0 <= _GEN_0;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2264 & _GEN_2265) begin // @[stationary_dpe.scala 95:32]
          Station2_0_1 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_0_1 <= _GEN_1;
        end
      end else begin
        Station2_0_1 <= _GEN_1;
      end
    end else begin
      Station2_0_1 <= _GEN_1;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2264 & _GEN_2267) begin // @[stationary_dpe.scala 95:32]
          Station2_0_2 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_0_2 <= _GEN_2;
        end
      end else begin
        Station2_0_2 <= _GEN_2;
      end
    end else begin
      Station2_0_2 <= _GEN_2;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2264 & _GEN_2269) begin // @[stationary_dpe.scala 95:32]
          Station2_0_3 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_0_3 <= _GEN_3;
        end
      end else begin
        Station2_0_3 <= _GEN_3;
      end
    end else begin
      Station2_0_3 <= _GEN_3;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2264 & _GEN_2271) begin // @[stationary_dpe.scala 95:32]
          Station2_0_4 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_0_4 <= _GEN_4;
        end
      end else begin
        Station2_0_4 <= _GEN_4;
      end
    end else begin
      Station2_0_4 <= _GEN_4;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2264 & _GEN_2273) begin // @[stationary_dpe.scala 95:32]
          Station2_0_5 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_0_5 <= _GEN_5;
        end
      end else begin
        Station2_0_5 <= _GEN_5;
      end
    end else begin
      Station2_0_5 <= _GEN_5;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2264 & _GEN_2275) begin // @[stationary_dpe.scala 95:32]
          Station2_0_6 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_0_6 <= _GEN_6;
        end
      end else begin
        Station2_0_6 <= _GEN_6;
      end
    end else begin
      Station2_0_6 <= _GEN_6;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2264 & _GEN_2277) begin // @[stationary_dpe.scala 95:32]
          Station2_0_7 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_0_7 <= _GEN_7;
        end
      end else begin
        Station2_0_7 <= _GEN_7;
      end
    end else begin
      Station2_0_7 <= _GEN_7;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2278 & _GEN_2279) begin // @[stationary_dpe.scala 95:32]
          Station2_1_0 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_1_0 <= _GEN_8;
        end
      end else begin
        Station2_1_0 <= _GEN_8;
      end
    end else begin
      Station2_1_0 <= _GEN_8;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2278 & _GEN_2265) begin // @[stationary_dpe.scala 95:32]
          Station2_1_1 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_1_1 <= _GEN_9;
        end
      end else begin
        Station2_1_1 <= _GEN_9;
      end
    end else begin
      Station2_1_1 <= _GEN_9;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2278 & _GEN_2267) begin // @[stationary_dpe.scala 95:32]
          Station2_1_2 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_1_2 <= _GEN_10;
        end
      end else begin
        Station2_1_2 <= _GEN_10;
      end
    end else begin
      Station2_1_2 <= _GEN_10;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2278 & _GEN_2269) begin // @[stationary_dpe.scala 95:32]
          Station2_1_3 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_1_3 <= _GEN_11;
        end
      end else begin
        Station2_1_3 <= _GEN_11;
      end
    end else begin
      Station2_1_3 <= _GEN_11;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2278 & _GEN_2271) begin // @[stationary_dpe.scala 95:32]
          Station2_1_4 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_1_4 <= _GEN_12;
        end
      end else begin
        Station2_1_4 <= _GEN_12;
      end
    end else begin
      Station2_1_4 <= _GEN_12;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2278 & _GEN_2273) begin // @[stationary_dpe.scala 95:32]
          Station2_1_5 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_1_5 <= _GEN_13;
        end
      end else begin
        Station2_1_5 <= _GEN_13;
      end
    end else begin
      Station2_1_5 <= _GEN_13;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2278 & _GEN_2275) begin // @[stationary_dpe.scala 95:32]
          Station2_1_6 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_1_6 <= _GEN_14;
        end
      end else begin
        Station2_1_6 <= _GEN_14;
      end
    end else begin
      Station2_1_6 <= _GEN_14;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2278 & _GEN_2277) begin // @[stationary_dpe.scala 95:32]
          Station2_1_7 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_1_7 <= _GEN_15;
        end
      end else begin
        Station2_1_7 <= _GEN_15;
      end
    end else begin
      Station2_1_7 <= _GEN_15;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2294 & _GEN_2279) begin // @[stationary_dpe.scala 95:32]
          Station2_2_0 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_2_0 <= _GEN_16;
        end
      end else begin
        Station2_2_0 <= _GEN_16;
      end
    end else begin
      Station2_2_0 <= _GEN_16;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2294 & _GEN_2265) begin // @[stationary_dpe.scala 95:32]
          Station2_2_1 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_2_1 <= _GEN_17;
        end
      end else begin
        Station2_2_1 <= _GEN_17;
      end
    end else begin
      Station2_2_1 <= _GEN_17;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2294 & _GEN_2267) begin // @[stationary_dpe.scala 95:32]
          Station2_2_2 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_2_2 <= _GEN_18;
        end
      end else begin
        Station2_2_2 <= _GEN_18;
      end
    end else begin
      Station2_2_2 <= _GEN_18;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2294 & _GEN_2269) begin // @[stationary_dpe.scala 95:32]
          Station2_2_3 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_2_3 <= _GEN_19;
        end
      end else begin
        Station2_2_3 <= _GEN_19;
      end
    end else begin
      Station2_2_3 <= _GEN_19;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2294 & _GEN_2271) begin // @[stationary_dpe.scala 95:32]
          Station2_2_4 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_2_4 <= _GEN_20;
        end
      end else begin
        Station2_2_4 <= _GEN_20;
      end
    end else begin
      Station2_2_4 <= _GEN_20;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2294 & _GEN_2273) begin // @[stationary_dpe.scala 95:32]
          Station2_2_5 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_2_5 <= _GEN_21;
        end
      end else begin
        Station2_2_5 <= _GEN_21;
      end
    end else begin
      Station2_2_5 <= _GEN_21;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2294 & _GEN_2275) begin // @[stationary_dpe.scala 95:32]
          Station2_2_6 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_2_6 <= _GEN_22;
        end
      end else begin
        Station2_2_6 <= _GEN_22;
      end
    end else begin
      Station2_2_6 <= _GEN_22;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2294 & _GEN_2277) begin // @[stationary_dpe.scala 95:32]
          Station2_2_7 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_2_7 <= _GEN_23;
        end
      end else begin
        Station2_2_7 <= _GEN_23;
      end
    end else begin
      Station2_2_7 <= _GEN_23;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2310 & _GEN_2279) begin // @[stationary_dpe.scala 95:32]
          Station2_3_0 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_3_0 <= _GEN_24;
        end
      end else begin
        Station2_3_0 <= _GEN_24;
      end
    end else begin
      Station2_3_0 <= _GEN_24;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2310 & _GEN_2265) begin // @[stationary_dpe.scala 95:32]
          Station2_3_1 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_3_1 <= _GEN_25;
        end
      end else begin
        Station2_3_1 <= _GEN_25;
      end
    end else begin
      Station2_3_1 <= _GEN_25;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2310 & _GEN_2267) begin // @[stationary_dpe.scala 95:32]
          Station2_3_2 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_3_2 <= _GEN_26;
        end
      end else begin
        Station2_3_2 <= _GEN_26;
      end
    end else begin
      Station2_3_2 <= _GEN_26;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2310 & _GEN_2269) begin // @[stationary_dpe.scala 95:32]
          Station2_3_3 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_3_3 <= _GEN_27;
        end
      end else begin
        Station2_3_3 <= _GEN_27;
      end
    end else begin
      Station2_3_3 <= _GEN_27;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2310 & _GEN_2271) begin // @[stationary_dpe.scala 95:32]
          Station2_3_4 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_3_4 <= _GEN_28;
        end
      end else begin
        Station2_3_4 <= _GEN_28;
      end
    end else begin
      Station2_3_4 <= _GEN_28;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2310 & _GEN_2273) begin // @[stationary_dpe.scala 95:32]
          Station2_3_5 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_3_5 <= _GEN_29;
        end
      end else begin
        Station2_3_5 <= _GEN_29;
      end
    end else begin
      Station2_3_5 <= _GEN_29;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2310 & _GEN_2275) begin // @[stationary_dpe.scala 95:32]
          Station2_3_6 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_3_6 <= _GEN_30;
        end
      end else begin
        Station2_3_6 <= _GEN_30;
      end
    end else begin
      Station2_3_6 <= _GEN_30;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2310 & _GEN_2277) begin // @[stationary_dpe.scala 95:32]
          Station2_3_7 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_3_7 <= _GEN_31;
        end
      end else begin
        Station2_3_7 <= _GEN_31;
      end
    end else begin
      Station2_3_7 <= _GEN_31;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2326 & _GEN_2279) begin // @[stationary_dpe.scala 95:32]
          Station2_4_0 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_4_0 <= _GEN_32;
        end
      end else begin
        Station2_4_0 <= _GEN_32;
      end
    end else begin
      Station2_4_0 <= _GEN_32;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2326 & _GEN_2265) begin // @[stationary_dpe.scala 95:32]
          Station2_4_1 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_4_1 <= _GEN_33;
        end
      end else begin
        Station2_4_1 <= _GEN_33;
      end
    end else begin
      Station2_4_1 <= _GEN_33;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2326 & _GEN_2267) begin // @[stationary_dpe.scala 95:32]
          Station2_4_2 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_4_2 <= _GEN_34;
        end
      end else begin
        Station2_4_2 <= _GEN_34;
      end
    end else begin
      Station2_4_2 <= _GEN_34;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2326 & _GEN_2269) begin // @[stationary_dpe.scala 95:32]
          Station2_4_3 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_4_3 <= _GEN_35;
        end
      end else begin
        Station2_4_3 <= _GEN_35;
      end
    end else begin
      Station2_4_3 <= _GEN_35;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2326 & _GEN_2271) begin // @[stationary_dpe.scala 95:32]
          Station2_4_4 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_4_4 <= _GEN_36;
        end
      end else begin
        Station2_4_4 <= _GEN_36;
      end
    end else begin
      Station2_4_4 <= _GEN_36;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2326 & _GEN_2273) begin // @[stationary_dpe.scala 95:32]
          Station2_4_5 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_4_5 <= _GEN_37;
        end
      end else begin
        Station2_4_5 <= _GEN_37;
      end
    end else begin
      Station2_4_5 <= _GEN_37;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2326 & _GEN_2275) begin // @[stationary_dpe.scala 95:32]
          Station2_4_6 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_4_6 <= _GEN_38;
        end
      end else begin
        Station2_4_6 <= _GEN_38;
      end
    end else begin
      Station2_4_6 <= _GEN_38;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2326 & _GEN_2277) begin // @[stationary_dpe.scala 95:32]
          Station2_4_7 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_4_7 <= _GEN_39;
        end
      end else begin
        Station2_4_7 <= _GEN_39;
      end
    end else begin
      Station2_4_7 <= _GEN_39;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2342 & _GEN_2279) begin // @[stationary_dpe.scala 95:32]
          Station2_5_0 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_5_0 <= _GEN_40;
        end
      end else begin
        Station2_5_0 <= _GEN_40;
      end
    end else begin
      Station2_5_0 <= _GEN_40;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2342 & _GEN_2265) begin // @[stationary_dpe.scala 95:32]
          Station2_5_1 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_5_1 <= _GEN_41;
        end
      end else begin
        Station2_5_1 <= _GEN_41;
      end
    end else begin
      Station2_5_1 <= _GEN_41;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2342 & _GEN_2267) begin // @[stationary_dpe.scala 95:32]
          Station2_5_2 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_5_2 <= _GEN_42;
        end
      end else begin
        Station2_5_2 <= _GEN_42;
      end
    end else begin
      Station2_5_2 <= _GEN_42;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2342 & _GEN_2269) begin // @[stationary_dpe.scala 95:32]
          Station2_5_3 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_5_3 <= _GEN_43;
        end
      end else begin
        Station2_5_3 <= _GEN_43;
      end
    end else begin
      Station2_5_3 <= _GEN_43;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2342 & _GEN_2271) begin // @[stationary_dpe.scala 95:32]
          Station2_5_4 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_5_4 <= _GEN_44;
        end
      end else begin
        Station2_5_4 <= _GEN_44;
      end
    end else begin
      Station2_5_4 <= _GEN_44;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2342 & _GEN_2273) begin // @[stationary_dpe.scala 95:32]
          Station2_5_5 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_5_5 <= _GEN_45;
        end
      end else begin
        Station2_5_5 <= _GEN_45;
      end
    end else begin
      Station2_5_5 <= _GEN_45;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2342 & _GEN_2275) begin // @[stationary_dpe.scala 95:32]
          Station2_5_6 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_5_6 <= _GEN_46;
        end
      end else begin
        Station2_5_6 <= _GEN_46;
      end
    end else begin
      Station2_5_6 <= _GEN_46;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2342 & _GEN_2277) begin // @[stationary_dpe.scala 95:32]
          Station2_5_7 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_5_7 <= _GEN_47;
        end
      end else begin
        Station2_5_7 <= _GEN_47;
      end
    end else begin
      Station2_5_7 <= _GEN_47;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2358 & _GEN_2279) begin // @[stationary_dpe.scala 95:32]
          Station2_6_0 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_6_0 <= _GEN_48;
        end
      end else begin
        Station2_6_0 <= _GEN_48;
      end
    end else begin
      Station2_6_0 <= _GEN_48;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2358 & _GEN_2265) begin // @[stationary_dpe.scala 95:32]
          Station2_6_1 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_6_1 <= _GEN_49;
        end
      end else begin
        Station2_6_1 <= _GEN_49;
      end
    end else begin
      Station2_6_1 <= _GEN_49;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2358 & _GEN_2267) begin // @[stationary_dpe.scala 95:32]
          Station2_6_2 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_6_2 <= _GEN_50;
        end
      end else begin
        Station2_6_2 <= _GEN_50;
      end
    end else begin
      Station2_6_2 <= _GEN_50;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2358 & _GEN_2269) begin // @[stationary_dpe.scala 95:32]
          Station2_6_3 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_6_3 <= _GEN_51;
        end
      end else begin
        Station2_6_3 <= _GEN_51;
      end
    end else begin
      Station2_6_3 <= _GEN_51;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2358 & _GEN_2271) begin // @[stationary_dpe.scala 95:32]
          Station2_6_4 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_6_4 <= _GEN_52;
        end
      end else begin
        Station2_6_4 <= _GEN_52;
      end
    end else begin
      Station2_6_4 <= _GEN_52;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2358 & _GEN_2273) begin // @[stationary_dpe.scala 95:32]
          Station2_6_5 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_6_5 <= _GEN_53;
        end
      end else begin
        Station2_6_5 <= _GEN_53;
      end
    end else begin
      Station2_6_5 <= _GEN_53;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2358 & _GEN_2275) begin // @[stationary_dpe.scala 95:32]
          Station2_6_6 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_6_6 <= _GEN_54;
        end
      end else begin
        Station2_6_6 <= _GEN_54;
      end
    end else begin
      Station2_6_6 <= _GEN_54;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2358 & _GEN_2277) begin // @[stationary_dpe.scala 95:32]
          Station2_6_7 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_6_7 <= _GEN_55;
        end
      end else begin
        Station2_6_7 <= _GEN_55;
      end
    end else begin
      Station2_6_7 <= _GEN_55;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2374 & _GEN_2279) begin // @[stationary_dpe.scala 95:32]
          Station2_7_0 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_7_0 <= _GEN_56;
        end
      end else begin
        Station2_7_0 <= _GEN_56;
      end
    end else begin
      Station2_7_0 <= _GEN_56;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2374 & _GEN_2265) begin // @[stationary_dpe.scala 95:32]
          Station2_7_1 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_7_1 <= _GEN_57;
        end
      end else begin
        Station2_7_1 <= _GEN_57;
      end
    end else begin
      Station2_7_1 <= _GEN_57;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2374 & _GEN_2267) begin // @[stationary_dpe.scala 95:32]
          Station2_7_2 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_7_2 <= _GEN_58;
        end
      end else begin
        Station2_7_2 <= _GEN_58;
      end
    end else begin
      Station2_7_2 <= _GEN_58;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2374 & _GEN_2269) begin // @[stationary_dpe.scala 95:32]
          Station2_7_3 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_7_3 <= _GEN_59;
        end
      end else begin
        Station2_7_3 <= _GEN_59;
      end
    end else begin
      Station2_7_3 <= _GEN_59;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2374 & _GEN_2271) begin // @[stationary_dpe.scala 95:32]
          Station2_7_4 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_7_4 <= _GEN_60;
        end
      end else begin
        Station2_7_4 <= _GEN_60;
      end
    end else begin
      Station2_7_4 <= _GEN_60;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2374 & _GEN_2273) begin // @[stationary_dpe.scala 95:32]
          Station2_7_5 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_7_5 <= _GEN_61;
        end
      end else begin
        Station2_7_5 <= _GEN_61;
      end
    end else begin
      Station2_7_5 <= _GEN_61;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2374 & _GEN_2275) begin // @[stationary_dpe.scala 95:32]
          Station2_7_6 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_7_6 <= _GEN_62;
        end
      end else begin
        Station2_7_6 <= _GEN_62;
      end
    end else begin
      Station2_7_6 <= _GEN_62;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2374 & _GEN_2277) begin // @[stationary_dpe.scala 95:32]
          Station2_7_7 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_7_7 <= _GEN_63;
        end
      end else begin
        Station2_7_7 <= _GEN_63;
      end
    end else begin
      Station2_7_7 <= _GEN_63;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2264 & _GEN_2279) begin // @[stationary_dpe.scala 116:32]
          Station3_0_0 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_0_0 <= _GEN_64;
        end
      end else begin
        Station3_0_0 <= _GEN_64;
      end
    end else begin
      Station3_0_0 <= _GEN_64;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2264 & _GEN_2265) begin // @[stationary_dpe.scala 116:32]
          Station3_0_1 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_0_1 <= _GEN_65;
        end
      end else begin
        Station3_0_1 <= _GEN_65;
      end
    end else begin
      Station3_0_1 <= _GEN_65;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2264 & _GEN_2267) begin // @[stationary_dpe.scala 116:32]
          Station3_0_2 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_0_2 <= _GEN_66;
        end
      end else begin
        Station3_0_2 <= _GEN_66;
      end
    end else begin
      Station3_0_2 <= _GEN_66;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2264 & _GEN_2269) begin // @[stationary_dpe.scala 116:32]
          Station3_0_3 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_0_3 <= _GEN_67;
        end
      end else begin
        Station3_0_3 <= _GEN_67;
      end
    end else begin
      Station3_0_3 <= _GEN_67;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2264 & _GEN_2271) begin // @[stationary_dpe.scala 116:32]
          Station3_0_4 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_0_4 <= _GEN_68;
        end
      end else begin
        Station3_0_4 <= _GEN_68;
      end
    end else begin
      Station3_0_4 <= _GEN_68;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2264 & _GEN_2273) begin // @[stationary_dpe.scala 116:32]
          Station3_0_5 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_0_5 <= _GEN_69;
        end
      end else begin
        Station3_0_5 <= _GEN_69;
      end
    end else begin
      Station3_0_5 <= _GEN_69;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2264 & _GEN_2275) begin // @[stationary_dpe.scala 116:32]
          Station3_0_6 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_0_6 <= _GEN_70;
        end
      end else begin
        Station3_0_6 <= _GEN_70;
      end
    end else begin
      Station3_0_6 <= _GEN_70;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2264 & _GEN_2277) begin // @[stationary_dpe.scala 116:32]
          Station3_0_7 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_0_7 <= _GEN_71;
        end
      end else begin
        Station3_0_7 <= _GEN_71;
      end
    end else begin
      Station3_0_7 <= _GEN_71;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2278 & _GEN_2279) begin // @[stationary_dpe.scala 116:32]
          Station3_1_0 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_1_0 <= _GEN_72;
        end
      end else begin
        Station3_1_0 <= _GEN_72;
      end
    end else begin
      Station3_1_0 <= _GEN_72;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2278 & _GEN_2265) begin // @[stationary_dpe.scala 116:32]
          Station3_1_1 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_1_1 <= _GEN_73;
        end
      end else begin
        Station3_1_1 <= _GEN_73;
      end
    end else begin
      Station3_1_1 <= _GEN_73;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2278 & _GEN_2267) begin // @[stationary_dpe.scala 116:32]
          Station3_1_2 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_1_2 <= _GEN_74;
        end
      end else begin
        Station3_1_2 <= _GEN_74;
      end
    end else begin
      Station3_1_2 <= _GEN_74;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2278 & _GEN_2269) begin // @[stationary_dpe.scala 116:32]
          Station3_1_3 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_1_3 <= _GEN_75;
        end
      end else begin
        Station3_1_3 <= _GEN_75;
      end
    end else begin
      Station3_1_3 <= _GEN_75;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2278 & _GEN_2271) begin // @[stationary_dpe.scala 116:32]
          Station3_1_4 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_1_4 <= _GEN_76;
        end
      end else begin
        Station3_1_4 <= _GEN_76;
      end
    end else begin
      Station3_1_4 <= _GEN_76;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2278 & _GEN_2273) begin // @[stationary_dpe.scala 116:32]
          Station3_1_5 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_1_5 <= _GEN_77;
        end
      end else begin
        Station3_1_5 <= _GEN_77;
      end
    end else begin
      Station3_1_5 <= _GEN_77;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2278 & _GEN_2275) begin // @[stationary_dpe.scala 116:32]
          Station3_1_6 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_1_6 <= _GEN_78;
        end
      end else begin
        Station3_1_6 <= _GEN_78;
      end
    end else begin
      Station3_1_6 <= _GEN_78;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2278 & _GEN_2277) begin // @[stationary_dpe.scala 116:32]
          Station3_1_7 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_1_7 <= _GEN_79;
        end
      end else begin
        Station3_1_7 <= _GEN_79;
      end
    end else begin
      Station3_1_7 <= _GEN_79;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2294 & _GEN_2279) begin // @[stationary_dpe.scala 116:32]
          Station3_2_0 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_2_0 <= _GEN_80;
        end
      end else begin
        Station3_2_0 <= _GEN_80;
      end
    end else begin
      Station3_2_0 <= _GEN_80;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2294 & _GEN_2265) begin // @[stationary_dpe.scala 116:32]
          Station3_2_1 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_2_1 <= _GEN_81;
        end
      end else begin
        Station3_2_1 <= _GEN_81;
      end
    end else begin
      Station3_2_1 <= _GEN_81;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2294 & _GEN_2267) begin // @[stationary_dpe.scala 116:32]
          Station3_2_2 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_2_2 <= _GEN_82;
        end
      end else begin
        Station3_2_2 <= _GEN_82;
      end
    end else begin
      Station3_2_2 <= _GEN_82;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2294 & _GEN_2269) begin // @[stationary_dpe.scala 116:32]
          Station3_2_3 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_2_3 <= _GEN_83;
        end
      end else begin
        Station3_2_3 <= _GEN_83;
      end
    end else begin
      Station3_2_3 <= _GEN_83;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2294 & _GEN_2271) begin // @[stationary_dpe.scala 116:32]
          Station3_2_4 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_2_4 <= _GEN_84;
        end
      end else begin
        Station3_2_4 <= _GEN_84;
      end
    end else begin
      Station3_2_4 <= _GEN_84;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2294 & _GEN_2273) begin // @[stationary_dpe.scala 116:32]
          Station3_2_5 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_2_5 <= _GEN_85;
        end
      end else begin
        Station3_2_5 <= _GEN_85;
      end
    end else begin
      Station3_2_5 <= _GEN_85;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2294 & _GEN_2275) begin // @[stationary_dpe.scala 116:32]
          Station3_2_6 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_2_6 <= _GEN_86;
        end
      end else begin
        Station3_2_6 <= _GEN_86;
      end
    end else begin
      Station3_2_6 <= _GEN_86;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2294 & _GEN_2277) begin // @[stationary_dpe.scala 116:32]
          Station3_2_7 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_2_7 <= _GEN_87;
        end
      end else begin
        Station3_2_7 <= _GEN_87;
      end
    end else begin
      Station3_2_7 <= _GEN_87;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2310 & _GEN_2279) begin // @[stationary_dpe.scala 116:32]
          Station3_3_0 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_3_0 <= _GEN_88;
        end
      end else begin
        Station3_3_0 <= _GEN_88;
      end
    end else begin
      Station3_3_0 <= _GEN_88;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2310 & _GEN_2265) begin // @[stationary_dpe.scala 116:32]
          Station3_3_1 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_3_1 <= _GEN_89;
        end
      end else begin
        Station3_3_1 <= _GEN_89;
      end
    end else begin
      Station3_3_1 <= _GEN_89;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2310 & _GEN_2267) begin // @[stationary_dpe.scala 116:32]
          Station3_3_2 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_3_2 <= _GEN_90;
        end
      end else begin
        Station3_3_2 <= _GEN_90;
      end
    end else begin
      Station3_3_2 <= _GEN_90;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2310 & _GEN_2269) begin // @[stationary_dpe.scala 116:32]
          Station3_3_3 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_3_3 <= _GEN_91;
        end
      end else begin
        Station3_3_3 <= _GEN_91;
      end
    end else begin
      Station3_3_3 <= _GEN_91;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2310 & _GEN_2271) begin // @[stationary_dpe.scala 116:32]
          Station3_3_4 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_3_4 <= _GEN_92;
        end
      end else begin
        Station3_3_4 <= _GEN_92;
      end
    end else begin
      Station3_3_4 <= _GEN_92;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2310 & _GEN_2273) begin // @[stationary_dpe.scala 116:32]
          Station3_3_5 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_3_5 <= _GEN_93;
        end
      end else begin
        Station3_3_5 <= _GEN_93;
      end
    end else begin
      Station3_3_5 <= _GEN_93;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2310 & _GEN_2275) begin // @[stationary_dpe.scala 116:32]
          Station3_3_6 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_3_6 <= _GEN_94;
        end
      end else begin
        Station3_3_6 <= _GEN_94;
      end
    end else begin
      Station3_3_6 <= _GEN_94;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2310 & _GEN_2277) begin // @[stationary_dpe.scala 116:32]
          Station3_3_7 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_3_7 <= _GEN_95;
        end
      end else begin
        Station3_3_7 <= _GEN_95;
      end
    end else begin
      Station3_3_7 <= _GEN_95;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2326 & _GEN_2279) begin // @[stationary_dpe.scala 116:32]
          Station3_4_0 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_4_0 <= _GEN_96;
        end
      end else begin
        Station3_4_0 <= _GEN_96;
      end
    end else begin
      Station3_4_0 <= _GEN_96;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2326 & _GEN_2265) begin // @[stationary_dpe.scala 116:32]
          Station3_4_1 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_4_1 <= _GEN_97;
        end
      end else begin
        Station3_4_1 <= _GEN_97;
      end
    end else begin
      Station3_4_1 <= _GEN_97;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2326 & _GEN_2267) begin // @[stationary_dpe.scala 116:32]
          Station3_4_2 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_4_2 <= _GEN_98;
        end
      end else begin
        Station3_4_2 <= _GEN_98;
      end
    end else begin
      Station3_4_2 <= _GEN_98;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2326 & _GEN_2269) begin // @[stationary_dpe.scala 116:32]
          Station3_4_3 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_4_3 <= _GEN_99;
        end
      end else begin
        Station3_4_3 <= _GEN_99;
      end
    end else begin
      Station3_4_3 <= _GEN_99;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2326 & _GEN_2271) begin // @[stationary_dpe.scala 116:32]
          Station3_4_4 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_4_4 <= _GEN_100;
        end
      end else begin
        Station3_4_4 <= _GEN_100;
      end
    end else begin
      Station3_4_4 <= _GEN_100;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2326 & _GEN_2273) begin // @[stationary_dpe.scala 116:32]
          Station3_4_5 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_4_5 <= _GEN_101;
        end
      end else begin
        Station3_4_5 <= _GEN_101;
      end
    end else begin
      Station3_4_5 <= _GEN_101;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2326 & _GEN_2275) begin // @[stationary_dpe.scala 116:32]
          Station3_4_6 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_4_6 <= _GEN_102;
        end
      end else begin
        Station3_4_6 <= _GEN_102;
      end
    end else begin
      Station3_4_6 <= _GEN_102;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2326 & _GEN_2277) begin // @[stationary_dpe.scala 116:32]
          Station3_4_7 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_4_7 <= _GEN_103;
        end
      end else begin
        Station3_4_7 <= _GEN_103;
      end
    end else begin
      Station3_4_7 <= _GEN_103;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2342 & _GEN_2279) begin // @[stationary_dpe.scala 116:32]
          Station3_5_0 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_5_0 <= _GEN_104;
        end
      end else begin
        Station3_5_0 <= _GEN_104;
      end
    end else begin
      Station3_5_0 <= _GEN_104;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2342 & _GEN_2265) begin // @[stationary_dpe.scala 116:32]
          Station3_5_1 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_5_1 <= _GEN_105;
        end
      end else begin
        Station3_5_1 <= _GEN_105;
      end
    end else begin
      Station3_5_1 <= _GEN_105;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2342 & _GEN_2267) begin // @[stationary_dpe.scala 116:32]
          Station3_5_2 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_5_2 <= _GEN_106;
        end
      end else begin
        Station3_5_2 <= _GEN_106;
      end
    end else begin
      Station3_5_2 <= _GEN_106;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2342 & _GEN_2269) begin // @[stationary_dpe.scala 116:32]
          Station3_5_3 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_5_3 <= _GEN_107;
        end
      end else begin
        Station3_5_3 <= _GEN_107;
      end
    end else begin
      Station3_5_3 <= _GEN_107;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2342 & _GEN_2271) begin // @[stationary_dpe.scala 116:32]
          Station3_5_4 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_5_4 <= _GEN_108;
        end
      end else begin
        Station3_5_4 <= _GEN_108;
      end
    end else begin
      Station3_5_4 <= _GEN_108;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2342 & _GEN_2273) begin // @[stationary_dpe.scala 116:32]
          Station3_5_5 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_5_5 <= _GEN_109;
        end
      end else begin
        Station3_5_5 <= _GEN_109;
      end
    end else begin
      Station3_5_5 <= _GEN_109;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2342 & _GEN_2275) begin // @[stationary_dpe.scala 116:32]
          Station3_5_6 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_5_6 <= _GEN_110;
        end
      end else begin
        Station3_5_6 <= _GEN_110;
      end
    end else begin
      Station3_5_6 <= _GEN_110;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2342 & _GEN_2277) begin // @[stationary_dpe.scala 116:32]
          Station3_5_7 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_5_7 <= _GEN_111;
        end
      end else begin
        Station3_5_7 <= _GEN_111;
      end
    end else begin
      Station3_5_7 <= _GEN_111;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2358 & _GEN_2279) begin // @[stationary_dpe.scala 116:32]
          Station3_6_0 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_6_0 <= _GEN_112;
        end
      end else begin
        Station3_6_0 <= _GEN_112;
      end
    end else begin
      Station3_6_0 <= _GEN_112;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2358 & _GEN_2265) begin // @[stationary_dpe.scala 116:32]
          Station3_6_1 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_6_1 <= _GEN_113;
        end
      end else begin
        Station3_6_1 <= _GEN_113;
      end
    end else begin
      Station3_6_1 <= _GEN_113;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2358 & _GEN_2267) begin // @[stationary_dpe.scala 116:32]
          Station3_6_2 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_6_2 <= _GEN_114;
        end
      end else begin
        Station3_6_2 <= _GEN_114;
      end
    end else begin
      Station3_6_2 <= _GEN_114;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2358 & _GEN_2269) begin // @[stationary_dpe.scala 116:32]
          Station3_6_3 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_6_3 <= _GEN_115;
        end
      end else begin
        Station3_6_3 <= _GEN_115;
      end
    end else begin
      Station3_6_3 <= _GEN_115;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2358 & _GEN_2271) begin // @[stationary_dpe.scala 116:32]
          Station3_6_4 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_6_4 <= _GEN_116;
        end
      end else begin
        Station3_6_4 <= _GEN_116;
      end
    end else begin
      Station3_6_4 <= _GEN_116;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2358 & _GEN_2273) begin // @[stationary_dpe.scala 116:32]
          Station3_6_5 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_6_5 <= _GEN_117;
        end
      end else begin
        Station3_6_5 <= _GEN_117;
      end
    end else begin
      Station3_6_5 <= _GEN_117;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2358 & _GEN_2275) begin // @[stationary_dpe.scala 116:32]
          Station3_6_6 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_6_6 <= _GEN_118;
        end
      end else begin
        Station3_6_6 <= _GEN_118;
      end
    end else begin
      Station3_6_6 <= _GEN_118;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2358 & _GEN_2277) begin // @[stationary_dpe.scala 116:32]
          Station3_6_7 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_6_7 <= _GEN_119;
        end
      end else begin
        Station3_6_7 <= _GEN_119;
      end
    end else begin
      Station3_6_7 <= _GEN_119;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2374 & _GEN_2279) begin // @[stationary_dpe.scala 116:32]
          Station3_7_0 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_7_0 <= _GEN_120;
        end
      end else begin
        Station3_7_0 <= _GEN_120;
      end
    end else begin
      Station3_7_0 <= _GEN_120;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2374 & _GEN_2265) begin // @[stationary_dpe.scala 116:32]
          Station3_7_1 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_7_1 <= _GEN_121;
        end
      end else begin
        Station3_7_1 <= _GEN_121;
      end
    end else begin
      Station3_7_1 <= _GEN_121;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2374 & _GEN_2267) begin // @[stationary_dpe.scala 116:32]
          Station3_7_2 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_7_2 <= _GEN_122;
        end
      end else begin
        Station3_7_2 <= _GEN_122;
      end
    end else begin
      Station3_7_2 <= _GEN_122;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2374 & _GEN_2269) begin // @[stationary_dpe.scala 116:32]
          Station3_7_3 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_7_3 <= _GEN_123;
        end
      end else begin
        Station3_7_3 <= _GEN_123;
      end
    end else begin
      Station3_7_3 <= _GEN_123;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2374 & _GEN_2271) begin // @[stationary_dpe.scala 116:32]
          Station3_7_4 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_7_4 <= _GEN_124;
        end
      end else begin
        Station3_7_4 <= _GEN_124;
      end
    end else begin
      Station3_7_4 <= _GEN_124;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2374 & _GEN_2273) begin // @[stationary_dpe.scala 116:32]
          Station3_7_5 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_7_5 <= _GEN_125;
        end
      end else begin
        Station3_7_5 <= _GEN_125;
      end
    end else begin
      Station3_7_5 <= _GEN_125;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2374 & _GEN_2275) begin // @[stationary_dpe.scala 116:32]
          Station3_7_6 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_7_6 <= _GEN_126;
        end
      end else begin
        Station3_7_6 <= _GEN_126;
      end
    end else begin
      Station3_7_6 <= _GEN_126;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2374 & _GEN_2277) begin // @[stationary_dpe.scala 116:32]
          Station3_7_7 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_7_7 <= _GEN_127;
        end
      end else begin
        Station3_7_7 <= _GEN_127;
      end
    end else begin
      Station3_7_7 <= _GEN_127;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2264 & _GEN_2279) begin // @[stationary_dpe.scala 128:32]
          Station4_0_0 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_0_0 <= _GEN_128;
        end
      end else begin
        Station4_0_0 <= _GEN_128;
      end
    end else begin
      Station4_0_0 <= _GEN_128;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2264 & _GEN_2265) begin // @[stationary_dpe.scala 128:32]
          Station4_0_1 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_0_1 <= _GEN_129;
        end
      end else begin
        Station4_0_1 <= _GEN_129;
      end
    end else begin
      Station4_0_1 <= _GEN_129;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2264 & _GEN_2267) begin // @[stationary_dpe.scala 128:32]
          Station4_0_2 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_0_2 <= _GEN_130;
        end
      end else begin
        Station4_0_2 <= _GEN_130;
      end
    end else begin
      Station4_0_2 <= _GEN_130;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2264 & _GEN_2269) begin // @[stationary_dpe.scala 128:32]
          Station4_0_3 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_0_3 <= _GEN_131;
        end
      end else begin
        Station4_0_3 <= _GEN_131;
      end
    end else begin
      Station4_0_3 <= _GEN_131;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2264 & _GEN_2271) begin // @[stationary_dpe.scala 128:32]
          Station4_0_4 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_0_4 <= _GEN_132;
        end
      end else begin
        Station4_0_4 <= _GEN_132;
      end
    end else begin
      Station4_0_4 <= _GEN_132;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2264 & _GEN_2273) begin // @[stationary_dpe.scala 128:32]
          Station4_0_5 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_0_5 <= _GEN_133;
        end
      end else begin
        Station4_0_5 <= _GEN_133;
      end
    end else begin
      Station4_0_5 <= _GEN_133;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2264 & _GEN_2275) begin // @[stationary_dpe.scala 128:32]
          Station4_0_6 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_0_6 <= _GEN_134;
        end
      end else begin
        Station4_0_6 <= _GEN_134;
      end
    end else begin
      Station4_0_6 <= _GEN_134;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2264 & _GEN_2277) begin // @[stationary_dpe.scala 128:32]
          Station4_0_7 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_0_7 <= _GEN_135;
        end
      end else begin
        Station4_0_7 <= _GEN_135;
      end
    end else begin
      Station4_0_7 <= _GEN_135;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2278 & _GEN_2279) begin // @[stationary_dpe.scala 128:32]
          Station4_1_0 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_1_0 <= _GEN_136;
        end
      end else begin
        Station4_1_0 <= _GEN_136;
      end
    end else begin
      Station4_1_0 <= _GEN_136;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2278 & _GEN_2265) begin // @[stationary_dpe.scala 128:32]
          Station4_1_1 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_1_1 <= _GEN_137;
        end
      end else begin
        Station4_1_1 <= _GEN_137;
      end
    end else begin
      Station4_1_1 <= _GEN_137;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2278 & _GEN_2267) begin // @[stationary_dpe.scala 128:32]
          Station4_1_2 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_1_2 <= _GEN_138;
        end
      end else begin
        Station4_1_2 <= _GEN_138;
      end
    end else begin
      Station4_1_2 <= _GEN_138;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2278 & _GEN_2269) begin // @[stationary_dpe.scala 128:32]
          Station4_1_3 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_1_3 <= _GEN_139;
        end
      end else begin
        Station4_1_3 <= _GEN_139;
      end
    end else begin
      Station4_1_3 <= _GEN_139;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2278 & _GEN_2271) begin // @[stationary_dpe.scala 128:32]
          Station4_1_4 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_1_4 <= _GEN_140;
        end
      end else begin
        Station4_1_4 <= _GEN_140;
      end
    end else begin
      Station4_1_4 <= _GEN_140;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2278 & _GEN_2273) begin // @[stationary_dpe.scala 128:32]
          Station4_1_5 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_1_5 <= _GEN_141;
        end
      end else begin
        Station4_1_5 <= _GEN_141;
      end
    end else begin
      Station4_1_5 <= _GEN_141;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2278 & _GEN_2275) begin // @[stationary_dpe.scala 128:32]
          Station4_1_6 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_1_6 <= _GEN_142;
        end
      end else begin
        Station4_1_6 <= _GEN_142;
      end
    end else begin
      Station4_1_6 <= _GEN_142;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2278 & _GEN_2277) begin // @[stationary_dpe.scala 128:32]
          Station4_1_7 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_1_7 <= _GEN_143;
        end
      end else begin
        Station4_1_7 <= _GEN_143;
      end
    end else begin
      Station4_1_7 <= _GEN_143;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2294 & _GEN_2279) begin // @[stationary_dpe.scala 128:32]
          Station4_2_0 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_2_0 <= _GEN_144;
        end
      end else begin
        Station4_2_0 <= _GEN_144;
      end
    end else begin
      Station4_2_0 <= _GEN_144;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2294 & _GEN_2265) begin // @[stationary_dpe.scala 128:32]
          Station4_2_1 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_2_1 <= _GEN_145;
        end
      end else begin
        Station4_2_1 <= _GEN_145;
      end
    end else begin
      Station4_2_1 <= _GEN_145;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2294 & _GEN_2267) begin // @[stationary_dpe.scala 128:32]
          Station4_2_2 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_2_2 <= _GEN_146;
        end
      end else begin
        Station4_2_2 <= _GEN_146;
      end
    end else begin
      Station4_2_2 <= _GEN_146;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2294 & _GEN_2269) begin // @[stationary_dpe.scala 128:32]
          Station4_2_3 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_2_3 <= _GEN_147;
        end
      end else begin
        Station4_2_3 <= _GEN_147;
      end
    end else begin
      Station4_2_3 <= _GEN_147;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2294 & _GEN_2271) begin // @[stationary_dpe.scala 128:32]
          Station4_2_4 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_2_4 <= _GEN_148;
        end
      end else begin
        Station4_2_4 <= _GEN_148;
      end
    end else begin
      Station4_2_4 <= _GEN_148;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2294 & _GEN_2273) begin // @[stationary_dpe.scala 128:32]
          Station4_2_5 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_2_5 <= _GEN_149;
        end
      end else begin
        Station4_2_5 <= _GEN_149;
      end
    end else begin
      Station4_2_5 <= _GEN_149;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2294 & _GEN_2275) begin // @[stationary_dpe.scala 128:32]
          Station4_2_6 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_2_6 <= _GEN_150;
        end
      end else begin
        Station4_2_6 <= _GEN_150;
      end
    end else begin
      Station4_2_6 <= _GEN_150;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2294 & _GEN_2277) begin // @[stationary_dpe.scala 128:32]
          Station4_2_7 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_2_7 <= _GEN_151;
        end
      end else begin
        Station4_2_7 <= _GEN_151;
      end
    end else begin
      Station4_2_7 <= _GEN_151;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2310 & _GEN_2279) begin // @[stationary_dpe.scala 128:32]
          Station4_3_0 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_3_0 <= _GEN_152;
        end
      end else begin
        Station4_3_0 <= _GEN_152;
      end
    end else begin
      Station4_3_0 <= _GEN_152;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2310 & _GEN_2265) begin // @[stationary_dpe.scala 128:32]
          Station4_3_1 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_3_1 <= _GEN_153;
        end
      end else begin
        Station4_3_1 <= _GEN_153;
      end
    end else begin
      Station4_3_1 <= _GEN_153;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2310 & _GEN_2267) begin // @[stationary_dpe.scala 128:32]
          Station4_3_2 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_3_2 <= _GEN_154;
        end
      end else begin
        Station4_3_2 <= _GEN_154;
      end
    end else begin
      Station4_3_2 <= _GEN_154;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2310 & _GEN_2269) begin // @[stationary_dpe.scala 128:32]
          Station4_3_3 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_3_3 <= _GEN_155;
        end
      end else begin
        Station4_3_3 <= _GEN_155;
      end
    end else begin
      Station4_3_3 <= _GEN_155;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2310 & _GEN_2271) begin // @[stationary_dpe.scala 128:32]
          Station4_3_4 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_3_4 <= _GEN_156;
        end
      end else begin
        Station4_3_4 <= _GEN_156;
      end
    end else begin
      Station4_3_4 <= _GEN_156;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2310 & _GEN_2273) begin // @[stationary_dpe.scala 128:32]
          Station4_3_5 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_3_5 <= _GEN_157;
        end
      end else begin
        Station4_3_5 <= _GEN_157;
      end
    end else begin
      Station4_3_5 <= _GEN_157;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2310 & _GEN_2275) begin // @[stationary_dpe.scala 128:32]
          Station4_3_6 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_3_6 <= _GEN_158;
        end
      end else begin
        Station4_3_6 <= _GEN_158;
      end
    end else begin
      Station4_3_6 <= _GEN_158;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2310 & _GEN_2277) begin // @[stationary_dpe.scala 128:32]
          Station4_3_7 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_3_7 <= _GEN_159;
        end
      end else begin
        Station4_3_7 <= _GEN_159;
      end
    end else begin
      Station4_3_7 <= _GEN_159;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2326 & _GEN_2279) begin // @[stationary_dpe.scala 128:32]
          Station4_4_0 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_4_0 <= _GEN_160;
        end
      end else begin
        Station4_4_0 <= _GEN_160;
      end
    end else begin
      Station4_4_0 <= _GEN_160;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2326 & _GEN_2265) begin // @[stationary_dpe.scala 128:32]
          Station4_4_1 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_4_1 <= _GEN_161;
        end
      end else begin
        Station4_4_1 <= _GEN_161;
      end
    end else begin
      Station4_4_1 <= _GEN_161;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2326 & _GEN_2267) begin // @[stationary_dpe.scala 128:32]
          Station4_4_2 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_4_2 <= _GEN_162;
        end
      end else begin
        Station4_4_2 <= _GEN_162;
      end
    end else begin
      Station4_4_2 <= _GEN_162;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2326 & _GEN_2269) begin // @[stationary_dpe.scala 128:32]
          Station4_4_3 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_4_3 <= _GEN_163;
        end
      end else begin
        Station4_4_3 <= _GEN_163;
      end
    end else begin
      Station4_4_3 <= _GEN_163;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2326 & _GEN_2271) begin // @[stationary_dpe.scala 128:32]
          Station4_4_4 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_4_4 <= _GEN_164;
        end
      end else begin
        Station4_4_4 <= _GEN_164;
      end
    end else begin
      Station4_4_4 <= _GEN_164;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2326 & _GEN_2273) begin // @[stationary_dpe.scala 128:32]
          Station4_4_5 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_4_5 <= _GEN_165;
        end
      end else begin
        Station4_4_5 <= _GEN_165;
      end
    end else begin
      Station4_4_5 <= _GEN_165;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2326 & _GEN_2275) begin // @[stationary_dpe.scala 128:32]
          Station4_4_6 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_4_6 <= _GEN_166;
        end
      end else begin
        Station4_4_6 <= _GEN_166;
      end
    end else begin
      Station4_4_6 <= _GEN_166;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2326 & _GEN_2277) begin // @[stationary_dpe.scala 128:32]
          Station4_4_7 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_4_7 <= _GEN_167;
        end
      end else begin
        Station4_4_7 <= _GEN_167;
      end
    end else begin
      Station4_4_7 <= _GEN_167;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2342 & _GEN_2279) begin // @[stationary_dpe.scala 128:32]
          Station4_5_0 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_5_0 <= _GEN_168;
        end
      end else begin
        Station4_5_0 <= _GEN_168;
      end
    end else begin
      Station4_5_0 <= _GEN_168;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2342 & _GEN_2265) begin // @[stationary_dpe.scala 128:32]
          Station4_5_1 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_5_1 <= _GEN_169;
        end
      end else begin
        Station4_5_1 <= _GEN_169;
      end
    end else begin
      Station4_5_1 <= _GEN_169;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2342 & _GEN_2267) begin // @[stationary_dpe.scala 128:32]
          Station4_5_2 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_5_2 <= _GEN_170;
        end
      end else begin
        Station4_5_2 <= _GEN_170;
      end
    end else begin
      Station4_5_2 <= _GEN_170;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2342 & _GEN_2269) begin // @[stationary_dpe.scala 128:32]
          Station4_5_3 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_5_3 <= _GEN_171;
        end
      end else begin
        Station4_5_3 <= _GEN_171;
      end
    end else begin
      Station4_5_3 <= _GEN_171;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2342 & _GEN_2271) begin // @[stationary_dpe.scala 128:32]
          Station4_5_4 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_5_4 <= _GEN_172;
        end
      end else begin
        Station4_5_4 <= _GEN_172;
      end
    end else begin
      Station4_5_4 <= _GEN_172;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2342 & _GEN_2273) begin // @[stationary_dpe.scala 128:32]
          Station4_5_5 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_5_5 <= _GEN_173;
        end
      end else begin
        Station4_5_5 <= _GEN_173;
      end
    end else begin
      Station4_5_5 <= _GEN_173;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2342 & _GEN_2275) begin // @[stationary_dpe.scala 128:32]
          Station4_5_6 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_5_6 <= _GEN_174;
        end
      end else begin
        Station4_5_6 <= _GEN_174;
      end
    end else begin
      Station4_5_6 <= _GEN_174;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2342 & _GEN_2277) begin // @[stationary_dpe.scala 128:32]
          Station4_5_7 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_5_7 <= _GEN_175;
        end
      end else begin
        Station4_5_7 <= _GEN_175;
      end
    end else begin
      Station4_5_7 <= _GEN_175;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2358 & _GEN_2279) begin // @[stationary_dpe.scala 128:32]
          Station4_6_0 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_6_0 <= _GEN_176;
        end
      end else begin
        Station4_6_0 <= _GEN_176;
      end
    end else begin
      Station4_6_0 <= _GEN_176;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2358 & _GEN_2265) begin // @[stationary_dpe.scala 128:32]
          Station4_6_1 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_6_1 <= _GEN_177;
        end
      end else begin
        Station4_6_1 <= _GEN_177;
      end
    end else begin
      Station4_6_1 <= _GEN_177;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2358 & _GEN_2267) begin // @[stationary_dpe.scala 128:32]
          Station4_6_2 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_6_2 <= _GEN_178;
        end
      end else begin
        Station4_6_2 <= _GEN_178;
      end
    end else begin
      Station4_6_2 <= _GEN_178;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2358 & _GEN_2269) begin // @[stationary_dpe.scala 128:32]
          Station4_6_3 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_6_3 <= _GEN_179;
        end
      end else begin
        Station4_6_3 <= _GEN_179;
      end
    end else begin
      Station4_6_3 <= _GEN_179;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2358 & _GEN_2271) begin // @[stationary_dpe.scala 128:32]
          Station4_6_4 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_6_4 <= _GEN_180;
        end
      end else begin
        Station4_6_4 <= _GEN_180;
      end
    end else begin
      Station4_6_4 <= _GEN_180;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2358 & _GEN_2273) begin // @[stationary_dpe.scala 128:32]
          Station4_6_5 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_6_5 <= _GEN_181;
        end
      end else begin
        Station4_6_5 <= _GEN_181;
      end
    end else begin
      Station4_6_5 <= _GEN_181;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2358 & _GEN_2275) begin // @[stationary_dpe.scala 128:32]
          Station4_6_6 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_6_6 <= _GEN_182;
        end
      end else begin
        Station4_6_6 <= _GEN_182;
      end
    end else begin
      Station4_6_6 <= _GEN_182;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2358 & _GEN_2277) begin // @[stationary_dpe.scala 128:32]
          Station4_6_7 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_6_7 <= _GEN_183;
        end
      end else begin
        Station4_6_7 <= _GEN_183;
      end
    end else begin
      Station4_6_7 <= _GEN_183;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2374 & _GEN_2279) begin // @[stationary_dpe.scala 128:32]
          Station4_7_0 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_7_0 <= _GEN_184;
        end
      end else begin
        Station4_7_0 <= _GEN_184;
      end
    end else begin
      Station4_7_0 <= _GEN_184;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2374 & _GEN_2265) begin // @[stationary_dpe.scala 128:32]
          Station4_7_1 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_7_1 <= _GEN_185;
        end
      end else begin
        Station4_7_1 <= _GEN_185;
      end
    end else begin
      Station4_7_1 <= _GEN_185;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2374 & _GEN_2267) begin // @[stationary_dpe.scala 128:32]
          Station4_7_2 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_7_2 <= _GEN_186;
        end
      end else begin
        Station4_7_2 <= _GEN_186;
      end
    end else begin
      Station4_7_2 <= _GEN_186;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2374 & _GEN_2269) begin // @[stationary_dpe.scala 128:32]
          Station4_7_3 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_7_3 <= _GEN_187;
        end
      end else begin
        Station4_7_3 <= _GEN_187;
      end
    end else begin
      Station4_7_3 <= _GEN_187;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2374 & _GEN_2271) begin // @[stationary_dpe.scala 128:32]
          Station4_7_4 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_7_4 <= _GEN_188;
        end
      end else begin
        Station4_7_4 <= _GEN_188;
      end
    end else begin
      Station4_7_4 <= _GEN_188;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2374 & _GEN_2273) begin // @[stationary_dpe.scala 128:32]
          Station4_7_5 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_7_5 <= _GEN_189;
        end
      end else begin
        Station4_7_5 <= _GEN_189;
      end
    end else begin
      Station4_7_5 <= _GEN_189;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2374 & _GEN_2275) begin // @[stationary_dpe.scala 128:32]
          Station4_7_6 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_7_6 <= _GEN_190;
        end
      end else begin
        Station4_7_6 <= _GEN_190;
      end
    end else begin
      Station4_7_6 <= _GEN_190;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2374 & _GEN_2277) begin // @[stationary_dpe.scala 128:32]
          Station4_7_7 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_7_7 <= _GEN_191;
        end
      end else begin
        Station4_7_7 <= _GEN_191;
      end
    end else begin
      Station4_7_7 <= _GEN_191;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2264 & _GEN_2279) begin // @[stationary_dpe.scala 140:32]
          Station5_0_0 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_0_0 <= _GEN_192;
        end
      end else begin
        Station5_0_0 <= _GEN_192;
      end
    end else begin
      Station5_0_0 <= _GEN_192;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2264 & _GEN_2265) begin // @[stationary_dpe.scala 140:32]
          Station5_0_1 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_0_1 <= _GEN_193;
        end
      end else begin
        Station5_0_1 <= _GEN_193;
      end
    end else begin
      Station5_0_1 <= _GEN_193;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2264 & _GEN_2267) begin // @[stationary_dpe.scala 140:32]
          Station5_0_2 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_0_2 <= _GEN_194;
        end
      end else begin
        Station5_0_2 <= _GEN_194;
      end
    end else begin
      Station5_0_2 <= _GEN_194;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2264 & _GEN_2269) begin // @[stationary_dpe.scala 140:32]
          Station5_0_3 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_0_3 <= _GEN_195;
        end
      end else begin
        Station5_0_3 <= _GEN_195;
      end
    end else begin
      Station5_0_3 <= _GEN_195;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2264 & _GEN_2271) begin // @[stationary_dpe.scala 140:32]
          Station5_0_4 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_0_4 <= _GEN_196;
        end
      end else begin
        Station5_0_4 <= _GEN_196;
      end
    end else begin
      Station5_0_4 <= _GEN_196;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2264 & _GEN_2273) begin // @[stationary_dpe.scala 140:32]
          Station5_0_5 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_0_5 <= _GEN_197;
        end
      end else begin
        Station5_0_5 <= _GEN_197;
      end
    end else begin
      Station5_0_5 <= _GEN_197;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2264 & _GEN_2275) begin // @[stationary_dpe.scala 140:32]
          Station5_0_6 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_0_6 <= _GEN_198;
        end
      end else begin
        Station5_0_6 <= _GEN_198;
      end
    end else begin
      Station5_0_6 <= _GEN_198;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2264 & _GEN_2277) begin // @[stationary_dpe.scala 140:32]
          Station5_0_7 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_0_7 <= _GEN_199;
        end
      end else begin
        Station5_0_7 <= _GEN_199;
      end
    end else begin
      Station5_0_7 <= _GEN_199;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2278 & _GEN_2279) begin // @[stationary_dpe.scala 140:32]
          Station5_1_0 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_1_0 <= _GEN_200;
        end
      end else begin
        Station5_1_0 <= _GEN_200;
      end
    end else begin
      Station5_1_0 <= _GEN_200;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2278 & _GEN_2265) begin // @[stationary_dpe.scala 140:32]
          Station5_1_1 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_1_1 <= _GEN_201;
        end
      end else begin
        Station5_1_1 <= _GEN_201;
      end
    end else begin
      Station5_1_1 <= _GEN_201;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2278 & _GEN_2267) begin // @[stationary_dpe.scala 140:32]
          Station5_1_2 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_1_2 <= _GEN_202;
        end
      end else begin
        Station5_1_2 <= _GEN_202;
      end
    end else begin
      Station5_1_2 <= _GEN_202;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2278 & _GEN_2269) begin // @[stationary_dpe.scala 140:32]
          Station5_1_3 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_1_3 <= _GEN_203;
        end
      end else begin
        Station5_1_3 <= _GEN_203;
      end
    end else begin
      Station5_1_3 <= _GEN_203;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2278 & _GEN_2271) begin // @[stationary_dpe.scala 140:32]
          Station5_1_4 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_1_4 <= _GEN_204;
        end
      end else begin
        Station5_1_4 <= _GEN_204;
      end
    end else begin
      Station5_1_4 <= _GEN_204;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2278 & _GEN_2273) begin // @[stationary_dpe.scala 140:32]
          Station5_1_5 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_1_5 <= _GEN_205;
        end
      end else begin
        Station5_1_5 <= _GEN_205;
      end
    end else begin
      Station5_1_5 <= _GEN_205;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2278 & _GEN_2275) begin // @[stationary_dpe.scala 140:32]
          Station5_1_6 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_1_6 <= _GEN_206;
        end
      end else begin
        Station5_1_6 <= _GEN_206;
      end
    end else begin
      Station5_1_6 <= _GEN_206;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2278 & _GEN_2277) begin // @[stationary_dpe.scala 140:32]
          Station5_1_7 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_1_7 <= _GEN_207;
        end
      end else begin
        Station5_1_7 <= _GEN_207;
      end
    end else begin
      Station5_1_7 <= _GEN_207;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2294 & _GEN_2279) begin // @[stationary_dpe.scala 140:32]
          Station5_2_0 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_2_0 <= _GEN_208;
        end
      end else begin
        Station5_2_0 <= _GEN_208;
      end
    end else begin
      Station5_2_0 <= _GEN_208;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2294 & _GEN_2265) begin // @[stationary_dpe.scala 140:32]
          Station5_2_1 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_2_1 <= _GEN_209;
        end
      end else begin
        Station5_2_1 <= _GEN_209;
      end
    end else begin
      Station5_2_1 <= _GEN_209;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2294 & _GEN_2267) begin // @[stationary_dpe.scala 140:32]
          Station5_2_2 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_2_2 <= _GEN_210;
        end
      end else begin
        Station5_2_2 <= _GEN_210;
      end
    end else begin
      Station5_2_2 <= _GEN_210;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2294 & _GEN_2269) begin // @[stationary_dpe.scala 140:32]
          Station5_2_3 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_2_3 <= _GEN_211;
        end
      end else begin
        Station5_2_3 <= _GEN_211;
      end
    end else begin
      Station5_2_3 <= _GEN_211;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2294 & _GEN_2271) begin // @[stationary_dpe.scala 140:32]
          Station5_2_4 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_2_4 <= _GEN_212;
        end
      end else begin
        Station5_2_4 <= _GEN_212;
      end
    end else begin
      Station5_2_4 <= _GEN_212;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2294 & _GEN_2273) begin // @[stationary_dpe.scala 140:32]
          Station5_2_5 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_2_5 <= _GEN_213;
        end
      end else begin
        Station5_2_5 <= _GEN_213;
      end
    end else begin
      Station5_2_5 <= _GEN_213;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2294 & _GEN_2275) begin // @[stationary_dpe.scala 140:32]
          Station5_2_6 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_2_6 <= _GEN_214;
        end
      end else begin
        Station5_2_6 <= _GEN_214;
      end
    end else begin
      Station5_2_6 <= _GEN_214;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2294 & _GEN_2277) begin // @[stationary_dpe.scala 140:32]
          Station5_2_7 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_2_7 <= _GEN_215;
        end
      end else begin
        Station5_2_7 <= _GEN_215;
      end
    end else begin
      Station5_2_7 <= _GEN_215;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2310 & _GEN_2279) begin // @[stationary_dpe.scala 140:32]
          Station5_3_0 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_3_0 <= _GEN_216;
        end
      end else begin
        Station5_3_0 <= _GEN_216;
      end
    end else begin
      Station5_3_0 <= _GEN_216;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2310 & _GEN_2265) begin // @[stationary_dpe.scala 140:32]
          Station5_3_1 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_3_1 <= _GEN_217;
        end
      end else begin
        Station5_3_1 <= _GEN_217;
      end
    end else begin
      Station5_3_1 <= _GEN_217;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2310 & _GEN_2267) begin // @[stationary_dpe.scala 140:32]
          Station5_3_2 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_3_2 <= _GEN_218;
        end
      end else begin
        Station5_3_2 <= _GEN_218;
      end
    end else begin
      Station5_3_2 <= _GEN_218;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2310 & _GEN_2269) begin // @[stationary_dpe.scala 140:32]
          Station5_3_3 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_3_3 <= _GEN_219;
        end
      end else begin
        Station5_3_3 <= _GEN_219;
      end
    end else begin
      Station5_3_3 <= _GEN_219;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2310 & _GEN_2271) begin // @[stationary_dpe.scala 140:32]
          Station5_3_4 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_3_4 <= _GEN_220;
        end
      end else begin
        Station5_3_4 <= _GEN_220;
      end
    end else begin
      Station5_3_4 <= _GEN_220;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2310 & _GEN_2273) begin // @[stationary_dpe.scala 140:32]
          Station5_3_5 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_3_5 <= _GEN_221;
        end
      end else begin
        Station5_3_5 <= _GEN_221;
      end
    end else begin
      Station5_3_5 <= _GEN_221;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2310 & _GEN_2275) begin // @[stationary_dpe.scala 140:32]
          Station5_3_6 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_3_6 <= _GEN_222;
        end
      end else begin
        Station5_3_6 <= _GEN_222;
      end
    end else begin
      Station5_3_6 <= _GEN_222;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2310 & _GEN_2277) begin // @[stationary_dpe.scala 140:32]
          Station5_3_7 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_3_7 <= _GEN_223;
        end
      end else begin
        Station5_3_7 <= _GEN_223;
      end
    end else begin
      Station5_3_7 <= _GEN_223;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2326 & _GEN_2279) begin // @[stationary_dpe.scala 140:32]
          Station5_4_0 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_4_0 <= _GEN_224;
        end
      end else begin
        Station5_4_0 <= _GEN_224;
      end
    end else begin
      Station5_4_0 <= _GEN_224;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2326 & _GEN_2265) begin // @[stationary_dpe.scala 140:32]
          Station5_4_1 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_4_1 <= _GEN_225;
        end
      end else begin
        Station5_4_1 <= _GEN_225;
      end
    end else begin
      Station5_4_1 <= _GEN_225;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2326 & _GEN_2267) begin // @[stationary_dpe.scala 140:32]
          Station5_4_2 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_4_2 <= _GEN_226;
        end
      end else begin
        Station5_4_2 <= _GEN_226;
      end
    end else begin
      Station5_4_2 <= _GEN_226;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2326 & _GEN_2269) begin // @[stationary_dpe.scala 140:32]
          Station5_4_3 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_4_3 <= _GEN_227;
        end
      end else begin
        Station5_4_3 <= _GEN_227;
      end
    end else begin
      Station5_4_3 <= _GEN_227;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2326 & _GEN_2271) begin // @[stationary_dpe.scala 140:32]
          Station5_4_4 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_4_4 <= _GEN_228;
        end
      end else begin
        Station5_4_4 <= _GEN_228;
      end
    end else begin
      Station5_4_4 <= _GEN_228;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2326 & _GEN_2273) begin // @[stationary_dpe.scala 140:32]
          Station5_4_5 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_4_5 <= _GEN_229;
        end
      end else begin
        Station5_4_5 <= _GEN_229;
      end
    end else begin
      Station5_4_5 <= _GEN_229;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2326 & _GEN_2275) begin // @[stationary_dpe.scala 140:32]
          Station5_4_6 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_4_6 <= _GEN_230;
        end
      end else begin
        Station5_4_6 <= _GEN_230;
      end
    end else begin
      Station5_4_6 <= _GEN_230;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2326 & _GEN_2277) begin // @[stationary_dpe.scala 140:32]
          Station5_4_7 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_4_7 <= _GEN_231;
        end
      end else begin
        Station5_4_7 <= _GEN_231;
      end
    end else begin
      Station5_4_7 <= _GEN_231;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2342 & _GEN_2279) begin // @[stationary_dpe.scala 140:32]
          Station5_5_0 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_5_0 <= _GEN_232;
        end
      end else begin
        Station5_5_0 <= _GEN_232;
      end
    end else begin
      Station5_5_0 <= _GEN_232;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2342 & _GEN_2265) begin // @[stationary_dpe.scala 140:32]
          Station5_5_1 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_5_1 <= _GEN_233;
        end
      end else begin
        Station5_5_1 <= _GEN_233;
      end
    end else begin
      Station5_5_1 <= _GEN_233;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2342 & _GEN_2267) begin // @[stationary_dpe.scala 140:32]
          Station5_5_2 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_5_2 <= _GEN_234;
        end
      end else begin
        Station5_5_2 <= _GEN_234;
      end
    end else begin
      Station5_5_2 <= _GEN_234;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2342 & _GEN_2269) begin // @[stationary_dpe.scala 140:32]
          Station5_5_3 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_5_3 <= _GEN_235;
        end
      end else begin
        Station5_5_3 <= _GEN_235;
      end
    end else begin
      Station5_5_3 <= _GEN_235;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2342 & _GEN_2271) begin // @[stationary_dpe.scala 140:32]
          Station5_5_4 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_5_4 <= _GEN_236;
        end
      end else begin
        Station5_5_4 <= _GEN_236;
      end
    end else begin
      Station5_5_4 <= _GEN_236;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2342 & _GEN_2273) begin // @[stationary_dpe.scala 140:32]
          Station5_5_5 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_5_5 <= _GEN_237;
        end
      end else begin
        Station5_5_5 <= _GEN_237;
      end
    end else begin
      Station5_5_5 <= _GEN_237;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2342 & _GEN_2275) begin // @[stationary_dpe.scala 140:32]
          Station5_5_6 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_5_6 <= _GEN_238;
        end
      end else begin
        Station5_5_6 <= _GEN_238;
      end
    end else begin
      Station5_5_6 <= _GEN_238;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2342 & _GEN_2277) begin // @[stationary_dpe.scala 140:32]
          Station5_5_7 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_5_7 <= _GEN_239;
        end
      end else begin
        Station5_5_7 <= _GEN_239;
      end
    end else begin
      Station5_5_7 <= _GEN_239;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2358 & _GEN_2279) begin // @[stationary_dpe.scala 140:32]
          Station5_6_0 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_6_0 <= _GEN_240;
        end
      end else begin
        Station5_6_0 <= _GEN_240;
      end
    end else begin
      Station5_6_0 <= _GEN_240;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2358 & _GEN_2265) begin // @[stationary_dpe.scala 140:32]
          Station5_6_1 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_6_1 <= _GEN_241;
        end
      end else begin
        Station5_6_1 <= _GEN_241;
      end
    end else begin
      Station5_6_1 <= _GEN_241;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2358 & _GEN_2267) begin // @[stationary_dpe.scala 140:32]
          Station5_6_2 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_6_2 <= _GEN_242;
        end
      end else begin
        Station5_6_2 <= _GEN_242;
      end
    end else begin
      Station5_6_2 <= _GEN_242;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2358 & _GEN_2269) begin // @[stationary_dpe.scala 140:32]
          Station5_6_3 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_6_3 <= _GEN_243;
        end
      end else begin
        Station5_6_3 <= _GEN_243;
      end
    end else begin
      Station5_6_3 <= _GEN_243;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2358 & _GEN_2271) begin // @[stationary_dpe.scala 140:32]
          Station5_6_4 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_6_4 <= _GEN_244;
        end
      end else begin
        Station5_6_4 <= _GEN_244;
      end
    end else begin
      Station5_6_4 <= _GEN_244;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2358 & _GEN_2273) begin // @[stationary_dpe.scala 140:32]
          Station5_6_5 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_6_5 <= _GEN_245;
        end
      end else begin
        Station5_6_5 <= _GEN_245;
      end
    end else begin
      Station5_6_5 <= _GEN_245;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2358 & _GEN_2275) begin // @[stationary_dpe.scala 140:32]
          Station5_6_6 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_6_6 <= _GEN_246;
        end
      end else begin
        Station5_6_6 <= _GEN_246;
      end
    end else begin
      Station5_6_6 <= _GEN_246;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2358 & _GEN_2277) begin // @[stationary_dpe.scala 140:32]
          Station5_6_7 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_6_7 <= _GEN_247;
        end
      end else begin
        Station5_6_7 <= _GEN_247;
      end
    end else begin
      Station5_6_7 <= _GEN_247;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2374 & _GEN_2279) begin // @[stationary_dpe.scala 140:32]
          Station5_7_0 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_7_0 <= _GEN_248;
        end
      end else begin
        Station5_7_0 <= _GEN_248;
      end
    end else begin
      Station5_7_0 <= _GEN_248;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2374 & _GEN_2265) begin // @[stationary_dpe.scala 140:32]
          Station5_7_1 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_7_1 <= _GEN_249;
        end
      end else begin
        Station5_7_1 <= _GEN_249;
      end
    end else begin
      Station5_7_1 <= _GEN_249;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2374 & _GEN_2267) begin // @[stationary_dpe.scala 140:32]
          Station5_7_2 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_7_2 <= _GEN_250;
        end
      end else begin
        Station5_7_2 <= _GEN_250;
      end
    end else begin
      Station5_7_2 <= _GEN_250;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2374 & _GEN_2269) begin // @[stationary_dpe.scala 140:32]
          Station5_7_3 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_7_3 <= _GEN_251;
        end
      end else begin
        Station5_7_3 <= _GEN_251;
      end
    end else begin
      Station5_7_3 <= _GEN_251;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2374 & _GEN_2271) begin // @[stationary_dpe.scala 140:32]
          Station5_7_4 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_7_4 <= _GEN_252;
        end
      end else begin
        Station5_7_4 <= _GEN_252;
      end
    end else begin
      Station5_7_4 <= _GEN_252;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2374 & _GEN_2273) begin // @[stationary_dpe.scala 140:32]
          Station5_7_5 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_7_5 <= _GEN_253;
        end
      end else begin
        Station5_7_5 <= _GEN_253;
      end
    end else begin
      Station5_7_5 <= _GEN_253;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2374 & _GEN_2275) begin // @[stationary_dpe.scala 140:32]
          Station5_7_6 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_7_6 <= _GEN_254;
        end
      end else begin
        Station5_7_6 <= _GEN_254;
      end
    end else begin
      Station5_7_6 <= _GEN_254;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2374 & _GEN_2277) begin // @[stationary_dpe.scala 140:32]
          Station5_7_7 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_7_7 <= _GEN_255;
        end
      end else begin
        Station5_7_7 <= _GEN_255;
      end
    end else begin
      Station5_7_7 <= _GEN_255;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2264 & _GEN_2279) begin // @[stationary_dpe.scala 152:32]
          Station6_0_0 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_0_0 <= _GEN_256;
        end
      end else begin
        Station6_0_0 <= _GEN_256;
      end
    end else begin
      Station6_0_0 <= _GEN_256;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2264 & _GEN_2265) begin // @[stationary_dpe.scala 152:32]
          Station6_0_1 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_0_1 <= _GEN_257;
        end
      end else begin
        Station6_0_1 <= _GEN_257;
      end
    end else begin
      Station6_0_1 <= _GEN_257;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2264 & _GEN_2267) begin // @[stationary_dpe.scala 152:32]
          Station6_0_2 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_0_2 <= _GEN_258;
        end
      end else begin
        Station6_0_2 <= _GEN_258;
      end
    end else begin
      Station6_0_2 <= _GEN_258;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2264 & _GEN_2269) begin // @[stationary_dpe.scala 152:32]
          Station6_0_3 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_0_3 <= _GEN_259;
        end
      end else begin
        Station6_0_3 <= _GEN_259;
      end
    end else begin
      Station6_0_3 <= _GEN_259;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2264 & _GEN_2271) begin // @[stationary_dpe.scala 152:32]
          Station6_0_4 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_0_4 <= _GEN_260;
        end
      end else begin
        Station6_0_4 <= _GEN_260;
      end
    end else begin
      Station6_0_4 <= _GEN_260;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2264 & _GEN_2273) begin // @[stationary_dpe.scala 152:32]
          Station6_0_5 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_0_5 <= _GEN_261;
        end
      end else begin
        Station6_0_5 <= _GEN_261;
      end
    end else begin
      Station6_0_5 <= _GEN_261;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2264 & _GEN_2275) begin // @[stationary_dpe.scala 152:32]
          Station6_0_6 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_0_6 <= _GEN_262;
        end
      end else begin
        Station6_0_6 <= _GEN_262;
      end
    end else begin
      Station6_0_6 <= _GEN_262;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2264 & _GEN_2277) begin // @[stationary_dpe.scala 152:32]
          Station6_0_7 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_0_7 <= _GEN_263;
        end
      end else begin
        Station6_0_7 <= _GEN_263;
      end
    end else begin
      Station6_0_7 <= _GEN_263;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2278 & _GEN_2279) begin // @[stationary_dpe.scala 152:32]
          Station6_1_0 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_1_0 <= _GEN_264;
        end
      end else begin
        Station6_1_0 <= _GEN_264;
      end
    end else begin
      Station6_1_0 <= _GEN_264;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2278 & _GEN_2265) begin // @[stationary_dpe.scala 152:32]
          Station6_1_1 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_1_1 <= _GEN_265;
        end
      end else begin
        Station6_1_1 <= _GEN_265;
      end
    end else begin
      Station6_1_1 <= _GEN_265;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2278 & _GEN_2267) begin // @[stationary_dpe.scala 152:32]
          Station6_1_2 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_1_2 <= _GEN_266;
        end
      end else begin
        Station6_1_2 <= _GEN_266;
      end
    end else begin
      Station6_1_2 <= _GEN_266;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2278 & _GEN_2269) begin // @[stationary_dpe.scala 152:32]
          Station6_1_3 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_1_3 <= _GEN_267;
        end
      end else begin
        Station6_1_3 <= _GEN_267;
      end
    end else begin
      Station6_1_3 <= _GEN_267;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2278 & _GEN_2271) begin // @[stationary_dpe.scala 152:32]
          Station6_1_4 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_1_4 <= _GEN_268;
        end
      end else begin
        Station6_1_4 <= _GEN_268;
      end
    end else begin
      Station6_1_4 <= _GEN_268;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2278 & _GEN_2273) begin // @[stationary_dpe.scala 152:32]
          Station6_1_5 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_1_5 <= _GEN_269;
        end
      end else begin
        Station6_1_5 <= _GEN_269;
      end
    end else begin
      Station6_1_5 <= _GEN_269;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2278 & _GEN_2275) begin // @[stationary_dpe.scala 152:32]
          Station6_1_6 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_1_6 <= _GEN_270;
        end
      end else begin
        Station6_1_6 <= _GEN_270;
      end
    end else begin
      Station6_1_6 <= _GEN_270;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2278 & _GEN_2277) begin // @[stationary_dpe.scala 152:32]
          Station6_1_7 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_1_7 <= _GEN_271;
        end
      end else begin
        Station6_1_7 <= _GEN_271;
      end
    end else begin
      Station6_1_7 <= _GEN_271;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2294 & _GEN_2279) begin // @[stationary_dpe.scala 152:32]
          Station6_2_0 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_2_0 <= _GEN_272;
        end
      end else begin
        Station6_2_0 <= _GEN_272;
      end
    end else begin
      Station6_2_0 <= _GEN_272;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2294 & _GEN_2265) begin // @[stationary_dpe.scala 152:32]
          Station6_2_1 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_2_1 <= _GEN_273;
        end
      end else begin
        Station6_2_1 <= _GEN_273;
      end
    end else begin
      Station6_2_1 <= _GEN_273;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2294 & _GEN_2267) begin // @[stationary_dpe.scala 152:32]
          Station6_2_2 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_2_2 <= _GEN_274;
        end
      end else begin
        Station6_2_2 <= _GEN_274;
      end
    end else begin
      Station6_2_2 <= _GEN_274;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2294 & _GEN_2269) begin // @[stationary_dpe.scala 152:32]
          Station6_2_3 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_2_3 <= _GEN_275;
        end
      end else begin
        Station6_2_3 <= _GEN_275;
      end
    end else begin
      Station6_2_3 <= _GEN_275;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2294 & _GEN_2271) begin // @[stationary_dpe.scala 152:32]
          Station6_2_4 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_2_4 <= _GEN_276;
        end
      end else begin
        Station6_2_4 <= _GEN_276;
      end
    end else begin
      Station6_2_4 <= _GEN_276;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2294 & _GEN_2273) begin // @[stationary_dpe.scala 152:32]
          Station6_2_5 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_2_5 <= _GEN_277;
        end
      end else begin
        Station6_2_5 <= _GEN_277;
      end
    end else begin
      Station6_2_5 <= _GEN_277;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2294 & _GEN_2275) begin // @[stationary_dpe.scala 152:32]
          Station6_2_6 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_2_6 <= _GEN_278;
        end
      end else begin
        Station6_2_6 <= _GEN_278;
      end
    end else begin
      Station6_2_6 <= _GEN_278;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2294 & _GEN_2277) begin // @[stationary_dpe.scala 152:32]
          Station6_2_7 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_2_7 <= _GEN_279;
        end
      end else begin
        Station6_2_7 <= _GEN_279;
      end
    end else begin
      Station6_2_7 <= _GEN_279;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2310 & _GEN_2279) begin // @[stationary_dpe.scala 152:32]
          Station6_3_0 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_3_0 <= _GEN_280;
        end
      end else begin
        Station6_3_0 <= _GEN_280;
      end
    end else begin
      Station6_3_0 <= _GEN_280;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2310 & _GEN_2265) begin // @[stationary_dpe.scala 152:32]
          Station6_3_1 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_3_1 <= _GEN_281;
        end
      end else begin
        Station6_3_1 <= _GEN_281;
      end
    end else begin
      Station6_3_1 <= _GEN_281;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2310 & _GEN_2267) begin // @[stationary_dpe.scala 152:32]
          Station6_3_2 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_3_2 <= _GEN_282;
        end
      end else begin
        Station6_3_2 <= _GEN_282;
      end
    end else begin
      Station6_3_2 <= _GEN_282;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2310 & _GEN_2269) begin // @[stationary_dpe.scala 152:32]
          Station6_3_3 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_3_3 <= _GEN_283;
        end
      end else begin
        Station6_3_3 <= _GEN_283;
      end
    end else begin
      Station6_3_3 <= _GEN_283;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2310 & _GEN_2271) begin // @[stationary_dpe.scala 152:32]
          Station6_3_4 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_3_4 <= _GEN_284;
        end
      end else begin
        Station6_3_4 <= _GEN_284;
      end
    end else begin
      Station6_3_4 <= _GEN_284;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2310 & _GEN_2273) begin // @[stationary_dpe.scala 152:32]
          Station6_3_5 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_3_5 <= _GEN_285;
        end
      end else begin
        Station6_3_5 <= _GEN_285;
      end
    end else begin
      Station6_3_5 <= _GEN_285;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2310 & _GEN_2275) begin // @[stationary_dpe.scala 152:32]
          Station6_3_6 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_3_6 <= _GEN_286;
        end
      end else begin
        Station6_3_6 <= _GEN_286;
      end
    end else begin
      Station6_3_6 <= _GEN_286;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2310 & _GEN_2277) begin // @[stationary_dpe.scala 152:32]
          Station6_3_7 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_3_7 <= _GEN_287;
        end
      end else begin
        Station6_3_7 <= _GEN_287;
      end
    end else begin
      Station6_3_7 <= _GEN_287;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2326 & _GEN_2279) begin // @[stationary_dpe.scala 152:32]
          Station6_4_0 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_4_0 <= _GEN_288;
        end
      end else begin
        Station6_4_0 <= _GEN_288;
      end
    end else begin
      Station6_4_0 <= _GEN_288;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2326 & _GEN_2265) begin // @[stationary_dpe.scala 152:32]
          Station6_4_1 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_4_1 <= _GEN_289;
        end
      end else begin
        Station6_4_1 <= _GEN_289;
      end
    end else begin
      Station6_4_1 <= _GEN_289;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2326 & _GEN_2267) begin // @[stationary_dpe.scala 152:32]
          Station6_4_2 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_4_2 <= _GEN_290;
        end
      end else begin
        Station6_4_2 <= _GEN_290;
      end
    end else begin
      Station6_4_2 <= _GEN_290;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2326 & _GEN_2269) begin // @[stationary_dpe.scala 152:32]
          Station6_4_3 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_4_3 <= _GEN_291;
        end
      end else begin
        Station6_4_3 <= _GEN_291;
      end
    end else begin
      Station6_4_3 <= _GEN_291;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2326 & _GEN_2271) begin // @[stationary_dpe.scala 152:32]
          Station6_4_4 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_4_4 <= _GEN_292;
        end
      end else begin
        Station6_4_4 <= _GEN_292;
      end
    end else begin
      Station6_4_4 <= _GEN_292;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2326 & _GEN_2273) begin // @[stationary_dpe.scala 152:32]
          Station6_4_5 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_4_5 <= _GEN_293;
        end
      end else begin
        Station6_4_5 <= _GEN_293;
      end
    end else begin
      Station6_4_5 <= _GEN_293;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2326 & _GEN_2275) begin // @[stationary_dpe.scala 152:32]
          Station6_4_6 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_4_6 <= _GEN_294;
        end
      end else begin
        Station6_4_6 <= _GEN_294;
      end
    end else begin
      Station6_4_6 <= _GEN_294;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2326 & _GEN_2277) begin // @[stationary_dpe.scala 152:32]
          Station6_4_7 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_4_7 <= _GEN_295;
        end
      end else begin
        Station6_4_7 <= _GEN_295;
      end
    end else begin
      Station6_4_7 <= _GEN_295;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2342 & _GEN_2279) begin // @[stationary_dpe.scala 152:32]
          Station6_5_0 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_5_0 <= _GEN_296;
        end
      end else begin
        Station6_5_0 <= _GEN_296;
      end
    end else begin
      Station6_5_0 <= _GEN_296;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2342 & _GEN_2265) begin // @[stationary_dpe.scala 152:32]
          Station6_5_1 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_5_1 <= _GEN_297;
        end
      end else begin
        Station6_5_1 <= _GEN_297;
      end
    end else begin
      Station6_5_1 <= _GEN_297;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2342 & _GEN_2267) begin // @[stationary_dpe.scala 152:32]
          Station6_5_2 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_5_2 <= _GEN_298;
        end
      end else begin
        Station6_5_2 <= _GEN_298;
      end
    end else begin
      Station6_5_2 <= _GEN_298;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2342 & _GEN_2269) begin // @[stationary_dpe.scala 152:32]
          Station6_5_3 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_5_3 <= _GEN_299;
        end
      end else begin
        Station6_5_3 <= _GEN_299;
      end
    end else begin
      Station6_5_3 <= _GEN_299;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2342 & _GEN_2271) begin // @[stationary_dpe.scala 152:32]
          Station6_5_4 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_5_4 <= _GEN_300;
        end
      end else begin
        Station6_5_4 <= _GEN_300;
      end
    end else begin
      Station6_5_4 <= _GEN_300;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2342 & _GEN_2273) begin // @[stationary_dpe.scala 152:32]
          Station6_5_5 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_5_5 <= _GEN_301;
        end
      end else begin
        Station6_5_5 <= _GEN_301;
      end
    end else begin
      Station6_5_5 <= _GEN_301;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2342 & _GEN_2275) begin // @[stationary_dpe.scala 152:32]
          Station6_5_6 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_5_6 <= _GEN_302;
        end
      end else begin
        Station6_5_6 <= _GEN_302;
      end
    end else begin
      Station6_5_6 <= _GEN_302;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2342 & _GEN_2277) begin // @[stationary_dpe.scala 152:32]
          Station6_5_7 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_5_7 <= _GEN_303;
        end
      end else begin
        Station6_5_7 <= _GEN_303;
      end
    end else begin
      Station6_5_7 <= _GEN_303;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2358 & _GEN_2279) begin // @[stationary_dpe.scala 152:32]
          Station6_6_0 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_6_0 <= _GEN_304;
        end
      end else begin
        Station6_6_0 <= _GEN_304;
      end
    end else begin
      Station6_6_0 <= _GEN_304;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2358 & _GEN_2265) begin // @[stationary_dpe.scala 152:32]
          Station6_6_1 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_6_1 <= _GEN_305;
        end
      end else begin
        Station6_6_1 <= _GEN_305;
      end
    end else begin
      Station6_6_1 <= _GEN_305;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2358 & _GEN_2267) begin // @[stationary_dpe.scala 152:32]
          Station6_6_2 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_6_2 <= _GEN_306;
        end
      end else begin
        Station6_6_2 <= _GEN_306;
      end
    end else begin
      Station6_6_2 <= _GEN_306;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2358 & _GEN_2269) begin // @[stationary_dpe.scala 152:32]
          Station6_6_3 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_6_3 <= _GEN_307;
        end
      end else begin
        Station6_6_3 <= _GEN_307;
      end
    end else begin
      Station6_6_3 <= _GEN_307;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2358 & _GEN_2271) begin // @[stationary_dpe.scala 152:32]
          Station6_6_4 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_6_4 <= _GEN_308;
        end
      end else begin
        Station6_6_4 <= _GEN_308;
      end
    end else begin
      Station6_6_4 <= _GEN_308;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2358 & _GEN_2273) begin // @[stationary_dpe.scala 152:32]
          Station6_6_5 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_6_5 <= _GEN_309;
        end
      end else begin
        Station6_6_5 <= _GEN_309;
      end
    end else begin
      Station6_6_5 <= _GEN_309;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2358 & _GEN_2275) begin // @[stationary_dpe.scala 152:32]
          Station6_6_6 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_6_6 <= _GEN_310;
        end
      end else begin
        Station6_6_6 <= _GEN_310;
      end
    end else begin
      Station6_6_6 <= _GEN_310;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2358 & _GEN_2277) begin // @[stationary_dpe.scala 152:32]
          Station6_6_7 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_6_7 <= _GEN_311;
        end
      end else begin
        Station6_6_7 <= _GEN_311;
      end
    end else begin
      Station6_6_7 <= _GEN_311;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2374 & _GEN_2279) begin // @[stationary_dpe.scala 152:32]
          Station6_7_0 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_7_0 <= _GEN_312;
        end
      end else begin
        Station6_7_0 <= _GEN_312;
      end
    end else begin
      Station6_7_0 <= _GEN_312;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2374 & _GEN_2265) begin // @[stationary_dpe.scala 152:32]
          Station6_7_1 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_7_1 <= _GEN_313;
        end
      end else begin
        Station6_7_1 <= _GEN_313;
      end
    end else begin
      Station6_7_1 <= _GEN_313;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2374 & _GEN_2267) begin // @[stationary_dpe.scala 152:32]
          Station6_7_2 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_7_2 <= _GEN_314;
        end
      end else begin
        Station6_7_2 <= _GEN_314;
      end
    end else begin
      Station6_7_2 <= _GEN_314;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2374 & _GEN_2269) begin // @[stationary_dpe.scala 152:32]
          Station6_7_3 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_7_3 <= _GEN_315;
        end
      end else begin
        Station6_7_3 <= _GEN_315;
      end
    end else begin
      Station6_7_3 <= _GEN_315;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2374 & _GEN_2271) begin // @[stationary_dpe.scala 152:32]
          Station6_7_4 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_7_4 <= _GEN_316;
        end
      end else begin
        Station6_7_4 <= _GEN_316;
      end
    end else begin
      Station6_7_4 <= _GEN_316;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2374 & _GEN_2273) begin // @[stationary_dpe.scala 152:32]
          Station6_7_5 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_7_5 <= _GEN_317;
        end
      end else begin
        Station6_7_5 <= _GEN_317;
      end
    end else begin
      Station6_7_5 <= _GEN_317;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2374 & _GEN_2275) begin // @[stationary_dpe.scala 152:32]
          Station6_7_6 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_7_6 <= _GEN_318;
        end
      end else begin
        Station6_7_6 <= _GEN_318;
      end
    end else begin
      Station6_7_6 <= _GEN_318;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2374 & _GEN_2277) begin // @[stationary_dpe.scala 152:32]
          Station6_7_7 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_7_7 <= _GEN_319;
        end
      end else begin
        Station6_7_7 <= _GEN_319;
      end
    end else begin
      Station6_7_7 <= _GEN_319;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2264 & _GEN_2279) begin // @[stationary_dpe.scala 164:32]
          Station7_0_0 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_0_0 <= _GEN_320;
        end
      end else begin
        Station7_0_0 <= _GEN_320;
      end
    end else begin
      Station7_0_0 <= _GEN_320;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2264 & _GEN_2265) begin // @[stationary_dpe.scala 164:32]
          Station7_0_1 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_0_1 <= _GEN_321;
        end
      end else begin
        Station7_0_1 <= _GEN_321;
      end
    end else begin
      Station7_0_1 <= _GEN_321;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2264 & _GEN_2267) begin // @[stationary_dpe.scala 164:32]
          Station7_0_2 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_0_2 <= _GEN_322;
        end
      end else begin
        Station7_0_2 <= _GEN_322;
      end
    end else begin
      Station7_0_2 <= _GEN_322;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2264 & _GEN_2269) begin // @[stationary_dpe.scala 164:32]
          Station7_0_3 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_0_3 <= _GEN_323;
        end
      end else begin
        Station7_0_3 <= _GEN_323;
      end
    end else begin
      Station7_0_3 <= _GEN_323;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2264 & _GEN_2271) begin // @[stationary_dpe.scala 164:32]
          Station7_0_4 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_0_4 <= _GEN_324;
        end
      end else begin
        Station7_0_4 <= _GEN_324;
      end
    end else begin
      Station7_0_4 <= _GEN_324;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2264 & _GEN_2273) begin // @[stationary_dpe.scala 164:32]
          Station7_0_5 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_0_5 <= _GEN_325;
        end
      end else begin
        Station7_0_5 <= _GEN_325;
      end
    end else begin
      Station7_0_5 <= _GEN_325;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2264 & _GEN_2275) begin // @[stationary_dpe.scala 164:32]
          Station7_0_6 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_0_6 <= _GEN_326;
        end
      end else begin
        Station7_0_6 <= _GEN_326;
      end
    end else begin
      Station7_0_6 <= _GEN_326;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2264 & _GEN_2277) begin // @[stationary_dpe.scala 164:32]
          Station7_0_7 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_0_7 <= _GEN_327;
        end
      end else begin
        Station7_0_7 <= _GEN_327;
      end
    end else begin
      Station7_0_7 <= _GEN_327;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2278 & _GEN_2279) begin // @[stationary_dpe.scala 164:32]
          Station7_1_0 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_1_0 <= _GEN_328;
        end
      end else begin
        Station7_1_0 <= _GEN_328;
      end
    end else begin
      Station7_1_0 <= _GEN_328;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2278 & _GEN_2265) begin // @[stationary_dpe.scala 164:32]
          Station7_1_1 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_1_1 <= _GEN_329;
        end
      end else begin
        Station7_1_1 <= _GEN_329;
      end
    end else begin
      Station7_1_1 <= _GEN_329;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2278 & _GEN_2267) begin // @[stationary_dpe.scala 164:32]
          Station7_1_2 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_1_2 <= _GEN_330;
        end
      end else begin
        Station7_1_2 <= _GEN_330;
      end
    end else begin
      Station7_1_2 <= _GEN_330;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2278 & _GEN_2269) begin // @[stationary_dpe.scala 164:32]
          Station7_1_3 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_1_3 <= _GEN_331;
        end
      end else begin
        Station7_1_3 <= _GEN_331;
      end
    end else begin
      Station7_1_3 <= _GEN_331;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2278 & _GEN_2271) begin // @[stationary_dpe.scala 164:32]
          Station7_1_4 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_1_4 <= _GEN_332;
        end
      end else begin
        Station7_1_4 <= _GEN_332;
      end
    end else begin
      Station7_1_4 <= _GEN_332;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2278 & _GEN_2273) begin // @[stationary_dpe.scala 164:32]
          Station7_1_5 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_1_5 <= _GEN_333;
        end
      end else begin
        Station7_1_5 <= _GEN_333;
      end
    end else begin
      Station7_1_5 <= _GEN_333;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2278 & _GEN_2275) begin // @[stationary_dpe.scala 164:32]
          Station7_1_6 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_1_6 <= _GEN_334;
        end
      end else begin
        Station7_1_6 <= _GEN_334;
      end
    end else begin
      Station7_1_6 <= _GEN_334;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2278 & _GEN_2277) begin // @[stationary_dpe.scala 164:32]
          Station7_1_7 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_1_7 <= _GEN_335;
        end
      end else begin
        Station7_1_7 <= _GEN_335;
      end
    end else begin
      Station7_1_7 <= _GEN_335;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2294 & _GEN_2279) begin // @[stationary_dpe.scala 164:32]
          Station7_2_0 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_2_0 <= _GEN_336;
        end
      end else begin
        Station7_2_0 <= _GEN_336;
      end
    end else begin
      Station7_2_0 <= _GEN_336;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2294 & _GEN_2265) begin // @[stationary_dpe.scala 164:32]
          Station7_2_1 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_2_1 <= _GEN_337;
        end
      end else begin
        Station7_2_1 <= _GEN_337;
      end
    end else begin
      Station7_2_1 <= _GEN_337;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2294 & _GEN_2267) begin // @[stationary_dpe.scala 164:32]
          Station7_2_2 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_2_2 <= _GEN_338;
        end
      end else begin
        Station7_2_2 <= _GEN_338;
      end
    end else begin
      Station7_2_2 <= _GEN_338;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2294 & _GEN_2269) begin // @[stationary_dpe.scala 164:32]
          Station7_2_3 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_2_3 <= _GEN_339;
        end
      end else begin
        Station7_2_3 <= _GEN_339;
      end
    end else begin
      Station7_2_3 <= _GEN_339;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2294 & _GEN_2271) begin // @[stationary_dpe.scala 164:32]
          Station7_2_4 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_2_4 <= _GEN_340;
        end
      end else begin
        Station7_2_4 <= _GEN_340;
      end
    end else begin
      Station7_2_4 <= _GEN_340;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2294 & _GEN_2273) begin // @[stationary_dpe.scala 164:32]
          Station7_2_5 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_2_5 <= _GEN_341;
        end
      end else begin
        Station7_2_5 <= _GEN_341;
      end
    end else begin
      Station7_2_5 <= _GEN_341;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2294 & _GEN_2275) begin // @[stationary_dpe.scala 164:32]
          Station7_2_6 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_2_6 <= _GEN_342;
        end
      end else begin
        Station7_2_6 <= _GEN_342;
      end
    end else begin
      Station7_2_6 <= _GEN_342;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2294 & _GEN_2277) begin // @[stationary_dpe.scala 164:32]
          Station7_2_7 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_2_7 <= _GEN_343;
        end
      end else begin
        Station7_2_7 <= _GEN_343;
      end
    end else begin
      Station7_2_7 <= _GEN_343;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2310 & _GEN_2279) begin // @[stationary_dpe.scala 164:32]
          Station7_3_0 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_3_0 <= _GEN_344;
        end
      end else begin
        Station7_3_0 <= _GEN_344;
      end
    end else begin
      Station7_3_0 <= _GEN_344;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2310 & _GEN_2265) begin // @[stationary_dpe.scala 164:32]
          Station7_3_1 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_3_1 <= _GEN_345;
        end
      end else begin
        Station7_3_1 <= _GEN_345;
      end
    end else begin
      Station7_3_1 <= _GEN_345;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2310 & _GEN_2267) begin // @[stationary_dpe.scala 164:32]
          Station7_3_2 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_3_2 <= _GEN_346;
        end
      end else begin
        Station7_3_2 <= _GEN_346;
      end
    end else begin
      Station7_3_2 <= _GEN_346;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2310 & _GEN_2269) begin // @[stationary_dpe.scala 164:32]
          Station7_3_3 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_3_3 <= _GEN_347;
        end
      end else begin
        Station7_3_3 <= _GEN_347;
      end
    end else begin
      Station7_3_3 <= _GEN_347;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2310 & _GEN_2271) begin // @[stationary_dpe.scala 164:32]
          Station7_3_4 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_3_4 <= _GEN_348;
        end
      end else begin
        Station7_3_4 <= _GEN_348;
      end
    end else begin
      Station7_3_4 <= _GEN_348;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2310 & _GEN_2273) begin // @[stationary_dpe.scala 164:32]
          Station7_3_5 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_3_5 <= _GEN_349;
        end
      end else begin
        Station7_3_5 <= _GEN_349;
      end
    end else begin
      Station7_3_5 <= _GEN_349;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2310 & _GEN_2275) begin // @[stationary_dpe.scala 164:32]
          Station7_3_6 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_3_6 <= _GEN_350;
        end
      end else begin
        Station7_3_6 <= _GEN_350;
      end
    end else begin
      Station7_3_6 <= _GEN_350;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2310 & _GEN_2277) begin // @[stationary_dpe.scala 164:32]
          Station7_3_7 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_3_7 <= _GEN_351;
        end
      end else begin
        Station7_3_7 <= _GEN_351;
      end
    end else begin
      Station7_3_7 <= _GEN_351;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2326 & _GEN_2279) begin // @[stationary_dpe.scala 164:32]
          Station7_4_0 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_4_0 <= _GEN_352;
        end
      end else begin
        Station7_4_0 <= _GEN_352;
      end
    end else begin
      Station7_4_0 <= _GEN_352;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2326 & _GEN_2265) begin // @[stationary_dpe.scala 164:32]
          Station7_4_1 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_4_1 <= _GEN_353;
        end
      end else begin
        Station7_4_1 <= _GEN_353;
      end
    end else begin
      Station7_4_1 <= _GEN_353;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2326 & _GEN_2267) begin // @[stationary_dpe.scala 164:32]
          Station7_4_2 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_4_2 <= _GEN_354;
        end
      end else begin
        Station7_4_2 <= _GEN_354;
      end
    end else begin
      Station7_4_2 <= _GEN_354;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2326 & _GEN_2269) begin // @[stationary_dpe.scala 164:32]
          Station7_4_3 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_4_3 <= _GEN_355;
        end
      end else begin
        Station7_4_3 <= _GEN_355;
      end
    end else begin
      Station7_4_3 <= _GEN_355;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2326 & _GEN_2271) begin // @[stationary_dpe.scala 164:32]
          Station7_4_4 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_4_4 <= _GEN_356;
        end
      end else begin
        Station7_4_4 <= _GEN_356;
      end
    end else begin
      Station7_4_4 <= _GEN_356;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2326 & _GEN_2273) begin // @[stationary_dpe.scala 164:32]
          Station7_4_5 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_4_5 <= _GEN_357;
        end
      end else begin
        Station7_4_5 <= _GEN_357;
      end
    end else begin
      Station7_4_5 <= _GEN_357;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2326 & _GEN_2275) begin // @[stationary_dpe.scala 164:32]
          Station7_4_6 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_4_6 <= _GEN_358;
        end
      end else begin
        Station7_4_6 <= _GEN_358;
      end
    end else begin
      Station7_4_6 <= _GEN_358;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2326 & _GEN_2277) begin // @[stationary_dpe.scala 164:32]
          Station7_4_7 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_4_7 <= _GEN_359;
        end
      end else begin
        Station7_4_7 <= _GEN_359;
      end
    end else begin
      Station7_4_7 <= _GEN_359;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2342 & _GEN_2279) begin // @[stationary_dpe.scala 164:32]
          Station7_5_0 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_5_0 <= _GEN_360;
        end
      end else begin
        Station7_5_0 <= _GEN_360;
      end
    end else begin
      Station7_5_0 <= _GEN_360;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2342 & _GEN_2265) begin // @[stationary_dpe.scala 164:32]
          Station7_5_1 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_5_1 <= _GEN_361;
        end
      end else begin
        Station7_5_1 <= _GEN_361;
      end
    end else begin
      Station7_5_1 <= _GEN_361;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2342 & _GEN_2267) begin // @[stationary_dpe.scala 164:32]
          Station7_5_2 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_5_2 <= _GEN_362;
        end
      end else begin
        Station7_5_2 <= _GEN_362;
      end
    end else begin
      Station7_5_2 <= _GEN_362;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2342 & _GEN_2269) begin // @[stationary_dpe.scala 164:32]
          Station7_5_3 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_5_3 <= _GEN_363;
        end
      end else begin
        Station7_5_3 <= _GEN_363;
      end
    end else begin
      Station7_5_3 <= _GEN_363;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2342 & _GEN_2271) begin // @[stationary_dpe.scala 164:32]
          Station7_5_4 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_5_4 <= _GEN_364;
        end
      end else begin
        Station7_5_4 <= _GEN_364;
      end
    end else begin
      Station7_5_4 <= _GEN_364;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2342 & _GEN_2273) begin // @[stationary_dpe.scala 164:32]
          Station7_5_5 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_5_5 <= _GEN_365;
        end
      end else begin
        Station7_5_5 <= _GEN_365;
      end
    end else begin
      Station7_5_5 <= _GEN_365;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2342 & _GEN_2275) begin // @[stationary_dpe.scala 164:32]
          Station7_5_6 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_5_6 <= _GEN_366;
        end
      end else begin
        Station7_5_6 <= _GEN_366;
      end
    end else begin
      Station7_5_6 <= _GEN_366;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2342 & _GEN_2277) begin // @[stationary_dpe.scala 164:32]
          Station7_5_7 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_5_7 <= _GEN_367;
        end
      end else begin
        Station7_5_7 <= _GEN_367;
      end
    end else begin
      Station7_5_7 <= _GEN_367;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2358 & _GEN_2279) begin // @[stationary_dpe.scala 164:32]
          Station7_6_0 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_6_0 <= _GEN_368;
        end
      end else begin
        Station7_6_0 <= _GEN_368;
      end
    end else begin
      Station7_6_0 <= _GEN_368;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2358 & _GEN_2265) begin // @[stationary_dpe.scala 164:32]
          Station7_6_1 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_6_1 <= _GEN_369;
        end
      end else begin
        Station7_6_1 <= _GEN_369;
      end
    end else begin
      Station7_6_1 <= _GEN_369;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2358 & _GEN_2267) begin // @[stationary_dpe.scala 164:32]
          Station7_6_2 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_6_2 <= _GEN_370;
        end
      end else begin
        Station7_6_2 <= _GEN_370;
      end
    end else begin
      Station7_6_2 <= _GEN_370;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2358 & _GEN_2269) begin // @[stationary_dpe.scala 164:32]
          Station7_6_3 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_6_3 <= _GEN_371;
        end
      end else begin
        Station7_6_3 <= _GEN_371;
      end
    end else begin
      Station7_6_3 <= _GEN_371;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2358 & _GEN_2271) begin // @[stationary_dpe.scala 164:32]
          Station7_6_4 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_6_4 <= _GEN_372;
        end
      end else begin
        Station7_6_4 <= _GEN_372;
      end
    end else begin
      Station7_6_4 <= _GEN_372;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2358 & _GEN_2273) begin // @[stationary_dpe.scala 164:32]
          Station7_6_5 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_6_5 <= _GEN_373;
        end
      end else begin
        Station7_6_5 <= _GEN_373;
      end
    end else begin
      Station7_6_5 <= _GEN_373;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2358 & _GEN_2275) begin // @[stationary_dpe.scala 164:32]
          Station7_6_6 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_6_6 <= _GEN_374;
        end
      end else begin
        Station7_6_6 <= _GEN_374;
      end
    end else begin
      Station7_6_6 <= _GEN_374;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2358 & _GEN_2277) begin // @[stationary_dpe.scala 164:32]
          Station7_6_7 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_6_7 <= _GEN_375;
        end
      end else begin
        Station7_6_7 <= _GEN_375;
      end
    end else begin
      Station7_6_7 <= _GEN_375;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2374 & _GEN_2279) begin // @[stationary_dpe.scala 164:32]
          Station7_7_0 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_7_0 <= _GEN_376;
        end
      end else begin
        Station7_7_0 <= _GEN_376;
      end
    end else begin
      Station7_7_0 <= _GEN_376;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2374 & _GEN_2265) begin // @[stationary_dpe.scala 164:32]
          Station7_7_1 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_7_1 <= _GEN_377;
        end
      end else begin
        Station7_7_1 <= _GEN_377;
      end
    end else begin
      Station7_7_1 <= _GEN_377;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2374 & _GEN_2267) begin // @[stationary_dpe.scala 164:32]
          Station7_7_2 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_7_2 <= _GEN_378;
        end
      end else begin
        Station7_7_2 <= _GEN_378;
      end
    end else begin
      Station7_7_2 <= _GEN_378;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2374 & _GEN_2269) begin // @[stationary_dpe.scala 164:32]
          Station7_7_3 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_7_3 <= _GEN_379;
        end
      end else begin
        Station7_7_3 <= _GEN_379;
      end
    end else begin
      Station7_7_3 <= _GEN_379;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2374 & _GEN_2271) begin // @[stationary_dpe.scala 164:32]
          Station7_7_4 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_7_4 <= _GEN_380;
        end
      end else begin
        Station7_7_4 <= _GEN_380;
      end
    end else begin
      Station7_7_4 <= _GEN_380;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2374 & _GEN_2273) begin // @[stationary_dpe.scala 164:32]
          Station7_7_5 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_7_5 <= _GEN_381;
        end
      end else begin
        Station7_7_5 <= _GEN_381;
      end
    end else begin
      Station7_7_5 <= _GEN_381;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2374 & _GEN_2275) begin // @[stationary_dpe.scala 164:32]
          Station7_7_6 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_7_6 <= _GEN_382;
        end
      end else begin
        Station7_7_6 <= _GEN_382;
      end
    end else begin
      Station7_7_6 <= _GEN_382;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2374 & _GEN_2277) begin // @[stationary_dpe.scala 164:32]
          Station7_7_7 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_7_7 <= _GEN_383;
        end
      end else begin
        Station7_7_7 <= _GEN_383;
      end
    end else begin
      Station7_7_7 <= _GEN_383;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2264 & _GEN_2279) begin // @[stationary_dpe.scala 176:32]
          Station8_0_0 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_0_0 <= _GEN_384;
        end
      end else begin
        Station8_0_0 <= _GEN_384;
      end
    end else begin
      Station8_0_0 <= _GEN_384;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2264 & _GEN_2265) begin // @[stationary_dpe.scala 176:32]
          Station8_0_1 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_0_1 <= _GEN_385;
        end
      end else begin
        Station8_0_1 <= _GEN_385;
      end
    end else begin
      Station8_0_1 <= _GEN_385;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2264 & _GEN_2267) begin // @[stationary_dpe.scala 176:32]
          Station8_0_2 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_0_2 <= _GEN_386;
        end
      end else begin
        Station8_0_2 <= _GEN_386;
      end
    end else begin
      Station8_0_2 <= _GEN_386;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2264 & _GEN_2269) begin // @[stationary_dpe.scala 176:32]
          Station8_0_3 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_0_3 <= _GEN_387;
        end
      end else begin
        Station8_0_3 <= _GEN_387;
      end
    end else begin
      Station8_0_3 <= _GEN_387;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2264 & _GEN_2271) begin // @[stationary_dpe.scala 176:32]
          Station8_0_4 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_0_4 <= _GEN_388;
        end
      end else begin
        Station8_0_4 <= _GEN_388;
      end
    end else begin
      Station8_0_4 <= _GEN_388;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2264 & _GEN_2273) begin // @[stationary_dpe.scala 176:32]
          Station8_0_5 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_0_5 <= _GEN_389;
        end
      end else begin
        Station8_0_5 <= _GEN_389;
      end
    end else begin
      Station8_0_5 <= _GEN_389;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2264 & _GEN_2275) begin // @[stationary_dpe.scala 176:32]
          Station8_0_6 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_0_6 <= _GEN_390;
        end
      end else begin
        Station8_0_6 <= _GEN_390;
      end
    end else begin
      Station8_0_6 <= _GEN_390;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2264 & _GEN_2277) begin // @[stationary_dpe.scala 176:32]
          Station8_0_7 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_0_7 <= _GEN_391;
        end
      end else begin
        Station8_0_7 <= _GEN_391;
      end
    end else begin
      Station8_0_7 <= _GEN_391;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2278 & _GEN_2279) begin // @[stationary_dpe.scala 176:32]
          Station8_1_0 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_1_0 <= _GEN_392;
        end
      end else begin
        Station8_1_0 <= _GEN_392;
      end
    end else begin
      Station8_1_0 <= _GEN_392;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2278 & _GEN_2265) begin // @[stationary_dpe.scala 176:32]
          Station8_1_1 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_1_1 <= _GEN_393;
        end
      end else begin
        Station8_1_1 <= _GEN_393;
      end
    end else begin
      Station8_1_1 <= _GEN_393;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2278 & _GEN_2267) begin // @[stationary_dpe.scala 176:32]
          Station8_1_2 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_1_2 <= _GEN_394;
        end
      end else begin
        Station8_1_2 <= _GEN_394;
      end
    end else begin
      Station8_1_2 <= _GEN_394;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2278 & _GEN_2269) begin // @[stationary_dpe.scala 176:32]
          Station8_1_3 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_1_3 <= _GEN_395;
        end
      end else begin
        Station8_1_3 <= _GEN_395;
      end
    end else begin
      Station8_1_3 <= _GEN_395;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2278 & _GEN_2271) begin // @[stationary_dpe.scala 176:32]
          Station8_1_4 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_1_4 <= _GEN_396;
        end
      end else begin
        Station8_1_4 <= _GEN_396;
      end
    end else begin
      Station8_1_4 <= _GEN_396;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2278 & _GEN_2273) begin // @[stationary_dpe.scala 176:32]
          Station8_1_5 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_1_5 <= _GEN_397;
        end
      end else begin
        Station8_1_5 <= _GEN_397;
      end
    end else begin
      Station8_1_5 <= _GEN_397;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2278 & _GEN_2275) begin // @[stationary_dpe.scala 176:32]
          Station8_1_6 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_1_6 <= _GEN_398;
        end
      end else begin
        Station8_1_6 <= _GEN_398;
      end
    end else begin
      Station8_1_6 <= _GEN_398;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2278 & _GEN_2277) begin // @[stationary_dpe.scala 176:32]
          Station8_1_7 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_1_7 <= _GEN_399;
        end
      end else begin
        Station8_1_7 <= _GEN_399;
      end
    end else begin
      Station8_1_7 <= _GEN_399;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2294 & _GEN_2279) begin // @[stationary_dpe.scala 176:32]
          Station8_2_0 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_2_0 <= _GEN_400;
        end
      end else begin
        Station8_2_0 <= _GEN_400;
      end
    end else begin
      Station8_2_0 <= _GEN_400;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2294 & _GEN_2265) begin // @[stationary_dpe.scala 176:32]
          Station8_2_1 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_2_1 <= _GEN_401;
        end
      end else begin
        Station8_2_1 <= _GEN_401;
      end
    end else begin
      Station8_2_1 <= _GEN_401;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2294 & _GEN_2267) begin // @[stationary_dpe.scala 176:32]
          Station8_2_2 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_2_2 <= _GEN_402;
        end
      end else begin
        Station8_2_2 <= _GEN_402;
      end
    end else begin
      Station8_2_2 <= _GEN_402;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2294 & _GEN_2269) begin // @[stationary_dpe.scala 176:32]
          Station8_2_3 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_2_3 <= _GEN_403;
        end
      end else begin
        Station8_2_3 <= _GEN_403;
      end
    end else begin
      Station8_2_3 <= _GEN_403;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2294 & _GEN_2271) begin // @[stationary_dpe.scala 176:32]
          Station8_2_4 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_2_4 <= _GEN_404;
        end
      end else begin
        Station8_2_4 <= _GEN_404;
      end
    end else begin
      Station8_2_4 <= _GEN_404;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2294 & _GEN_2273) begin // @[stationary_dpe.scala 176:32]
          Station8_2_5 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_2_5 <= _GEN_405;
        end
      end else begin
        Station8_2_5 <= _GEN_405;
      end
    end else begin
      Station8_2_5 <= _GEN_405;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2294 & _GEN_2275) begin // @[stationary_dpe.scala 176:32]
          Station8_2_6 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_2_6 <= _GEN_406;
        end
      end else begin
        Station8_2_6 <= _GEN_406;
      end
    end else begin
      Station8_2_6 <= _GEN_406;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2294 & _GEN_2277) begin // @[stationary_dpe.scala 176:32]
          Station8_2_7 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_2_7 <= _GEN_407;
        end
      end else begin
        Station8_2_7 <= _GEN_407;
      end
    end else begin
      Station8_2_7 <= _GEN_407;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2310 & _GEN_2279) begin // @[stationary_dpe.scala 176:32]
          Station8_3_0 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_3_0 <= _GEN_408;
        end
      end else begin
        Station8_3_0 <= _GEN_408;
      end
    end else begin
      Station8_3_0 <= _GEN_408;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2310 & _GEN_2265) begin // @[stationary_dpe.scala 176:32]
          Station8_3_1 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_3_1 <= _GEN_409;
        end
      end else begin
        Station8_3_1 <= _GEN_409;
      end
    end else begin
      Station8_3_1 <= _GEN_409;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2310 & _GEN_2267) begin // @[stationary_dpe.scala 176:32]
          Station8_3_2 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_3_2 <= _GEN_410;
        end
      end else begin
        Station8_3_2 <= _GEN_410;
      end
    end else begin
      Station8_3_2 <= _GEN_410;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2310 & _GEN_2269) begin // @[stationary_dpe.scala 176:32]
          Station8_3_3 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_3_3 <= _GEN_411;
        end
      end else begin
        Station8_3_3 <= _GEN_411;
      end
    end else begin
      Station8_3_3 <= _GEN_411;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2310 & _GEN_2271) begin // @[stationary_dpe.scala 176:32]
          Station8_3_4 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_3_4 <= _GEN_412;
        end
      end else begin
        Station8_3_4 <= _GEN_412;
      end
    end else begin
      Station8_3_4 <= _GEN_412;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2310 & _GEN_2273) begin // @[stationary_dpe.scala 176:32]
          Station8_3_5 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_3_5 <= _GEN_413;
        end
      end else begin
        Station8_3_5 <= _GEN_413;
      end
    end else begin
      Station8_3_5 <= _GEN_413;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2310 & _GEN_2275) begin // @[stationary_dpe.scala 176:32]
          Station8_3_6 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_3_6 <= _GEN_414;
        end
      end else begin
        Station8_3_6 <= _GEN_414;
      end
    end else begin
      Station8_3_6 <= _GEN_414;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2310 & _GEN_2277) begin // @[stationary_dpe.scala 176:32]
          Station8_3_7 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_3_7 <= _GEN_415;
        end
      end else begin
        Station8_3_7 <= _GEN_415;
      end
    end else begin
      Station8_3_7 <= _GEN_415;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2326 & _GEN_2279) begin // @[stationary_dpe.scala 176:32]
          Station8_4_0 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_4_0 <= _GEN_416;
        end
      end else begin
        Station8_4_0 <= _GEN_416;
      end
    end else begin
      Station8_4_0 <= _GEN_416;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2326 & _GEN_2265) begin // @[stationary_dpe.scala 176:32]
          Station8_4_1 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_4_1 <= _GEN_417;
        end
      end else begin
        Station8_4_1 <= _GEN_417;
      end
    end else begin
      Station8_4_1 <= _GEN_417;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2326 & _GEN_2267) begin // @[stationary_dpe.scala 176:32]
          Station8_4_2 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_4_2 <= _GEN_418;
        end
      end else begin
        Station8_4_2 <= _GEN_418;
      end
    end else begin
      Station8_4_2 <= _GEN_418;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2326 & _GEN_2269) begin // @[stationary_dpe.scala 176:32]
          Station8_4_3 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_4_3 <= _GEN_419;
        end
      end else begin
        Station8_4_3 <= _GEN_419;
      end
    end else begin
      Station8_4_3 <= _GEN_419;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2326 & _GEN_2271) begin // @[stationary_dpe.scala 176:32]
          Station8_4_4 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_4_4 <= _GEN_420;
        end
      end else begin
        Station8_4_4 <= _GEN_420;
      end
    end else begin
      Station8_4_4 <= _GEN_420;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2326 & _GEN_2273) begin // @[stationary_dpe.scala 176:32]
          Station8_4_5 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_4_5 <= _GEN_421;
        end
      end else begin
        Station8_4_5 <= _GEN_421;
      end
    end else begin
      Station8_4_5 <= _GEN_421;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2326 & _GEN_2275) begin // @[stationary_dpe.scala 176:32]
          Station8_4_6 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_4_6 <= _GEN_422;
        end
      end else begin
        Station8_4_6 <= _GEN_422;
      end
    end else begin
      Station8_4_6 <= _GEN_422;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2326 & _GEN_2277) begin // @[stationary_dpe.scala 176:32]
          Station8_4_7 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_4_7 <= _GEN_423;
        end
      end else begin
        Station8_4_7 <= _GEN_423;
      end
    end else begin
      Station8_4_7 <= _GEN_423;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2342 & _GEN_2279) begin // @[stationary_dpe.scala 176:32]
          Station8_5_0 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_5_0 <= _GEN_424;
        end
      end else begin
        Station8_5_0 <= _GEN_424;
      end
    end else begin
      Station8_5_0 <= _GEN_424;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2342 & _GEN_2265) begin // @[stationary_dpe.scala 176:32]
          Station8_5_1 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_5_1 <= _GEN_425;
        end
      end else begin
        Station8_5_1 <= _GEN_425;
      end
    end else begin
      Station8_5_1 <= _GEN_425;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2342 & _GEN_2267) begin // @[stationary_dpe.scala 176:32]
          Station8_5_2 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_5_2 <= _GEN_426;
        end
      end else begin
        Station8_5_2 <= _GEN_426;
      end
    end else begin
      Station8_5_2 <= _GEN_426;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2342 & _GEN_2269) begin // @[stationary_dpe.scala 176:32]
          Station8_5_3 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_5_3 <= _GEN_427;
        end
      end else begin
        Station8_5_3 <= _GEN_427;
      end
    end else begin
      Station8_5_3 <= _GEN_427;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2342 & _GEN_2271) begin // @[stationary_dpe.scala 176:32]
          Station8_5_4 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_5_4 <= _GEN_428;
        end
      end else begin
        Station8_5_4 <= _GEN_428;
      end
    end else begin
      Station8_5_4 <= _GEN_428;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2342 & _GEN_2273) begin // @[stationary_dpe.scala 176:32]
          Station8_5_5 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_5_5 <= _GEN_429;
        end
      end else begin
        Station8_5_5 <= _GEN_429;
      end
    end else begin
      Station8_5_5 <= _GEN_429;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2342 & _GEN_2275) begin // @[stationary_dpe.scala 176:32]
          Station8_5_6 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_5_6 <= _GEN_430;
        end
      end else begin
        Station8_5_6 <= _GEN_430;
      end
    end else begin
      Station8_5_6 <= _GEN_430;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2342 & _GEN_2277) begin // @[stationary_dpe.scala 176:32]
          Station8_5_7 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_5_7 <= _GEN_431;
        end
      end else begin
        Station8_5_7 <= _GEN_431;
      end
    end else begin
      Station8_5_7 <= _GEN_431;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2358 & _GEN_2279) begin // @[stationary_dpe.scala 176:32]
          Station8_6_0 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_6_0 <= _GEN_432;
        end
      end else begin
        Station8_6_0 <= _GEN_432;
      end
    end else begin
      Station8_6_0 <= _GEN_432;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2358 & _GEN_2265) begin // @[stationary_dpe.scala 176:32]
          Station8_6_1 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_6_1 <= _GEN_433;
        end
      end else begin
        Station8_6_1 <= _GEN_433;
      end
    end else begin
      Station8_6_1 <= _GEN_433;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2358 & _GEN_2267) begin // @[stationary_dpe.scala 176:32]
          Station8_6_2 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_6_2 <= _GEN_434;
        end
      end else begin
        Station8_6_2 <= _GEN_434;
      end
    end else begin
      Station8_6_2 <= _GEN_434;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2358 & _GEN_2269) begin // @[stationary_dpe.scala 176:32]
          Station8_6_3 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_6_3 <= _GEN_435;
        end
      end else begin
        Station8_6_3 <= _GEN_435;
      end
    end else begin
      Station8_6_3 <= _GEN_435;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2358 & _GEN_2271) begin // @[stationary_dpe.scala 176:32]
          Station8_6_4 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_6_4 <= _GEN_436;
        end
      end else begin
        Station8_6_4 <= _GEN_436;
      end
    end else begin
      Station8_6_4 <= _GEN_436;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2358 & _GEN_2273) begin // @[stationary_dpe.scala 176:32]
          Station8_6_5 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_6_5 <= _GEN_437;
        end
      end else begin
        Station8_6_5 <= _GEN_437;
      end
    end else begin
      Station8_6_5 <= _GEN_437;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2358 & _GEN_2275) begin // @[stationary_dpe.scala 176:32]
          Station8_6_6 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_6_6 <= _GEN_438;
        end
      end else begin
        Station8_6_6 <= _GEN_438;
      end
    end else begin
      Station8_6_6 <= _GEN_438;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2358 & _GEN_2277) begin // @[stationary_dpe.scala 176:32]
          Station8_6_7 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_6_7 <= _GEN_439;
        end
      end else begin
        Station8_6_7 <= _GEN_439;
      end
    end else begin
      Station8_6_7 <= _GEN_439;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2374 & _GEN_2279) begin // @[stationary_dpe.scala 176:32]
          Station8_7_0 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_7_0 <= _GEN_440;
        end
      end else begin
        Station8_7_0 <= _GEN_440;
      end
    end else begin
      Station8_7_0 <= _GEN_440;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2374 & _GEN_2265) begin // @[stationary_dpe.scala 176:32]
          Station8_7_1 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_7_1 <= _GEN_441;
        end
      end else begin
        Station8_7_1 <= _GEN_441;
      end
    end else begin
      Station8_7_1 <= _GEN_441;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2374 & _GEN_2267) begin // @[stationary_dpe.scala 176:32]
          Station8_7_2 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_7_2 <= _GEN_442;
        end
      end else begin
        Station8_7_2 <= _GEN_442;
      end
    end else begin
      Station8_7_2 <= _GEN_442;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2374 & _GEN_2269) begin // @[stationary_dpe.scala 176:32]
          Station8_7_3 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_7_3 <= _GEN_443;
        end
      end else begin
        Station8_7_3 <= _GEN_443;
      end
    end else begin
      Station8_7_3 <= _GEN_443;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2374 & _GEN_2271) begin // @[stationary_dpe.scala 176:32]
          Station8_7_4 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_7_4 <= _GEN_444;
        end
      end else begin
        Station8_7_4 <= _GEN_444;
      end
    end else begin
      Station8_7_4 <= _GEN_444;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2374 & _GEN_2273) begin // @[stationary_dpe.scala 176:32]
          Station8_7_5 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_7_5 <= _GEN_445;
        end
      end else begin
        Station8_7_5 <= _GEN_445;
      end
    end else begin
      Station8_7_5 <= _GEN_445;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2374 & _GEN_2275) begin // @[stationary_dpe.scala 176:32]
          Station8_7_6 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_7_6 <= _GEN_446;
        end
      end else begin
        Station8_7_6 <= _GEN_446;
      end
    end else begin
      Station8_7_6 <= _GEN_446;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2374 & _GEN_2277) begin // @[stationary_dpe.scala 176:32]
          Station8_7_7 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_7_7 <= _GEN_447;
        end
      end else begin
        Station8_7_7 <= _GEN_447;
      end
    end else begin
      Station8_7_7 <= _GEN_447;
    end
    if (reset) begin // @[stationary_dpe.scala 79:20]
      i <= 32'h0; // @[stationary_dpe.scala 79:20]
    end else if (i < 32'h7 & j == 32'h7) begin // @[stationary_dpe.scala 222:74]
      i <= _i_T_1; // @[stationary_dpe.scala 223:11]
    end
    if (reset) begin // @[stationary_dpe.scala 80:20]
      j <= 32'h0; // @[stationary_dpe.scala 80:20]
    end else if (j < 32'h7 & i <= 32'h7) begin // @[stationary_dpe.scala 226:71]
      j <= _j_T_1; // @[stationary_dpe.scala 227:11]
    end else if (!(i == 32'h7 & _T_57)) begin // @[stationary_dpe.scala 229:81]
      j <= 32'h0; // @[stationary_dpe.scala 233:11]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  Station2_0_0 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  Station2_0_1 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  Station2_0_2 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  Station2_0_3 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  Station2_0_4 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  Station2_0_5 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  Station2_0_6 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  Station2_0_7 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  Station2_1_0 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  Station2_1_1 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  Station2_1_2 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  Station2_1_3 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  Station2_1_4 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  Station2_1_5 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  Station2_1_6 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  Station2_1_7 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  Station2_2_0 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  Station2_2_1 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  Station2_2_2 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  Station2_2_3 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  Station2_2_4 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  Station2_2_5 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  Station2_2_6 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  Station2_2_7 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  Station2_3_0 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  Station2_3_1 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  Station2_3_2 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  Station2_3_3 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  Station2_3_4 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  Station2_3_5 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  Station2_3_6 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  Station2_3_7 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  Station2_4_0 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  Station2_4_1 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  Station2_4_2 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  Station2_4_3 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  Station2_4_4 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  Station2_4_5 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  Station2_4_6 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  Station2_4_7 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  Station2_5_0 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  Station2_5_1 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  Station2_5_2 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  Station2_5_3 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  Station2_5_4 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  Station2_5_5 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  Station2_5_6 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  Station2_5_7 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  Station2_6_0 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  Station2_6_1 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  Station2_6_2 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  Station2_6_3 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  Station2_6_4 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  Station2_6_5 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  Station2_6_6 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  Station2_6_7 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  Station2_7_0 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  Station2_7_1 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  Station2_7_2 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  Station2_7_3 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  Station2_7_4 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  Station2_7_5 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  Station2_7_6 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  Station2_7_7 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  Station3_0_0 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  Station3_0_1 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  Station3_0_2 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  Station3_0_3 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  Station3_0_4 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  Station3_0_5 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  Station3_0_6 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  Station3_0_7 = _RAND_72[15:0];
  _RAND_73 = {1{`RANDOM}};
  Station3_1_0 = _RAND_73[15:0];
  _RAND_74 = {1{`RANDOM}};
  Station3_1_1 = _RAND_74[15:0];
  _RAND_75 = {1{`RANDOM}};
  Station3_1_2 = _RAND_75[15:0];
  _RAND_76 = {1{`RANDOM}};
  Station3_1_3 = _RAND_76[15:0];
  _RAND_77 = {1{`RANDOM}};
  Station3_1_4 = _RAND_77[15:0];
  _RAND_78 = {1{`RANDOM}};
  Station3_1_5 = _RAND_78[15:0];
  _RAND_79 = {1{`RANDOM}};
  Station3_1_6 = _RAND_79[15:0];
  _RAND_80 = {1{`RANDOM}};
  Station3_1_7 = _RAND_80[15:0];
  _RAND_81 = {1{`RANDOM}};
  Station3_2_0 = _RAND_81[15:0];
  _RAND_82 = {1{`RANDOM}};
  Station3_2_1 = _RAND_82[15:0];
  _RAND_83 = {1{`RANDOM}};
  Station3_2_2 = _RAND_83[15:0];
  _RAND_84 = {1{`RANDOM}};
  Station3_2_3 = _RAND_84[15:0];
  _RAND_85 = {1{`RANDOM}};
  Station3_2_4 = _RAND_85[15:0];
  _RAND_86 = {1{`RANDOM}};
  Station3_2_5 = _RAND_86[15:0];
  _RAND_87 = {1{`RANDOM}};
  Station3_2_6 = _RAND_87[15:0];
  _RAND_88 = {1{`RANDOM}};
  Station3_2_7 = _RAND_88[15:0];
  _RAND_89 = {1{`RANDOM}};
  Station3_3_0 = _RAND_89[15:0];
  _RAND_90 = {1{`RANDOM}};
  Station3_3_1 = _RAND_90[15:0];
  _RAND_91 = {1{`RANDOM}};
  Station3_3_2 = _RAND_91[15:0];
  _RAND_92 = {1{`RANDOM}};
  Station3_3_3 = _RAND_92[15:0];
  _RAND_93 = {1{`RANDOM}};
  Station3_3_4 = _RAND_93[15:0];
  _RAND_94 = {1{`RANDOM}};
  Station3_3_5 = _RAND_94[15:0];
  _RAND_95 = {1{`RANDOM}};
  Station3_3_6 = _RAND_95[15:0];
  _RAND_96 = {1{`RANDOM}};
  Station3_3_7 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  Station3_4_0 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  Station3_4_1 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  Station3_4_2 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  Station3_4_3 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  Station3_4_4 = _RAND_101[15:0];
  _RAND_102 = {1{`RANDOM}};
  Station3_4_5 = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  Station3_4_6 = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  Station3_4_7 = _RAND_104[15:0];
  _RAND_105 = {1{`RANDOM}};
  Station3_5_0 = _RAND_105[15:0];
  _RAND_106 = {1{`RANDOM}};
  Station3_5_1 = _RAND_106[15:0];
  _RAND_107 = {1{`RANDOM}};
  Station3_5_2 = _RAND_107[15:0];
  _RAND_108 = {1{`RANDOM}};
  Station3_5_3 = _RAND_108[15:0];
  _RAND_109 = {1{`RANDOM}};
  Station3_5_4 = _RAND_109[15:0];
  _RAND_110 = {1{`RANDOM}};
  Station3_5_5 = _RAND_110[15:0];
  _RAND_111 = {1{`RANDOM}};
  Station3_5_6 = _RAND_111[15:0];
  _RAND_112 = {1{`RANDOM}};
  Station3_5_7 = _RAND_112[15:0];
  _RAND_113 = {1{`RANDOM}};
  Station3_6_0 = _RAND_113[15:0];
  _RAND_114 = {1{`RANDOM}};
  Station3_6_1 = _RAND_114[15:0];
  _RAND_115 = {1{`RANDOM}};
  Station3_6_2 = _RAND_115[15:0];
  _RAND_116 = {1{`RANDOM}};
  Station3_6_3 = _RAND_116[15:0];
  _RAND_117 = {1{`RANDOM}};
  Station3_6_4 = _RAND_117[15:0];
  _RAND_118 = {1{`RANDOM}};
  Station3_6_5 = _RAND_118[15:0];
  _RAND_119 = {1{`RANDOM}};
  Station3_6_6 = _RAND_119[15:0];
  _RAND_120 = {1{`RANDOM}};
  Station3_6_7 = _RAND_120[15:0];
  _RAND_121 = {1{`RANDOM}};
  Station3_7_0 = _RAND_121[15:0];
  _RAND_122 = {1{`RANDOM}};
  Station3_7_1 = _RAND_122[15:0];
  _RAND_123 = {1{`RANDOM}};
  Station3_7_2 = _RAND_123[15:0];
  _RAND_124 = {1{`RANDOM}};
  Station3_7_3 = _RAND_124[15:0];
  _RAND_125 = {1{`RANDOM}};
  Station3_7_4 = _RAND_125[15:0];
  _RAND_126 = {1{`RANDOM}};
  Station3_7_5 = _RAND_126[15:0];
  _RAND_127 = {1{`RANDOM}};
  Station3_7_6 = _RAND_127[15:0];
  _RAND_128 = {1{`RANDOM}};
  Station3_7_7 = _RAND_128[15:0];
  _RAND_129 = {1{`RANDOM}};
  Station4_0_0 = _RAND_129[15:0];
  _RAND_130 = {1{`RANDOM}};
  Station4_0_1 = _RAND_130[15:0];
  _RAND_131 = {1{`RANDOM}};
  Station4_0_2 = _RAND_131[15:0];
  _RAND_132 = {1{`RANDOM}};
  Station4_0_3 = _RAND_132[15:0];
  _RAND_133 = {1{`RANDOM}};
  Station4_0_4 = _RAND_133[15:0];
  _RAND_134 = {1{`RANDOM}};
  Station4_0_5 = _RAND_134[15:0];
  _RAND_135 = {1{`RANDOM}};
  Station4_0_6 = _RAND_135[15:0];
  _RAND_136 = {1{`RANDOM}};
  Station4_0_7 = _RAND_136[15:0];
  _RAND_137 = {1{`RANDOM}};
  Station4_1_0 = _RAND_137[15:0];
  _RAND_138 = {1{`RANDOM}};
  Station4_1_1 = _RAND_138[15:0];
  _RAND_139 = {1{`RANDOM}};
  Station4_1_2 = _RAND_139[15:0];
  _RAND_140 = {1{`RANDOM}};
  Station4_1_3 = _RAND_140[15:0];
  _RAND_141 = {1{`RANDOM}};
  Station4_1_4 = _RAND_141[15:0];
  _RAND_142 = {1{`RANDOM}};
  Station4_1_5 = _RAND_142[15:0];
  _RAND_143 = {1{`RANDOM}};
  Station4_1_6 = _RAND_143[15:0];
  _RAND_144 = {1{`RANDOM}};
  Station4_1_7 = _RAND_144[15:0];
  _RAND_145 = {1{`RANDOM}};
  Station4_2_0 = _RAND_145[15:0];
  _RAND_146 = {1{`RANDOM}};
  Station4_2_1 = _RAND_146[15:0];
  _RAND_147 = {1{`RANDOM}};
  Station4_2_2 = _RAND_147[15:0];
  _RAND_148 = {1{`RANDOM}};
  Station4_2_3 = _RAND_148[15:0];
  _RAND_149 = {1{`RANDOM}};
  Station4_2_4 = _RAND_149[15:0];
  _RAND_150 = {1{`RANDOM}};
  Station4_2_5 = _RAND_150[15:0];
  _RAND_151 = {1{`RANDOM}};
  Station4_2_6 = _RAND_151[15:0];
  _RAND_152 = {1{`RANDOM}};
  Station4_2_7 = _RAND_152[15:0];
  _RAND_153 = {1{`RANDOM}};
  Station4_3_0 = _RAND_153[15:0];
  _RAND_154 = {1{`RANDOM}};
  Station4_3_1 = _RAND_154[15:0];
  _RAND_155 = {1{`RANDOM}};
  Station4_3_2 = _RAND_155[15:0];
  _RAND_156 = {1{`RANDOM}};
  Station4_3_3 = _RAND_156[15:0];
  _RAND_157 = {1{`RANDOM}};
  Station4_3_4 = _RAND_157[15:0];
  _RAND_158 = {1{`RANDOM}};
  Station4_3_5 = _RAND_158[15:0];
  _RAND_159 = {1{`RANDOM}};
  Station4_3_6 = _RAND_159[15:0];
  _RAND_160 = {1{`RANDOM}};
  Station4_3_7 = _RAND_160[15:0];
  _RAND_161 = {1{`RANDOM}};
  Station4_4_0 = _RAND_161[15:0];
  _RAND_162 = {1{`RANDOM}};
  Station4_4_1 = _RAND_162[15:0];
  _RAND_163 = {1{`RANDOM}};
  Station4_4_2 = _RAND_163[15:0];
  _RAND_164 = {1{`RANDOM}};
  Station4_4_3 = _RAND_164[15:0];
  _RAND_165 = {1{`RANDOM}};
  Station4_4_4 = _RAND_165[15:0];
  _RAND_166 = {1{`RANDOM}};
  Station4_4_5 = _RAND_166[15:0];
  _RAND_167 = {1{`RANDOM}};
  Station4_4_6 = _RAND_167[15:0];
  _RAND_168 = {1{`RANDOM}};
  Station4_4_7 = _RAND_168[15:0];
  _RAND_169 = {1{`RANDOM}};
  Station4_5_0 = _RAND_169[15:0];
  _RAND_170 = {1{`RANDOM}};
  Station4_5_1 = _RAND_170[15:0];
  _RAND_171 = {1{`RANDOM}};
  Station4_5_2 = _RAND_171[15:0];
  _RAND_172 = {1{`RANDOM}};
  Station4_5_3 = _RAND_172[15:0];
  _RAND_173 = {1{`RANDOM}};
  Station4_5_4 = _RAND_173[15:0];
  _RAND_174 = {1{`RANDOM}};
  Station4_5_5 = _RAND_174[15:0];
  _RAND_175 = {1{`RANDOM}};
  Station4_5_6 = _RAND_175[15:0];
  _RAND_176 = {1{`RANDOM}};
  Station4_5_7 = _RAND_176[15:0];
  _RAND_177 = {1{`RANDOM}};
  Station4_6_0 = _RAND_177[15:0];
  _RAND_178 = {1{`RANDOM}};
  Station4_6_1 = _RAND_178[15:0];
  _RAND_179 = {1{`RANDOM}};
  Station4_6_2 = _RAND_179[15:0];
  _RAND_180 = {1{`RANDOM}};
  Station4_6_3 = _RAND_180[15:0];
  _RAND_181 = {1{`RANDOM}};
  Station4_6_4 = _RAND_181[15:0];
  _RAND_182 = {1{`RANDOM}};
  Station4_6_5 = _RAND_182[15:0];
  _RAND_183 = {1{`RANDOM}};
  Station4_6_6 = _RAND_183[15:0];
  _RAND_184 = {1{`RANDOM}};
  Station4_6_7 = _RAND_184[15:0];
  _RAND_185 = {1{`RANDOM}};
  Station4_7_0 = _RAND_185[15:0];
  _RAND_186 = {1{`RANDOM}};
  Station4_7_1 = _RAND_186[15:0];
  _RAND_187 = {1{`RANDOM}};
  Station4_7_2 = _RAND_187[15:0];
  _RAND_188 = {1{`RANDOM}};
  Station4_7_3 = _RAND_188[15:0];
  _RAND_189 = {1{`RANDOM}};
  Station4_7_4 = _RAND_189[15:0];
  _RAND_190 = {1{`RANDOM}};
  Station4_7_5 = _RAND_190[15:0];
  _RAND_191 = {1{`RANDOM}};
  Station4_7_6 = _RAND_191[15:0];
  _RAND_192 = {1{`RANDOM}};
  Station4_7_7 = _RAND_192[15:0];
  _RAND_193 = {1{`RANDOM}};
  Station5_0_0 = _RAND_193[15:0];
  _RAND_194 = {1{`RANDOM}};
  Station5_0_1 = _RAND_194[15:0];
  _RAND_195 = {1{`RANDOM}};
  Station5_0_2 = _RAND_195[15:0];
  _RAND_196 = {1{`RANDOM}};
  Station5_0_3 = _RAND_196[15:0];
  _RAND_197 = {1{`RANDOM}};
  Station5_0_4 = _RAND_197[15:0];
  _RAND_198 = {1{`RANDOM}};
  Station5_0_5 = _RAND_198[15:0];
  _RAND_199 = {1{`RANDOM}};
  Station5_0_6 = _RAND_199[15:0];
  _RAND_200 = {1{`RANDOM}};
  Station5_0_7 = _RAND_200[15:0];
  _RAND_201 = {1{`RANDOM}};
  Station5_1_0 = _RAND_201[15:0];
  _RAND_202 = {1{`RANDOM}};
  Station5_1_1 = _RAND_202[15:0];
  _RAND_203 = {1{`RANDOM}};
  Station5_1_2 = _RAND_203[15:0];
  _RAND_204 = {1{`RANDOM}};
  Station5_1_3 = _RAND_204[15:0];
  _RAND_205 = {1{`RANDOM}};
  Station5_1_4 = _RAND_205[15:0];
  _RAND_206 = {1{`RANDOM}};
  Station5_1_5 = _RAND_206[15:0];
  _RAND_207 = {1{`RANDOM}};
  Station5_1_6 = _RAND_207[15:0];
  _RAND_208 = {1{`RANDOM}};
  Station5_1_7 = _RAND_208[15:0];
  _RAND_209 = {1{`RANDOM}};
  Station5_2_0 = _RAND_209[15:0];
  _RAND_210 = {1{`RANDOM}};
  Station5_2_1 = _RAND_210[15:0];
  _RAND_211 = {1{`RANDOM}};
  Station5_2_2 = _RAND_211[15:0];
  _RAND_212 = {1{`RANDOM}};
  Station5_2_3 = _RAND_212[15:0];
  _RAND_213 = {1{`RANDOM}};
  Station5_2_4 = _RAND_213[15:0];
  _RAND_214 = {1{`RANDOM}};
  Station5_2_5 = _RAND_214[15:0];
  _RAND_215 = {1{`RANDOM}};
  Station5_2_6 = _RAND_215[15:0];
  _RAND_216 = {1{`RANDOM}};
  Station5_2_7 = _RAND_216[15:0];
  _RAND_217 = {1{`RANDOM}};
  Station5_3_0 = _RAND_217[15:0];
  _RAND_218 = {1{`RANDOM}};
  Station5_3_1 = _RAND_218[15:0];
  _RAND_219 = {1{`RANDOM}};
  Station5_3_2 = _RAND_219[15:0];
  _RAND_220 = {1{`RANDOM}};
  Station5_3_3 = _RAND_220[15:0];
  _RAND_221 = {1{`RANDOM}};
  Station5_3_4 = _RAND_221[15:0];
  _RAND_222 = {1{`RANDOM}};
  Station5_3_5 = _RAND_222[15:0];
  _RAND_223 = {1{`RANDOM}};
  Station5_3_6 = _RAND_223[15:0];
  _RAND_224 = {1{`RANDOM}};
  Station5_3_7 = _RAND_224[15:0];
  _RAND_225 = {1{`RANDOM}};
  Station5_4_0 = _RAND_225[15:0];
  _RAND_226 = {1{`RANDOM}};
  Station5_4_1 = _RAND_226[15:0];
  _RAND_227 = {1{`RANDOM}};
  Station5_4_2 = _RAND_227[15:0];
  _RAND_228 = {1{`RANDOM}};
  Station5_4_3 = _RAND_228[15:0];
  _RAND_229 = {1{`RANDOM}};
  Station5_4_4 = _RAND_229[15:0];
  _RAND_230 = {1{`RANDOM}};
  Station5_4_5 = _RAND_230[15:0];
  _RAND_231 = {1{`RANDOM}};
  Station5_4_6 = _RAND_231[15:0];
  _RAND_232 = {1{`RANDOM}};
  Station5_4_7 = _RAND_232[15:0];
  _RAND_233 = {1{`RANDOM}};
  Station5_5_0 = _RAND_233[15:0];
  _RAND_234 = {1{`RANDOM}};
  Station5_5_1 = _RAND_234[15:0];
  _RAND_235 = {1{`RANDOM}};
  Station5_5_2 = _RAND_235[15:0];
  _RAND_236 = {1{`RANDOM}};
  Station5_5_3 = _RAND_236[15:0];
  _RAND_237 = {1{`RANDOM}};
  Station5_5_4 = _RAND_237[15:0];
  _RAND_238 = {1{`RANDOM}};
  Station5_5_5 = _RAND_238[15:0];
  _RAND_239 = {1{`RANDOM}};
  Station5_5_6 = _RAND_239[15:0];
  _RAND_240 = {1{`RANDOM}};
  Station5_5_7 = _RAND_240[15:0];
  _RAND_241 = {1{`RANDOM}};
  Station5_6_0 = _RAND_241[15:0];
  _RAND_242 = {1{`RANDOM}};
  Station5_6_1 = _RAND_242[15:0];
  _RAND_243 = {1{`RANDOM}};
  Station5_6_2 = _RAND_243[15:0];
  _RAND_244 = {1{`RANDOM}};
  Station5_6_3 = _RAND_244[15:0];
  _RAND_245 = {1{`RANDOM}};
  Station5_6_4 = _RAND_245[15:0];
  _RAND_246 = {1{`RANDOM}};
  Station5_6_5 = _RAND_246[15:0];
  _RAND_247 = {1{`RANDOM}};
  Station5_6_6 = _RAND_247[15:0];
  _RAND_248 = {1{`RANDOM}};
  Station5_6_7 = _RAND_248[15:0];
  _RAND_249 = {1{`RANDOM}};
  Station5_7_0 = _RAND_249[15:0];
  _RAND_250 = {1{`RANDOM}};
  Station5_7_1 = _RAND_250[15:0];
  _RAND_251 = {1{`RANDOM}};
  Station5_7_2 = _RAND_251[15:0];
  _RAND_252 = {1{`RANDOM}};
  Station5_7_3 = _RAND_252[15:0];
  _RAND_253 = {1{`RANDOM}};
  Station5_7_4 = _RAND_253[15:0];
  _RAND_254 = {1{`RANDOM}};
  Station5_7_5 = _RAND_254[15:0];
  _RAND_255 = {1{`RANDOM}};
  Station5_7_6 = _RAND_255[15:0];
  _RAND_256 = {1{`RANDOM}};
  Station5_7_7 = _RAND_256[15:0];
  _RAND_257 = {1{`RANDOM}};
  Station6_0_0 = _RAND_257[15:0];
  _RAND_258 = {1{`RANDOM}};
  Station6_0_1 = _RAND_258[15:0];
  _RAND_259 = {1{`RANDOM}};
  Station6_0_2 = _RAND_259[15:0];
  _RAND_260 = {1{`RANDOM}};
  Station6_0_3 = _RAND_260[15:0];
  _RAND_261 = {1{`RANDOM}};
  Station6_0_4 = _RAND_261[15:0];
  _RAND_262 = {1{`RANDOM}};
  Station6_0_5 = _RAND_262[15:0];
  _RAND_263 = {1{`RANDOM}};
  Station6_0_6 = _RAND_263[15:0];
  _RAND_264 = {1{`RANDOM}};
  Station6_0_7 = _RAND_264[15:0];
  _RAND_265 = {1{`RANDOM}};
  Station6_1_0 = _RAND_265[15:0];
  _RAND_266 = {1{`RANDOM}};
  Station6_1_1 = _RAND_266[15:0];
  _RAND_267 = {1{`RANDOM}};
  Station6_1_2 = _RAND_267[15:0];
  _RAND_268 = {1{`RANDOM}};
  Station6_1_3 = _RAND_268[15:0];
  _RAND_269 = {1{`RANDOM}};
  Station6_1_4 = _RAND_269[15:0];
  _RAND_270 = {1{`RANDOM}};
  Station6_1_5 = _RAND_270[15:0];
  _RAND_271 = {1{`RANDOM}};
  Station6_1_6 = _RAND_271[15:0];
  _RAND_272 = {1{`RANDOM}};
  Station6_1_7 = _RAND_272[15:0];
  _RAND_273 = {1{`RANDOM}};
  Station6_2_0 = _RAND_273[15:0];
  _RAND_274 = {1{`RANDOM}};
  Station6_2_1 = _RAND_274[15:0];
  _RAND_275 = {1{`RANDOM}};
  Station6_2_2 = _RAND_275[15:0];
  _RAND_276 = {1{`RANDOM}};
  Station6_2_3 = _RAND_276[15:0];
  _RAND_277 = {1{`RANDOM}};
  Station6_2_4 = _RAND_277[15:0];
  _RAND_278 = {1{`RANDOM}};
  Station6_2_5 = _RAND_278[15:0];
  _RAND_279 = {1{`RANDOM}};
  Station6_2_6 = _RAND_279[15:0];
  _RAND_280 = {1{`RANDOM}};
  Station6_2_7 = _RAND_280[15:0];
  _RAND_281 = {1{`RANDOM}};
  Station6_3_0 = _RAND_281[15:0];
  _RAND_282 = {1{`RANDOM}};
  Station6_3_1 = _RAND_282[15:0];
  _RAND_283 = {1{`RANDOM}};
  Station6_3_2 = _RAND_283[15:0];
  _RAND_284 = {1{`RANDOM}};
  Station6_3_3 = _RAND_284[15:0];
  _RAND_285 = {1{`RANDOM}};
  Station6_3_4 = _RAND_285[15:0];
  _RAND_286 = {1{`RANDOM}};
  Station6_3_5 = _RAND_286[15:0];
  _RAND_287 = {1{`RANDOM}};
  Station6_3_6 = _RAND_287[15:0];
  _RAND_288 = {1{`RANDOM}};
  Station6_3_7 = _RAND_288[15:0];
  _RAND_289 = {1{`RANDOM}};
  Station6_4_0 = _RAND_289[15:0];
  _RAND_290 = {1{`RANDOM}};
  Station6_4_1 = _RAND_290[15:0];
  _RAND_291 = {1{`RANDOM}};
  Station6_4_2 = _RAND_291[15:0];
  _RAND_292 = {1{`RANDOM}};
  Station6_4_3 = _RAND_292[15:0];
  _RAND_293 = {1{`RANDOM}};
  Station6_4_4 = _RAND_293[15:0];
  _RAND_294 = {1{`RANDOM}};
  Station6_4_5 = _RAND_294[15:0];
  _RAND_295 = {1{`RANDOM}};
  Station6_4_6 = _RAND_295[15:0];
  _RAND_296 = {1{`RANDOM}};
  Station6_4_7 = _RAND_296[15:0];
  _RAND_297 = {1{`RANDOM}};
  Station6_5_0 = _RAND_297[15:0];
  _RAND_298 = {1{`RANDOM}};
  Station6_5_1 = _RAND_298[15:0];
  _RAND_299 = {1{`RANDOM}};
  Station6_5_2 = _RAND_299[15:0];
  _RAND_300 = {1{`RANDOM}};
  Station6_5_3 = _RAND_300[15:0];
  _RAND_301 = {1{`RANDOM}};
  Station6_5_4 = _RAND_301[15:0];
  _RAND_302 = {1{`RANDOM}};
  Station6_5_5 = _RAND_302[15:0];
  _RAND_303 = {1{`RANDOM}};
  Station6_5_6 = _RAND_303[15:0];
  _RAND_304 = {1{`RANDOM}};
  Station6_5_7 = _RAND_304[15:0];
  _RAND_305 = {1{`RANDOM}};
  Station6_6_0 = _RAND_305[15:0];
  _RAND_306 = {1{`RANDOM}};
  Station6_6_1 = _RAND_306[15:0];
  _RAND_307 = {1{`RANDOM}};
  Station6_6_2 = _RAND_307[15:0];
  _RAND_308 = {1{`RANDOM}};
  Station6_6_3 = _RAND_308[15:0];
  _RAND_309 = {1{`RANDOM}};
  Station6_6_4 = _RAND_309[15:0];
  _RAND_310 = {1{`RANDOM}};
  Station6_6_5 = _RAND_310[15:0];
  _RAND_311 = {1{`RANDOM}};
  Station6_6_6 = _RAND_311[15:0];
  _RAND_312 = {1{`RANDOM}};
  Station6_6_7 = _RAND_312[15:0];
  _RAND_313 = {1{`RANDOM}};
  Station6_7_0 = _RAND_313[15:0];
  _RAND_314 = {1{`RANDOM}};
  Station6_7_1 = _RAND_314[15:0];
  _RAND_315 = {1{`RANDOM}};
  Station6_7_2 = _RAND_315[15:0];
  _RAND_316 = {1{`RANDOM}};
  Station6_7_3 = _RAND_316[15:0];
  _RAND_317 = {1{`RANDOM}};
  Station6_7_4 = _RAND_317[15:0];
  _RAND_318 = {1{`RANDOM}};
  Station6_7_5 = _RAND_318[15:0];
  _RAND_319 = {1{`RANDOM}};
  Station6_7_6 = _RAND_319[15:0];
  _RAND_320 = {1{`RANDOM}};
  Station6_7_7 = _RAND_320[15:0];
  _RAND_321 = {1{`RANDOM}};
  Station7_0_0 = _RAND_321[15:0];
  _RAND_322 = {1{`RANDOM}};
  Station7_0_1 = _RAND_322[15:0];
  _RAND_323 = {1{`RANDOM}};
  Station7_0_2 = _RAND_323[15:0];
  _RAND_324 = {1{`RANDOM}};
  Station7_0_3 = _RAND_324[15:0];
  _RAND_325 = {1{`RANDOM}};
  Station7_0_4 = _RAND_325[15:0];
  _RAND_326 = {1{`RANDOM}};
  Station7_0_5 = _RAND_326[15:0];
  _RAND_327 = {1{`RANDOM}};
  Station7_0_6 = _RAND_327[15:0];
  _RAND_328 = {1{`RANDOM}};
  Station7_0_7 = _RAND_328[15:0];
  _RAND_329 = {1{`RANDOM}};
  Station7_1_0 = _RAND_329[15:0];
  _RAND_330 = {1{`RANDOM}};
  Station7_1_1 = _RAND_330[15:0];
  _RAND_331 = {1{`RANDOM}};
  Station7_1_2 = _RAND_331[15:0];
  _RAND_332 = {1{`RANDOM}};
  Station7_1_3 = _RAND_332[15:0];
  _RAND_333 = {1{`RANDOM}};
  Station7_1_4 = _RAND_333[15:0];
  _RAND_334 = {1{`RANDOM}};
  Station7_1_5 = _RAND_334[15:0];
  _RAND_335 = {1{`RANDOM}};
  Station7_1_6 = _RAND_335[15:0];
  _RAND_336 = {1{`RANDOM}};
  Station7_1_7 = _RAND_336[15:0];
  _RAND_337 = {1{`RANDOM}};
  Station7_2_0 = _RAND_337[15:0];
  _RAND_338 = {1{`RANDOM}};
  Station7_2_1 = _RAND_338[15:0];
  _RAND_339 = {1{`RANDOM}};
  Station7_2_2 = _RAND_339[15:0];
  _RAND_340 = {1{`RANDOM}};
  Station7_2_3 = _RAND_340[15:0];
  _RAND_341 = {1{`RANDOM}};
  Station7_2_4 = _RAND_341[15:0];
  _RAND_342 = {1{`RANDOM}};
  Station7_2_5 = _RAND_342[15:0];
  _RAND_343 = {1{`RANDOM}};
  Station7_2_6 = _RAND_343[15:0];
  _RAND_344 = {1{`RANDOM}};
  Station7_2_7 = _RAND_344[15:0];
  _RAND_345 = {1{`RANDOM}};
  Station7_3_0 = _RAND_345[15:0];
  _RAND_346 = {1{`RANDOM}};
  Station7_3_1 = _RAND_346[15:0];
  _RAND_347 = {1{`RANDOM}};
  Station7_3_2 = _RAND_347[15:0];
  _RAND_348 = {1{`RANDOM}};
  Station7_3_3 = _RAND_348[15:0];
  _RAND_349 = {1{`RANDOM}};
  Station7_3_4 = _RAND_349[15:0];
  _RAND_350 = {1{`RANDOM}};
  Station7_3_5 = _RAND_350[15:0];
  _RAND_351 = {1{`RANDOM}};
  Station7_3_6 = _RAND_351[15:0];
  _RAND_352 = {1{`RANDOM}};
  Station7_3_7 = _RAND_352[15:0];
  _RAND_353 = {1{`RANDOM}};
  Station7_4_0 = _RAND_353[15:0];
  _RAND_354 = {1{`RANDOM}};
  Station7_4_1 = _RAND_354[15:0];
  _RAND_355 = {1{`RANDOM}};
  Station7_4_2 = _RAND_355[15:0];
  _RAND_356 = {1{`RANDOM}};
  Station7_4_3 = _RAND_356[15:0];
  _RAND_357 = {1{`RANDOM}};
  Station7_4_4 = _RAND_357[15:0];
  _RAND_358 = {1{`RANDOM}};
  Station7_4_5 = _RAND_358[15:0];
  _RAND_359 = {1{`RANDOM}};
  Station7_4_6 = _RAND_359[15:0];
  _RAND_360 = {1{`RANDOM}};
  Station7_4_7 = _RAND_360[15:0];
  _RAND_361 = {1{`RANDOM}};
  Station7_5_0 = _RAND_361[15:0];
  _RAND_362 = {1{`RANDOM}};
  Station7_5_1 = _RAND_362[15:0];
  _RAND_363 = {1{`RANDOM}};
  Station7_5_2 = _RAND_363[15:0];
  _RAND_364 = {1{`RANDOM}};
  Station7_5_3 = _RAND_364[15:0];
  _RAND_365 = {1{`RANDOM}};
  Station7_5_4 = _RAND_365[15:0];
  _RAND_366 = {1{`RANDOM}};
  Station7_5_5 = _RAND_366[15:0];
  _RAND_367 = {1{`RANDOM}};
  Station7_5_6 = _RAND_367[15:0];
  _RAND_368 = {1{`RANDOM}};
  Station7_5_7 = _RAND_368[15:0];
  _RAND_369 = {1{`RANDOM}};
  Station7_6_0 = _RAND_369[15:0];
  _RAND_370 = {1{`RANDOM}};
  Station7_6_1 = _RAND_370[15:0];
  _RAND_371 = {1{`RANDOM}};
  Station7_6_2 = _RAND_371[15:0];
  _RAND_372 = {1{`RANDOM}};
  Station7_6_3 = _RAND_372[15:0];
  _RAND_373 = {1{`RANDOM}};
  Station7_6_4 = _RAND_373[15:0];
  _RAND_374 = {1{`RANDOM}};
  Station7_6_5 = _RAND_374[15:0];
  _RAND_375 = {1{`RANDOM}};
  Station7_6_6 = _RAND_375[15:0];
  _RAND_376 = {1{`RANDOM}};
  Station7_6_7 = _RAND_376[15:0];
  _RAND_377 = {1{`RANDOM}};
  Station7_7_0 = _RAND_377[15:0];
  _RAND_378 = {1{`RANDOM}};
  Station7_7_1 = _RAND_378[15:0];
  _RAND_379 = {1{`RANDOM}};
  Station7_7_2 = _RAND_379[15:0];
  _RAND_380 = {1{`RANDOM}};
  Station7_7_3 = _RAND_380[15:0];
  _RAND_381 = {1{`RANDOM}};
  Station7_7_4 = _RAND_381[15:0];
  _RAND_382 = {1{`RANDOM}};
  Station7_7_5 = _RAND_382[15:0];
  _RAND_383 = {1{`RANDOM}};
  Station7_7_6 = _RAND_383[15:0];
  _RAND_384 = {1{`RANDOM}};
  Station7_7_7 = _RAND_384[15:0];
  _RAND_385 = {1{`RANDOM}};
  Station8_0_0 = _RAND_385[15:0];
  _RAND_386 = {1{`RANDOM}};
  Station8_0_1 = _RAND_386[15:0];
  _RAND_387 = {1{`RANDOM}};
  Station8_0_2 = _RAND_387[15:0];
  _RAND_388 = {1{`RANDOM}};
  Station8_0_3 = _RAND_388[15:0];
  _RAND_389 = {1{`RANDOM}};
  Station8_0_4 = _RAND_389[15:0];
  _RAND_390 = {1{`RANDOM}};
  Station8_0_5 = _RAND_390[15:0];
  _RAND_391 = {1{`RANDOM}};
  Station8_0_6 = _RAND_391[15:0];
  _RAND_392 = {1{`RANDOM}};
  Station8_0_7 = _RAND_392[15:0];
  _RAND_393 = {1{`RANDOM}};
  Station8_1_0 = _RAND_393[15:0];
  _RAND_394 = {1{`RANDOM}};
  Station8_1_1 = _RAND_394[15:0];
  _RAND_395 = {1{`RANDOM}};
  Station8_1_2 = _RAND_395[15:0];
  _RAND_396 = {1{`RANDOM}};
  Station8_1_3 = _RAND_396[15:0];
  _RAND_397 = {1{`RANDOM}};
  Station8_1_4 = _RAND_397[15:0];
  _RAND_398 = {1{`RANDOM}};
  Station8_1_5 = _RAND_398[15:0];
  _RAND_399 = {1{`RANDOM}};
  Station8_1_6 = _RAND_399[15:0];
  _RAND_400 = {1{`RANDOM}};
  Station8_1_7 = _RAND_400[15:0];
  _RAND_401 = {1{`RANDOM}};
  Station8_2_0 = _RAND_401[15:0];
  _RAND_402 = {1{`RANDOM}};
  Station8_2_1 = _RAND_402[15:0];
  _RAND_403 = {1{`RANDOM}};
  Station8_2_2 = _RAND_403[15:0];
  _RAND_404 = {1{`RANDOM}};
  Station8_2_3 = _RAND_404[15:0];
  _RAND_405 = {1{`RANDOM}};
  Station8_2_4 = _RAND_405[15:0];
  _RAND_406 = {1{`RANDOM}};
  Station8_2_5 = _RAND_406[15:0];
  _RAND_407 = {1{`RANDOM}};
  Station8_2_6 = _RAND_407[15:0];
  _RAND_408 = {1{`RANDOM}};
  Station8_2_7 = _RAND_408[15:0];
  _RAND_409 = {1{`RANDOM}};
  Station8_3_0 = _RAND_409[15:0];
  _RAND_410 = {1{`RANDOM}};
  Station8_3_1 = _RAND_410[15:0];
  _RAND_411 = {1{`RANDOM}};
  Station8_3_2 = _RAND_411[15:0];
  _RAND_412 = {1{`RANDOM}};
  Station8_3_3 = _RAND_412[15:0];
  _RAND_413 = {1{`RANDOM}};
  Station8_3_4 = _RAND_413[15:0];
  _RAND_414 = {1{`RANDOM}};
  Station8_3_5 = _RAND_414[15:0];
  _RAND_415 = {1{`RANDOM}};
  Station8_3_6 = _RAND_415[15:0];
  _RAND_416 = {1{`RANDOM}};
  Station8_3_7 = _RAND_416[15:0];
  _RAND_417 = {1{`RANDOM}};
  Station8_4_0 = _RAND_417[15:0];
  _RAND_418 = {1{`RANDOM}};
  Station8_4_1 = _RAND_418[15:0];
  _RAND_419 = {1{`RANDOM}};
  Station8_4_2 = _RAND_419[15:0];
  _RAND_420 = {1{`RANDOM}};
  Station8_4_3 = _RAND_420[15:0];
  _RAND_421 = {1{`RANDOM}};
  Station8_4_4 = _RAND_421[15:0];
  _RAND_422 = {1{`RANDOM}};
  Station8_4_5 = _RAND_422[15:0];
  _RAND_423 = {1{`RANDOM}};
  Station8_4_6 = _RAND_423[15:0];
  _RAND_424 = {1{`RANDOM}};
  Station8_4_7 = _RAND_424[15:0];
  _RAND_425 = {1{`RANDOM}};
  Station8_5_0 = _RAND_425[15:0];
  _RAND_426 = {1{`RANDOM}};
  Station8_5_1 = _RAND_426[15:0];
  _RAND_427 = {1{`RANDOM}};
  Station8_5_2 = _RAND_427[15:0];
  _RAND_428 = {1{`RANDOM}};
  Station8_5_3 = _RAND_428[15:0];
  _RAND_429 = {1{`RANDOM}};
  Station8_5_4 = _RAND_429[15:0];
  _RAND_430 = {1{`RANDOM}};
  Station8_5_5 = _RAND_430[15:0];
  _RAND_431 = {1{`RANDOM}};
  Station8_5_6 = _RAND_431[15:0];
  _RAND_432 = {1{`RANDOM}};
  Station8_5_7 = _RAND_432[15:0];
  _RAND_433 = {1{`RANDOM}};
  Station8_6_0 = _RAND_433[15:0];
  _RAND_434 = {1{`RANDOM}};
  Station8_6_1 = _RAND_434[15:0];
  _RAND_435 = {1{`RANDOM}};
  Station8_6_2 = _RAND_435[15:0];
  _RAND_436 = {1{`RANDOM}};
  Station8_6_3 = _RAND_436[15:0];
  _RAND_437 = {1{`RANDOM}};
  Station8_6_4 = _RAND_437[15:0];
  _RAND_438 = {1{`RANDOM}};
  Station8_6_5 = _RAND_438[15:0];
  _RAND_439 = {1{`RANDOM}};
  Station8_6_6 = _RAND_439[15:0];
  _RAND_440 = {1{`RANDOM}};
  Station8_6_7 = _RAND_440[15:0];
  _RAND_441 = {1{`RANDOM}};
  Station8_7_0 = _RAND_441[15:0];
  _RAND_442 = {1{`RANDOM}};
  Station8_7_1 = _RAND_442[15:0];
  _RAND_443 = {1{`RANDOM}};
  Station8_7_2 = _RAND_443[15:0];
  _RAND_444 = {1{`RANDOM}};
  Station8_7_3 = _RAND_444[15:0];
  _RAND_445 = {1{`RANDOM}};
  Station8_7_4 = _RAND_445[15:0];
  _RAND_446 = {1{`RANDOM}};
  Station8_7_5 = _RAND_446[15:0];
  _RAND_447 = {1{`RANDOM}};
  Station8_7_6 = _RAND_447[15:0];
  _RAND_448 = {1{`RANDOM}};
  Station8_7_7 = _RAND_448[15:0];
  _RAND_449 = {1{`RANDOM}};
  i = _RAND_449[31:0];
  _RAND_450 = {1{`RANDOM}};
  j = _RAND_450[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ivncontrol4(
  input         clock,
  input         reset,
  input  [15:0] io_Stationary_matrix_0_0,
  input  [15:0] io_Stationary_matrix_0_1,
  input  [15:0] io_Stationary_matrix_0_2,
  input  [15:0] io_Stationary_matrix_0_3,
  input  [15:0] io_Stationary_matrix_0_4,
  input  [15:0] io_Stationary_matrix_0_5,
  input  [15:0] io_Stationary_matrix_0_6,
  input  [15:0] io_Stationary_matrix_0_7,
  input  [15:0] io_Stationary_matrix_1_0,
  input  [15:0] io_Stationary_matrix_1_1,
  input  [15:0] io_Stationary_matrix_1_2,
  input  [15:0] io_Stationary_matrix_1_3,
  input  [15:0] io_Stationary_matrix_1_4,
  input  [15:0] io_Stationary_matrix_1_5,
  input  [15:0] io_Stationary_matrix_1_6,
  input  [15:0] io_Stationary_matrix_1_7,
  input  [15:0] io_Stationary_matrix_2_0,
  input  [15:0] io_Stationary_matrix_2_1,
  input  [15:0] io_Stationary_matrix_2_2,
  input  [15:0] io_Stationary_matrix_2_3,
  input  [15:0] io_Stationary_matrix_2_4,
  input  [15:0] io_Stationary_matrix_2_5,
  input  [15:0] io_Stationary_matrix_2_6,
  input  [15:0] io_Stationary_matrix_2_7,
  input  [15:0] io_Stationary_matrix_3_0,
  input  [15:0] io_Stationary_matrix_3_1,
  input  [15:0] io_Stationary_matrix_3_2,
  input  [15:0] io_Stationary_matrix_3_3,
  input  [15:0] io_Stationary_matrix_3_4,
  input  [15:0] io_Stationary_matrix_3_5,
  input  [15:0] io_Stationary_matrix_3_6,
  input  [15:0] io_Stationary_matrix_3_7,
  input  [15:0] io_Stationary_matrix_4_0,
  input  [15:0] io_Stationary_matrix_4_1,
  input  [15:0] io_Stationary_matrix_4_2,
  input  [15:0] io_Stationary_matrix_4_3,
  input  [15:0] io_Stationary_matrix_4_4,
  input  [15:0] io_Stationary_matrix_4_5,
  input  [15:0] io_Stationary_matrix_4_6,
  input  [15:0] io_Stationary_matrix_4_7,
  input  [15:0] io_Stationary_matrix_5_0,
  input  [15:0] io_Stationary_matrix_5_1,
  input  [15:0] io_Stationary_matrix_5_2,
  input  [15:0] io_Stationary_matrix_5_3,
  input  [15:0] io_Stationary_matrix_5_4,
  input  [15:0] io_Stationary_matrix_5_5,
  input  [15:0] io_Stationary_matrix_5_6,
  input  [15:0] io_Stationary_matrix_5_7,
  input  [15:0] io_Stationary_matrix_6_0,
  input  [15:0] io_Stationary_matrix_6_1,
  input  [15:0] io_Stationary_matrix_6_2,
  input  [15:0] io_Stationary_matrix_6_3,
  input  [15:0] io_Stationary_matrix_6_4,
  input  [15:0] io_Stationary_matrix_6_5,
  input  [15:0] io_Stationary_matrix_6_6,
  input  [15:0] io_Stationary_matrix_6_7,
  input  [15:0] io_Stationary_matrix_7_0,
  input  [15:0] io_Stationary_matrix_7_1,
  input  [15:0] io_Stationary_matrix_7_2,
  input  [15:0] io_Stationary_matrix_7_3,
  input  [15:0] io_Stationary_matrix_7_4,
  input  [15:0] io_Stationary_matrix_7_5,
  input  [15:0] io_Stationary_matrix_7_6,
  input  [15:0] io_Stationary_matrix_7_7,
  output [4:0]  io_o_vn_0,
  output [4:0]  io_o_vn_1,
  output [4:0]  io_o_vn_2,
  output [4:0]  io_o_vn_3,
  output [4:0]  io_o_vn2_0,
  output [4:0]  io_o_vn2_1,
  output [4:0]  io_o_vn2_2,
  output [4:0]  io_o_vn2_3,
  output        io_ProcessValid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
`endif // RANDOMIZE_REG_INIT
  reg [4:0] i_vn_0; // @[ivncontrol4.scala 16:23]
  reg [4:0] i_vn_1; // @[ivncontrol4.scala 16:23]
  reg [4:0] i_vn_2; // @[ivncontrol4.scala 16:23]
  reg [4:0] i_vn_3; // @[ivncontrol4.scala 16:23]
  reg [4:0] i_vn2_0; // @[ivncontrol4.scala 17:24]
  reg [4:0] i_vn2_1; // @[ivncontrol4.scala 17:24]
  reg [4:0] i_vn2_2; // @[ivncontrol4.scala 17:24]
  reg [4:0] i_vn2_3; // @[ivncontrol4.scala 17:24]
  reg [31:0] rowcount_0; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_1; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_2; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_3; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_4; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_5; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_6; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_7; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_8; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_9; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_10; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_11; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_12; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_13; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_14; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_15; // @[ivncontrol4.scala 21:27]
  reg [31:0] pin; // @[ivncontrol4.scala 31:22]
  reg [31:0] i; // @[ivncontrol4.scala 35:20]
  reg [31:0] j; // @[ivncontrol4.scala 36:20]
  wire  _k_T_1 = j == 32'h7; // @[ivncontrol4.scala 38:37]
  wire  _k_T_2 = i == 32'h7 & j == 32'h7; // @[ivncontrol4.scala 38:31]
  reg  k; // @[ivncontrol4.scala 38:20]
  reg  io_ProcessValid_REG; // @[ivncontrol4.scala 42:35]
  reg [31:0] mat_0_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_0_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_0_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_0_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_0_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_0_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_0_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_0_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] count_0; // @[ivncontrol4.scala 52:20]
  reg [31:0] count_1; // @[ivncontrol4.scala 52:20]
  reg [31:0] count_2; // @[ivncontrol4.scala 52:20]
  reg [31:0] count_3; // @[ivncontrol4.scala 52:20]
  reg [31:0] count_4; // @[ivncontrol4.scala 52:20]
  reg [31:0] count_5; // @[ivncontrol4.scala 52:20]
  reg [31:0] count_6; // @[ivncontrol4.scala 52:20]
  reg [31:0] count_7; // @[ivncontrol4.scala 52:20]
  wire [15:0] _GEN_66 = 3'h0 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_0_1 : io_Stationary_matrix_0_0; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_67 = 3'h0 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_0_2 : _GEN_66; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_68 = 3'h0 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_0_3 : _GEN_67; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_69 = 3'h0 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_0_4 : _GEN_68; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_70 = 3'h0 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_0_5 : _GEN_69; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_71 = 3'h0 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_0_6 : _GEN_70; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_72 = 3'h0 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_0_7 : _GEN_71; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_73 = 3'h1 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_1_0 : _GEN_72; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_74 = 3'h1 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_1_1 : _GEN_73; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_75 = 3'h1 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_1_2 : _GEN_74; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_76 = 3'h1 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_1_3 : _GEN_75; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_77 = 3'h1 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_1_4 : _GEN_76; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_78 = 3'h1 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_1_5 : _GEN_77; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_79 = 3'h1 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_1_6 : _GEN_78; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_80 = 3'h1 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_1_7 : _GEN_79; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_81 = 3'h2 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_2_0 : _GEN_80; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_82 = 3'h2 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_2_1 : _GEN_81; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_83 = 3'h2 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_2_2 : _GEN_82; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_84 = 3'h2 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_2_3 : _GEN_83; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_85 = 3'h2 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_2_4 : _GEN_84; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_86 = 3'h2 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_2_5 : _GEN_85; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_87 = 3'h2 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_2_6 : _GEN_86; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_88 = 3'h2 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_2_7 : _GEN_87; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_89 = 3'h3 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_3_0 : _GEN_88; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_90 = 3'h3 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_3_1 : _GEN_89; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_91 = 3'h3 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_3_2 : _GEN_90; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_92 = 3'h3 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_3_3 : _GEN_91; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_93 = 3'h3 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_3_4 : _GEN_92; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_94 = 3'h3 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_3_5 : _GEN_93; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_95 = 3'h3 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_3_6 : _GEN_94; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_96 = 3'h3 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_3_7 : _GEN_95; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_97 = 3'h4 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_4_0 : _GEN_96; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_98 = 3'h4 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_4_1 : _GEN_97; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_99 = 3'h4 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_4_2 : _GEN_98; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_100 = 3'h4 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_4_3 : _GEN_99; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_101 = 3'h4 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_4_4 : _GEN_100; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_102 = 3'h4 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_4_5 : _GEN_101; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_103 = 3'h4 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_4_6 : _GEN_102; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_104 = 3'h4 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_4_7 : _GEN_103; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_105 = 3'h5 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_5_0 : _GEN_104; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_106 = 3'h5 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_5_1 : _GEN_105; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_107 = 3'h5 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_5_2 : _GEN_106; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_108 = 3'h5 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_5_3 : _GEN_107; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_109 = 3'h5 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_5_4 : _GEN_108; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_110 = 3'h5 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_5_5 : _GEN_109; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_111 = 3'h5 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_5_6 : _GEN_110; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_112 = 3'h5 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_5_7 : _GEN_111; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_113 = 3'h6 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_6_0 : _GEN_112; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_114 = 3'h6 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_6_1 : _GEN_113; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_115 = 3'h6 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_6_2 : _GEN_114; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_116 = 3'h6 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_6_3 : _GEN_115; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_117 = 3'h6 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_6_4 : _GEN_116; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_118 = 3'h6 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_6_5 : _GEN_117; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_119 = 3'h6 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_6_6 : _GEN_118; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_120 = 3'h6 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_6_7 : _GEN_119; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_121 = 3'h7 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_7_0 : _GEN_120; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_122 = 3'h7 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_7_1 : _GEN_121; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_123 = 3'h7 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_7_2 : _GEN_122; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_124 = 3'h7 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_7_3 : _GEN_123; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_125 = 3'h7 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_7_4 : _GEN_124; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_126 = 3'h7 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_7_5 : _GEN_125; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_127 = 3'h7 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_7_6 : _GEN_126; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_128 = 3'h7 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_7_7 : _GEN_127; // @[ivncontrol4.scala 57:{15,15}]
  wire [31:0] _mat_T_3_T_4 = {{16'd0}, _GEN_128}; // @[ivncontrol4.scala 57:{15,15}]
  wire  _GEN_225 = count_7 >= 32'h8; // @[ivncontrol4.scala 66:28 67:16]
  wire  valid1 = count_7 >= 32'h8; // @[ivncontrol4.scala 66:28 67:16]
  wire [31:0] _GEN_194 = 3'h1 == i[2:0] ? count_1 : count_0; // @[ivncontrol4.scala 60:{33,33}]
  wire [31:0] _GEN_195 = 3'h2 == i[2:0] ? count_2 : _GEN_194; // @[ivncontrol4.scala 60:{33,33}]
  wire [31:0] _GEN_196 = 3'h3 == i[2:0] ? count_3 : _GEN_195; // @[ivncontrol4.scala 60:{33,33}]
  wire [31:0] _GEN_197 = 3'h4 == i[2:0] ? count_4 : _GEN_196; // @[ivncontrol4.scala 60:{33,33}]
  wire [31:0] _GEN_198 = 3'h5 == i[2:0] ? count_5 : _GEN_197; // @[ivncontrol4.scala 60:{33,33}]
  wire [31:0] _GEN_199 = 3'h6 == i[2:0] ? count_6 : _GEN_198; // @[ivncontrol4.scala 60:{33,33}]
  wire [31:0] _GEN_200 = 3'h7 == i[2:0] ? count_7 : _GEN_199; // @[ivncontrol4.scala 60:{33,33}]
  wire [31:0] _count_T_2 = _GEN_200 + 32'h1; // @[ivncontrol4.scala 60:33]
  wire [31:0] _i_T_1 = i + 32'h1; // @[ivncontrol4.scala 104:16]
  wire [31:0] _j_T_1 = j + 32'h1; // @[ivncontrol4.scala 108:16]
  wire  _GEN_244 = _k_T_2; // @[ivncontrol4.scala 136:75 137:14 139:14]
  wire [31:0] _GEN_245 = rowcount_0 != 32'h0 ? 32'h0 : pin; // @[ivncontrol4.scala 145:30 146:13 31:22]
  wire  _T_27 = rowcount_0 == 32'h0; // @[ivncontrol4.scala 148:23]
  wire [31:0] _GEN_246 = rowcount_0 == 32'h0 & rowcount_1 != 32'h0 ? 32'h1 : _GEN_245; // @[ivncontrol4.scala 148:54 149:13]
  wire  _T_32 = _T_27 & rowcount_1 == 32'h0; // @[ivncontrol4.scala 151:31]
  wire [31:0] _GEN_247 = _T_27 & rowcount_1 == 32'h0 & rowcount_2 != 32'h0 ? 32'h2 : _GEN_246; // @[ivncontrol4.scala 151:77 152:13]
  wire  _T_39 = _T_32 & rowcount_2 == 32'h0; // @[ivncontrol4.scala 154:54]
  wire [31:0] _GEN_248 = _T_32 & rowcount_2 == 32'h0 & rowcount_3 != 32'h0 ? 32'h3 : _GEN_247; // @[ivncontrol4.scala 154:100 155:13]
  wire  _T_48 = _T_39 & rowcount_3 == 32'h0; // @[ivncontrol4.scala 157:77]
  wire [31:0] _GEN_249 = _T_39 & rowcount_3 == 32'h0 & rowcount_4 != 32'h0 ? 32'h4 : _GEN_248; // @[ivncontrol4.scala 157:123 158:13]
  wire  _T_59 = _T_48 & rowcount_4 == 32'h0; // @[ivncontrol4.scala 160:100]
  wire  _T_72 = _T_59 & rowcount_5 == 32'h0; // @[ivncontrol4.scala 163:123]
  wire  valid = _k_T_2; // @[ivncontrol4.scala 136:75 137:14 139:14]
  wire [32:0] _T_91 = {{1'd0}, pin}; // @[ivncontrol4.scala 174:27]
  wire [31:0] _GEN_254 = 4'h1 == _T_91[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_255 = 4'h2 == _T_91[3:0] ? rowcount_2 : _GEN_254; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_256 = 4'h3 == _T_91[3:0] ? rowcount_3 : _GEN_255; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_257 = 4'h4 == _T_91[3:0] ? rowcount_4 : _GEN_256; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_258 = 4'h5 == _T_91[3:0] ? rowcount_5 : _GEN_257; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_259 = 4'h6 == _T_91[3:0] ? rowcount_6 : _GEN_258; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_260 = 4'h7 == _T_91[3:0] ? rowcount_7 : _GEN_259; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_261 = 4'h8 == _T_91[3:0] ? rowcount_8 : _GEN_260; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_262 = 4'h9 == _T_91[3:0] ? rowcount_9 : _GEN_261; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_263 = 4'ha == _T_91[3:0] ? rowcount_10 : _GEN_262; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_264 = 4'hb == _T_91[3:0] ? rowcount_11 : _GEN_263; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_265 = 4'hc == _T_91[3:0] ? rowcount_12 : _GEN_264; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_266 = 4'hd == _T_91[3:0] ? rowcount_13 : _GEN_265; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_267 = 4'he == _T_91[3:0] ? rowcount_14 : _GEN_266; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_268 = 4'hf == _T_91[3:0] ? rowcount_15 : _GEN_267; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_381 = _GEN_268 == 32'h1 ? _T_91[31:0] : 32'h18; // @[ivncontrol4.scala 125:17 224:50 225:21]
  wire [31:0] _GEN_382 = _GEN_268 == 32'h2 ? _T_91[31:0] : _GEN_381; // @[ivncontrol4.scala 220:51 221:21]
  wire [31:0] _GEN_383 = _GEN_268 == 32'h2 ? _T_91[31:0] : 32'h17; // @[ivncontrol4.scala 125:17 220:51 222:21]
  wire [31:0] _GEN_384 = _GEN_268 == 32'h3 ? _T_91[31:0] : _GEN_382; // @[ivncontrol4.scala 215:50 216:21]
  wire [31:0] _GEN_385 = _GEN_268 == 32'h3 ? _T_91[31:0] : _GEN_383; // @[ivncontrol4.scala 215:50 217:21]
  wire [31:0] _GEN_386 = _GEN_268 == 32'h3 ? _T_91[31:0] : 32'h5; // @[ivncontrol4.scala 125:17 215:50 218:21]
  wire [31:0] _GEN_387 = _GEN_268 == 32'h4 ? _T_91[31:0] : _GEN_384; // @[ivncontrol4.scala 207:50 208:21]
  wire [31:0] _GEN_388 = _GEN_268 == 32'h4 ? _T_91[31:0] : _GEN_385; // @[ivncontrol4.scala 207:50 209:21]
  wire [31:0] _GEN_389 = _GEN_268 == 32'h4 ? _T_91[31:0] : _GEN_386; // @[ivncontrol4.scala 207:50 210:21]
  wire [31:0] _GEN_390 = _GEN_268 == 32'h4 ? _T_91[31:0] : 32'h17; // @[ivncontrol4.scala 125:17 207:50 211:21]
  wire [31:0] _GEN_391 = _GEN_268 == 32'h5 ? _T_91[31:0] : _GEN_387; // @[ivncontrol4.scala 200:50 201:21]
  wire [31:0] _GEN_392 = _GEN_268 == 32'h5 ? _T_91[31:0] : _GEN_388; // @[ivncontrol4.scala 200:50 202:21]
  wire [31:0] _GEN_393 = _GEN_268 == 32'h5 ? _T_91[31:0] : _GEN_389; // @[ivncontrol4.scala 200:50 203:21]
  wire [31:0] _GEN_394 = _GEN_268 == 32'h5 ? _T_91[31:0] : _GEN_390; // @[ivncontrol4.scala 200:50 204:21]
  wire [31:0] _GEN_395 = _GEN_268 == 32'h5 ? _T_91[31:0] : 32'h2; // @[ivncontrol4.scala 126:18 200:50 205:22]
  wire [31:0] _GEN_396 = _GEN_268 == 32'h6 ? _T_91[31:0] : _GEN_391; // @[ivncontrol4.scala 192:52 193:21]
  wire [31:0] _GEN_397 = _GEN_268 == 32'h6 ? _T_91[31:0] : _GEN_392; // @[ivncontrol4.scala 192:52 194:21]
  wire [31:0] _GEN_398 = _GEN_268 == 32'h6 ? _T_91[31:0] : _GEN_393; // @[ivncontrol4.scala 192:52 195:21]
  wire [31:0] _GEN_399 = _GEN_268 == 32'h6 ? _T_91[31:0] : _GEN_394; // @[ivncontrol4.scala 192:52 196:21]
  wire [31:0] _GEN_400 = _GEN_268 == 32'h6 ? _T_91[31:0] : _GEN_395; // @[ivncontrol4.scala 192:52 197:22]
  wire [31:0] _GEN_401 = _GEN_268 == 32'h6 ? _T_91[31:0] : 32'h11; // @[ivncontrol4.scala 126:18 192:52 198:22]
  wire [31:0] _GEN_402 = _GEN_268 == 32'h7 ? _T_91[31:0] : _GEN_396; // @[ivncontrol4.scala 184:52 185:21]
  wire [31:0] _GEN_403 = _GEN_268 == 32'h7 ? _T_91[31:0] : _GEN_397; // @[ivncontrol4.scala 184:52 186:21]
  wire [31:0] _GEN_404 = _GEN_268 == 32'h7 ? _T_91[31:0] : _GEN_398; // @[ivncontrol4.scala 184:52 187:21]
  wire [31:0] _GEN_405 = _GEN_268 == 32'h7 ? _T_91[31:0] : _GEN_399; // @[ivncontrol4.scala 184:52 188:21]
  wire [31:0] _GEN_406 = _GEN_268 == 32'h7 ? _T_91[31:0] : _GEN_400; // @[ivncontrol4.scala 184:52 189:22]
  wire [31:0] _GEN_407 = _GEN_268 == 32'h7 ? _T_91[31:0] : _GEN_401; // @[ivncontrol4.scala 184:52 190:22]
  wire [31:0] _GEN_408 = _GEN_268 == 32'h7 ? _T_91[31:0] : 32'h16; // @[ivncontrol4.scala 126:18 184:52 191:22]
  wire [31:0] _GEN_409 = _GEN_268 >= 32'h8 ? _T_91[31:0] : _GEN_402; // @[ivncontrol4.scala 174:42 175:21]
  wire [31:0] _GEN_410 = _GEN_268 >= 32'h8 ? _T_91[31:0] : _GEN_403; // @[ivncontrol4.scala 174:42 176:21]
  wire [31:0] _GEN_411 = _GEN_268 >= 32'h8 ? _T_91[31:0] : _GEN_404; // @[ivncontrol4.scala 174:42 177:21]
  wire [31:0] _GEN_412 = _GEN_268 >= 32'h8 ? _T_91[31:0] : _GEN_405; // @[ivncontrol4.scala 174:42 178:21]
  wire [31:0] _GEN_413 = _GEN_268 >= 32'h8 ? _T_91[31:0] : _GEN_406; // @[ivncontrol4.scala 174:42 179:22]
  wire [31:0] _GEN_414 = _GEN_268 >= 32'h8 ? _T_91[31:0] : _GEN_407; // @[ivncontrol4.scala 174:42 180:22]
  wire [31:0] _GEN_415 = _GEN_268 >= 32'h8 ? _T_91[31:0] : _GEN_408; // @[ivncontrol4.scala 174:42 181:22]
  wire [31:0] _GEN_416 = _GEN_268 >= 32'h8 ? _T_91[31:0] : 32'h1d; // @[ivncontrol4.scala 126:18 174:42 182:22]
  wire [31:0] _T_127 = 32'h8 - _GEN_268; // @[ivncontrol4.scala 228:18]
  wire [31:0] _i_vn_1_T_15 = 32'h1 + pin; // @[ivncontrol4.scala 229:29]
  wire [31:0] _GEN_529 = _T_127 == 32'h1 ? _i_vn_1_T_15 : _GEN_416; // @[ivncontrol4.scala 269:54 272:22]
  wire [31:0] _GEN_530 = _T_127 == 32'h2 ? _i_vn_1_T_15 : _GEN_415; // @[ivncontrol4.scala 264:54 267:22]
  wire [31:0] _GEN_531 = _T_127 == 32'h2 ? _i_vn_1_T_15 : _GEN_529; // @[ivncontrol4.scala 264:54 268:22]
  wire [31:0] _GEN_532 = _T_127 == 32'h3 ? _i_vn_1_T_15 : _GEN_414; // @[ivncontrol4.scala 257:54 259:22]
  wire [31:0] _GEN_533 = _T_127 == 32'h3 ? _i_vn_1_T_15 : _GEN_530; // @[ivncontrol4.scala 257:54 260:22]
  wire [31:0] _GEN_534 = _T_127 == 32'h3 ? _i_vn_1_T_15 : _GEN_531; // @[ivncontrol4.scala 257:54 261:22]
  wire [31:0] _GEN_535 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_413; // @[ivncontrol4.scala 251:54 253:22]
  wire [31:0] _GEN_536 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_532; // @[ivncontrol4.scala 251:54 254:22]
  wire [31:0] _GEN_537 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_533; // @[ivncontrol4.scala 251:54 255:22]
  wire [31:0] _GEN_538 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_534; // @[ivncontrol4.scala 251:54 256:22]
  wire [31:0] _GEN_539 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_412; // @[ivncontrol4.scala 244:54 246:21]
  wire [31:0] _GEN_540 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_535; // @[ivncontrol4.scala 244:54 247:22]
  wire [31:0] _GEN_541 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_536; // @[ivncontrol4.scala 244:54 248:22]
  wire [31:0] _GEN_542 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_537; // @[ivncontrol4.scala 244:54 249:22]
  wire [31:0] _GEN_543 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_538; // @[ivncontrol4.scala 244:54 250:22]
  wire [31:0] _GEN_544 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_411; // @[ivncontrol4.scala 237:54 238:22]
  wire [31:0] _GEN_545 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_539; // @[ivncontrol4.scala 237:54 239:21]
  wire [31:0] _GEN_546 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_540; // @[ivncontrol4.scala 237:54 240:22]
  wire [31:0] _GEN_547 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_541; // @[ivncontrol4.scala 237:54 241:22]
  wire [31:0] _GEN_548 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_542; // @[ivncontrol4.scala 237:54 242:22]
  wire [31:0] _GEN_549 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_543; // @[ivncontrol4.scala 237:54 243:22]
  wire [31:0] _GEN_550 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_410; // @[ivncontrol4.scala 228:49 229:22]
  wire [31:0] _GEN_551 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_544; // @[ivncontrol4.scala 228:49 230:21]
  wire [31:0] _GEN_552 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_545; // @[ivncontrol4.scala 228:49 231:21]
  wire [31:0] _GEN_553 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_546; // @[ivncontrol4.scala 228:49 232:22]
  wire [31:0] _GEN_554 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_547; // @[ivncontrol4.scala 228:49 233:22]
  wire [31:0] _GEN_555 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_548; // @[ivncontrol4.scala 228:49 234:22]
  wire [31:0] _GEN_556 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_549; // @[ivncontrol4.scala 228:49 235:22]
  wire [31:0] _GEN_574 = 4'h1 == _i_vn_1_T_15[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_575 = 4'h2 == _i_vn_1_T_15[3:0] ? rowcount_2 : _GEN_574; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_576 = 4'h3 == _i_vn_1_T_15[3:0] ? rowcount_3 : _GEN_575; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_577 = 4'h4 == _i_vn_1_T_15[3:0] ? rowcount_4 : _GEN_576; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_578 = 4'h5 == _i_vn_1_T_15[3:0] ? rowcount_5 : _GEN_577; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_579 = 4'h6 == _i_vn_1_T_15[3:0] ? rowcount_6 : _GEN_578; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_580 = 4'h7 == _i_vn_1_T_15[3:0] ? rowcount_7 : _GEN_579; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_581 = 4'h8 == _i_vn_1_T_15[3:0] ? rowcount_8 : _GEN_580; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_582 = 4'h9 == _i_vn_1_T_15[3:0] ? rowcount_9 : _GEN_581; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_583 = 4'ha == _i_vn_1_T_15[3:0] ? rowcount_10 : _GEN_582; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_584 = 4'hb == _i_vn_1_T_15[3:0] ? rowcount_11 : _GEN_583; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_585 = 4'hc == _i_vn_1_T_15[3:0] ? rowcount_12 : _GEN_584; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_586 = 4'hd == _i_vn_1_T_15[3:0] ? rowcount_13 : _GEN_585; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_587 = 4'he == _i_vn_1_T_15[3:0] ? rowcount_14 : _GEN_586; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_588 = 4'hf == _i_vn_1_T_15[3:0] ? rowcount_15 : _GEN_587; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _T_172 = _GEN_268 + _GEN_588; // @[ivncontrol4.scala 275:41]
  wire [31:0] _T_174 = 32'h8 - _T_172; // @[ivncontrol4.scala 275:18]
  wire [31:0] _i_vn_1_T_17 = 32'h2 + pin; // @[ivncontrol4.scala 276:29]
  wire [31:0] _GEN_781 = _T_174 == 32'h1 ? _i_vn_1_T_17 : _GEN_556; // @[ivncontrol4.scala 318:78 321:22]
  wire [31:0] _GEN_782 = _T_174 == 32'h2 ? _i_vn_1_T_17 : _GEN_555; // @[ivncontrol4.scala 312:76 315:22]
  wire [31:0] _GEN_783 = _T_174 == 32'h2 ? _i_vn_1_T_17 : _GEN_781; // @[ivncontrol4.scala 312:76 316:22]
  wire [31:0] _GEN_784 = _T_174 == 32'h3 ? _i_vn_1_T_17 : _GEN_554; // @[ivncontrol4.scala 305:78 307:23]
  wire [31:0] _GEN_785 = _T_174 == 32'h3 ? _i_vn_1_T_17 : _GEN_782; // @[ivncontrol4.scala 305:78 308:22]
  wire [31:0] _GEN_786 = _T_174 == 32'h3 ? _i_vn_1_T_17 : _GEN_783; // @[ivncontrol4.scala 305:78 309:22]
  wire [31:0] _GEN_787 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_553; // @[ivncontrol4.scala 299:78 301:22]
  wire [31:0] _GEN_788 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_784; // @[ivncontrol4.scala 299:78 302:22]
  wire [31:0] _GEN_789 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_785; // @[ivncontrol4.scala 299:78 303:22]
  wire [31:0] _GEN_790 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_786; // @[ivncontrol4.scala 299:78 304:22]
  wire [31:0] _GEN_791 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_552; // @[ivncontrol4.scala 292:76 294:23]
  wire [31:0] _GEN_792 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_787; // @[ivncontrol4.scala 292:76 295:22]
  wire [31:0] _GEN_793 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_788; // @[ivncontrol4.scala 292:76 296:22]
  wire [31:0] _GEN_794 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_789; // @[ivncontrol4.scala 292:76 297:22]
  wire [31:0] _GEN_795 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_790; // @[ivncontrol4.scala 292:76 298:22]
  wire [31:0] _GEN_796 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_551; // @[ivncontrol4.scala 284:77 286:22]
  wire [31:0] _GEN_797 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_791; // @[ivncontrol4.scala 284:77 287:21]
  wire [31:0] _GEN_798 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_792; // @[ivncontrol4.scala 284:77 288:22]
  wire [31:0] _GEN_799 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_793; // @[ivncontrol4.scala 284:77 289:22]
  wire [31:0] _GEN_800 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_794; // @[ivncontrol4.scala 284:77 290:22]
  wire [31:0] _GEN_801 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_795; // @[ivncontrol4.scala 284:77 291:22]
  wire [31:0] _GEN_802 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_550; // @[ivncontrol4.scala 275:73 276:22]
  wire [31:0] _GEN_803 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_796; // @[ivncontrol4.scala 275:73 277:21]
  wire [31:0] _GEN_804 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_797; // @[ivncontrol4.scala 275:73 278:21]
  wire [31:0] _GEN_805 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_798; // @[ivncontrol4.scala 275:73 279:22]
  wire [31:0] _GEN_806 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_799; // @[ivncontrol4.scala 275:73 280:22]
  wire [31:0] _GEN_807 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_800; // @[ivncontrol4.scala 275:73 281:22]
  wire [31:0] _GEN_808 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_801; // @[ivncontrol4.scala 275:73 282:22]
  wire [31:0] _GEN_842 = 4'h1 == _i_vn_1_T_17[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_843 = 4'h2 == _i_vn_1_T_17[3:0] ? rowcount_2 : _GEN_842; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_844 = 4'h3 == _i_vn_1_T_17[3:0] ? rowcount_3 : _GEN_843; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_845 = 4'h4 == _i_vn_1_T_17[3:0] ? rowcount_4 : _GEN_844; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_846 = 4'h5 == _i_vn_1_T_17[3:0] ? rowcount_5 : _GEN_845; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_847 = 4'h6 == _i_vn_1_T_17[3:0] ? rowcount_6 : _GEN_846; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_848 = 4'h7 == _i_vn_1_T_17[3:0] ? rowcount_7 : _GEN_847; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_849 = 4'h8 == _i_vn_1_T_17[3:0] ? rowcount_8 : _GEN_848; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_850 = 4'h9 == _i_vn_1_T_17[3:0] ? rowcount_9 : _GEN_849; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_851 = 4'ha == _i_vn_1_T_17[3:0] ? rowcount_10 : _GEN_850; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_852 = 4'hb == _i_vn_1_T_17[3:0] ? rowcount_11 : _GEN_851; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_853 = 4'hc == _i_vn_1_T_17[3:0] ? rowcount_12 : _GEN_852; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_854 = 4'hd == _i_vn_1_T_17[3:0] ? rowcount_13 : _GEN_853; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_855 = 4'he == _i_vn_1_T_17[3:0] ? rowcount_14 : _GEN_854; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_856 = 4'hf == _i_vn_1_T_17[3:0] ? rowcount_15 : _GEN_855; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _T_254 = _T_172 + _GEN_856; // @[ivncontrol4.scala 326:62]
  wire [31:0] _T_256 = 32'h8 - _T_254; // @[ivncontrol4.scala 326:17]
  wire [31:0] _i_vn_1_T_19 = 32'h3 + pin; // @[ivncontrol4.scala 327:29]
  wire [31:0] _GEN_1145 = _T_256 == 32'h1 ? _i_vn_1_T_19 : _GEN_808; // @[ivncontrol4.scala 369:100 372:22]
  wire [31:0] _GEN_1146 = _T_256 == 32'h2 ? _i_vn_1_T_19 : _GEN_807; // @[ivncontrol4.scala 363:98 366:22]
  wire [31:0] _GEN_1147 = _T_256 == 32'h2 ? _i_vn_1_T_19 : _GEN_1145; // @[ivncontrol4.scala 363:98 367:22]
  wire [31:0] _GEN_1148 = _T_256 == 32'h3 ? _i_vn_1_T_19 : _GEN_806; // @[ivncontrol4.scala 356:100 358:23]
  wire [31:0] _GEN_1149 = _T_256 == 32'h3 ? _i_vn_1_T_19 : _GEN_1146; // @[ivncontrol4.scala 356:100 359:22]
  wire [31:0] _GEN_1150 = _T_256 == 32'h3 ? _i_vn_1_T_19 : _GEN_1147; // @[ivncontrol4.scala 356:100 360:22]
  wire [31:0] _GEN_1151 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_805; // @[ivncontrol4.scala 350:100 352:22]
  wire [31:0] _GEN_1152 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_1148; // @[ivncontrol4.scala 350:100 353:22]
  wire [31:0] _GEN_1153 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_1149; // @[ivncontrol4.scala 350:100 354:22]
  wire [31:0] _GEN_1154 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_1150; // @[ivncontrol4.scala 350:100 355:22]
  wire [31:0] _GEN_1155 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_804; // @[ivncontrol4.scala 343:98 345:23]
  wire [31:0] _GEN_1156 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1151; // @[ivncontrol4.scala 343:98 346:22]
  wire [31:0] _GEN_1157 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1152; // @[ivncontrol4.scala 343:98 347:22]
  wire [31:0] _GEN_1158 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1153; // @[ivncontrol4.scala 343:98 348:22]
  wire [31:0] _GEN_1159 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1154; // @[ivncontrol4.scala 343:98 349:22]
  wire [31:0] _GEN_1160 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_803; // @[ivncontrol4.scala 335:99 337:22]
  wire [31:0] _GEN_1161 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1155; // @[ivncontrol4.scala 335:99 338:21]
  wire [31:0] _GEN_1162 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1156; // @[ivncontrol4.scala 335:99 339:22]
  wire [31:0] _GEN_1163 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1157; // @[ivncontrol4.scala 335:99 340:22]
  wire [31:0] _GEN_1164 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1158; // @[ivncontrol4.scala 335:99 341:22]
  wire [31:0] _GEN_1165 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1159; // @[ivncontrol4.scala 335:99 342:22]
  wire [31:0] _GEN_1166 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_802; // @[ivncontrol4.scala 326:94 327:22]
  wire [31:0] _GEN_1167 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1160; // @[ivncontrol4.scala 326:94 328:21]
  wire [31:0] _GEN_1168 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1161; // @[ivncontrol4.scala 326:94 329:21]
  wire [31:0] _GEN_1169 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1162; // @[ivncontrol4.scala 326:94 330:22]
  wire [31:0] _GEN_1170 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1163; // @[ivncontrol4.scala 326:94 331:22]
  wire [31:0] _GEN_1171 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1164; // @[ivncontrol4.scala 326:94 332:22]
  wire [31:0] _GEN_1172 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1165; // @[ivncontrol4.scala 326:94 333:22]
  wire [31:0] _GEN_1222 = 4'h1 == _i_vn_1_T_19[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1223 = 4'h2 == _i_vn_1_T_19[3:0] ? rowcount_2 : _GEN_1222; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1224 = 4'h3 == _i_vn_1_T_19[3:0] ? rowcount_3 : _GEN_1223; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1225 = 4'h4 == _i_vn_1_T_19[3:0] ? rowcount_4 : _GEN_1224; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1226 = 4'h5 == _i_vn_1_T_19[3:0] ? rowcount_5 : _GEN_1225; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1227 = 4'h6 == _i_vn_1_T_19[3:0] ? rowcount_6 : _GEN_1226; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1228 = 4'h7 == _i_vn_1_T_19[3:0] ? rowcount_7 : _GEN_1227; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1229 = 4'h8 == _i_vn_1_T_19[3:0] ? rowcount_8 : _GEN_1228; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1230 = 4'h9 == _i_vn_1_T_19[3:0] ? rowcount_9 : _GEN_1229; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1231 = 4'ha == _i_vn_1_T_19[3:0] ? rowcount_10 : _GEN_1230; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1232 = 4'hb == _i_vn_1_T_19[3:0] ? rowcount_11 : _GEN_1231; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1233 = 4'hc == _i_vn_1_T_19[3:0] ? rowcount_12 : _GEN_1232; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1234 = 4'hd == _i_vn_1_T_19[3:0] ? rowcount_13 : _GEN_1233; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1235 = 4'he == _i_vn_1_T_19[3:0] ? rowcount_14 : _GEN_1234; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1236 = 4'hf == _i_vn_1_T_19[3:0] ? rowcount_15 : _GEN_1235; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _T_371 = _T_254 + _GEN_1236; // @[ivncontrol4.scala 376:86]
  wire [31:0] _T_373 = 32'h8 - _T_371; // @[ivncontrol4.scala 376:19]
  wire [31:0] _i_vn_1_T_21 = 32'h4 + pin; // @[ivncontrol4.scala 377:29]
  wire [31:0] _GEN_1621 = _T_373 == 32'h1 ? _i_vn_1_T_21 : _GEN_1172; // @[ivncontrol4.scala 419:122 422:22]
  wire [31:0] _GEN_1622 = _T_373 == 32'h2 ? _i_vn_1_T_21 : _GEN_1171; // @[ivncontrol4.scala 413:121 416:22]
  wire [31:0] _GEN_1623 = _T_373 == 32'h2 ? _i_vn_1_T_21 : _GEN_1621; // @[ivncontrol4.scala 413:121 417:22]
  wire [31:0] _GEN_1624 = _T_373 == 32'h3 ? _i_vn_1_T_21 : _GEN_1170; // @[ivncontrol4.scala 406:123 408:23]
  wire [31:0] _GEN_1625 = _T_373 == 32'h3 ? _i_vn_1_T_21 : _GEN_1622; // @[ivncontrol4.scala 406:123 409:22]
  wire [31:0] _GEN_1626 = _T_373 == 32'h3 ? _i_vn_1_T_21 : _GEN_1623; // @[ivncontrol4.scala 406:123 410:22]
  wire [31:0] _GEN_1627 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1169; // @[ivncontrol4.scala 400:122 402:22]
  wire [31:0] _GEN_1628 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1624; // @[ivncontrol4.scala 400:122 403:22]
  wire [31:0] _GEN_1629 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1625; // @[ivncontrol4.scala 400:122 404:22]
  wire [31:0] _GEN_1630 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1626; // @[ivncontrol4.scala 400:122 405:22]
  wire [31:0] _GEN_1631 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1168; // @[ivncontrol4.scala 393:121 395:23]
  wire [31:0] _GEN_1632 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1627; // @[ivncontrol4.scala 393:121 396:22]
  wire [31:0] _GEN_1633 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1628; // @[ivncontrol4.scala 393:121 397:22]
  wire [31:0] _GEN_1634 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1629; // @[ivncontrol4.scala 393:121 398:22]
  wire [31:0] _GEN_1635 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1630; // @[ivncontrol4.scala 393:121 399:22]
  wire [31:0] _GEN_1636 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1167; // @[ivncontrol4.scala 385:121 387:22]
  wire [31:0] _GEN_1637 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1631; // @[ivncontrol4.scala 385:121 388:21]
  wire [31:0] _GEN_1638 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1632; // @[ivncontrol4.scala 385:121 389:22]
  wire [31:0] _GEN_1639 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1633; // @[ivncontrol4.scala 385:121 390:22]
  wire [31:0] _GEN_1640 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1634; // @[ivncontrol4.scala 385:121 391:22]
  wire [31:0] _GEN_1641 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1635; // @[ivncontrol4.scala 385:121 392:22]
  wire [31:0] _GEN_1642 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1166; // @[ivncontrol4.scala 376:118 377:22]
  wire [31:0] _GEN_1643 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1636; // @[ivncontrol4.scala 376:118 378:21]
  wire [31:0] _GEN_1644 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1637; // @[ivncontrol4.scala 376:118 379:21]
  wire [31:0] _GEN_1645 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1638; // @[ivncontrol4.scala 376:118 380:22]
  wire [31:0] _GEN_1646 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1639; // @[ivncontrol4.scala 376:118 381:22]
  wire [31:0] _GEN_1647 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1640; // @[ivncontrol4.scala 376:118 382:22]
  wire [31:0] _GEN_1648 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1641; // @[ivncontrol4.scala 376:118 383:22]
  wire [31:0] _GEN_1714 = 4'h1 == _i_vn_1_T_21[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1715 = 4'h2 == _i_vn_1_T_21[3:0] ? rowcount_2 : _GEN_1714; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1716 = 4'h3 == _i_vn_1_T_21[3:0] ? rowcount_3 : _GEN_1715; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1717 = 4'h4 == _i_vn_1_T_21[3:0] ? rowcount_4 : _GEN_1716; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1718 = 4'h5 == _i_vn_1_T_21[3:0] ? rowcount_5 : _GEN_1717; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1719 = 4'h6 == _i_vn_1_T_21[3:0] ? rowcount_6 : _GEN_1718; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1720 = 4'h7 == _i_vn_1_T_21[3:0] ? rowcount_7 : _GEN_1719; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1721 = 4'h8 == _i_vn_1_T_21[3:0] ? rowcount_8 : _GEN_1720; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1722 = 4'h9 == _i_vn_1_T_21[3:0] ? rowcount_9 : _GEN_1721; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1723 = 4'ha == _i_vn_1_T_21[3:0] ? rowcount_10 : _GEN_1722; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1724 = 4'hb == _i_vn_1_T_21[3:0] ? rowcount_11 : _GEN_1723; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1725 = 4'hc == _i_vn_1_T_21[3:0] ? rowcount_12 : _GEN_1724; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1726 = 4'hd == _i_vn_1_T_21[3:0] ? rowcount_13 : _GEN_1725; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1727 = 4'he == _i_vn_1_T_21[3:0] ? rowcount_14 : _GEN_1726; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1728 = 4'hf == _i_vn_1_T_21[3:0] ? rowcount_15 : _GEN_1727; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _T_523 = _T_371 + _GEN_1728; // @[ivncontrol4.scala 426:108]
  wire [31:0] _T_525 = 32'h8 - _T_523; // @[ivncontrol4.scala 426:19]
  wire [31:0] _i_vn_1_T_23 = 32'h5 + pin; // @[ivncontrol4.scala 427:29]
  wire [31:0] _GEN_2209 = _T_525 == 32'h1 ? _i_vn_1_T_23 : _GEN_1648; // @[ivncontrol4.scala 469:144 472:22]
  wire [31:0] _GEN_2210 = _T_525 == 32'h2 ? _i_vn_1_T_23 : _GEN_1647; // @[ivncontrol4.scala 463:143 466:22]
  wire [31:0] _GEN_2211 = _T_525 == 32'h2 ? _i_vn_1_T_23 : _GEN_2209; // @[ivncontrol4.scala 463:143 467:22]
  wire [31:0] _GEN_2212 = _T_525 == 32'h3 ? _i_vn_1_T_23 : _GEN_1646; // @[ivncontrol4.scala 456:145 458:23]
  wire [31:0] _GEN_2213 = _T_525 == 32'h3 ? _i_vn_1_T_23 : _GEN_2210; // @[ivncontrol4.scala 456:145 459:22]
  wire [31:0] _GEN_2214 = _T_525 == 32'h3 ? _i_vn_1_T_23 : _GEN_2211; // @[ivncontrol4.scala 456:145 460:22]
  wire [31:0] _GEN_2215 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_1645; // @[ivncontrol4.scala 450:143 452:22]
  wire [31:0] _GEN_2216 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_2212; // @[ivncontrol4.scala 450:143 453:22]
  wire [31:0] _GEN_2217 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_2213; // @[ivncontrol4.scala 450:143 454:22]
  wire [31:0] _GEN_2218 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_2214; // @[ivncontrol4.scala 450:143 455:22]
  wire [31:0] _GEN_2219 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_1644; // @[ivncontrol4.scala 443:143 445:23]
  wire [31:0] _GEN_2220 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2215; // @[ivncontrol4.scala 443:143 446:22]
  wire [31:0] _GEN_2221 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2216; // @[ivncontrol4.scala 443:143 447:22]
  wire [31:0] _GEN_2222 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2217; // @[ivncontrol4.scala 443:143 448:22]
  wire [31:0] _GEN_2223 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2218; // @[ivncontrol4.scala 443:143 449:22]
  wire [31:0] _GEN_2224 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_1643; // @[ivncontrol4.scala 435:143 437:22]
  wire [31:0] _GEN_2225 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2219; // @[ivncontrol4.scala 435:143 438:21]
  wire [31:0] _GEN_2226 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2220; // @[ivncontrol4.scala 435:143 439:22]
  wire [31:0] _GEN_2227 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2221; // @[ivncontrol4.scala 435:143 440:22]
  wire [31:0] _GEN_2228 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2222; // @[ivncontrol4.scala 435:143 441:22]
  wire [31:0] _GEN_2229 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2223; // @[ivncontrol4.scala 435:143 442:22]
  wire [31:0] _GEN_2230 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_1642; // @[ivncontrol4.scala 426:140 427:22]
  wire [31:0] _GEN_2231 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2224; // @[ivncontrol4.scala 426:140 428:21]
  wire [31:0] _GEN_2232 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2225; // @[ivncontrol4.scala 426:140 429:21]
  wire [31:0] _GEN_2233 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2226; // @[ivncontrol4.scala 426:140 430:22]
  wire [31:0] _GEN_2234 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2227; // @[ivncontrol4.scala 426:140 431:22]
  wire [31:0] _GEN_2235 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2228; // @[ivncontrol4.scala 426:140 432:22]
  wire [31:0] _GEN_2236 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2229; // @[ivncontrol4.scala 426:140 433:22]
  wire [31:0] _GEN_2318 = 4'h1 == _i_vn_1_T_23[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2319 = 4'h2 == _i_vn_1_T_23[3:0] ? rowcount_2 : _GEN_2318; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2320 = 4'h3 == _i_vn_1_T_23[3:0] ? rowcount_3 : _GEN_2319; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2321 = 4'h4 == _i_vn_1_T_23[3:0] ? rowcount_4 : _GEN_2320; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2322 = 4'h5 == _i_vn_1_T_23[3:0] ? rowcount_5 : _GEN_2321; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2323 = 4'h6 == _i_vn_1_T_23[3:0] ? rowcount_6 : _GEN_2322; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2324 = 4'h7 == _i_vn_1_T_23[3:0] ? rowcount_7 : _GEN_2323; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2325 = 4'h8 == _i_vn_1_T_23[3:0] ? rowcount_8 : _GEN_2324; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2326 = 4'h9 == _i_vn_1_T_23[3:0] ? rowcount_9 : _GEN_2325; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2327 = 4'ha == _i_vn_1_T_23[3:0] ? rowcount_10 : _GEN_2326; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2328 = 4'hb == _i_vn_1_T_23[3:0] ? rowcount_11 : _GEN_2327; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2329 = 4'hc == _i_vn_1_T_23[3:0] ? rowcount_12 : _GEN_2328; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2330 = 4'hd == _i_vn_1_T_23[3:0] ? rowcount_13 : _GEN_2329; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2331 = 4'he == _i_vn_1_T_23[3:0] ? rowcount_14 : _GEN_2330; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2332 = 4'hf == _i_vn_1_T_23[3:0] ? rowcount_15 : _GEN_2331; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _T_710 = _T_523 + _GEN_2332; // @[ivncontrol4.scala 477:130]
  wire [31:0] _T_712 = 32'h8 - _T_710; // @[ivncontrol4.scala 477:19]
  wire [31:0] _i_vn_1_T_25 = 32'h6 + pin; // @[ivncontrol4.scala 478:29]
  wire [31:0] _GEN_2909 = _T_712 == 32'h1 ? _i_vn_1_T_25 : _GEN_2236; // @[ivncontrol4.scala 520:166 523:22]
  wire [31:0] _GEN_2910 = _T_712 == 32'h2 ? _i_vn_1_T_25 : _GEN_2235; // @[ivncontrol4.scala 514:166 517:22]
  wire [31:0] _GEN_2911 = _T_712 == 32'h2 ? _i_vn_1_T_25 : _GEN_2909; // @[ivncontrol4.scala 514:166 518:22]
  wire [31:0] _GEN_2912 = _T_712 == 32'h3 ? _i_vn_1_T_25 : _GEN_2234; // @[ivncontrol4.scala 507:168 509:23]
  wire [31:0] _GEN_2913 = _T_712 == 32'h3 ? _i_vn_1_T_25 : _GEN_2910; // @[ivncontrol4.scala 507:168 510:22]
  wire [31:0] _GEN_2914 = _T_712 == 32'h3 ? _i_vn_1_T_25 : _GEN_2911; // @[ivncontrol4.scala 507:168 511:22]
  wire [31:0] _GEN_2915 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2233; // @[ivncontrol4.scala 501:166 503:22]
  wire [31:0] _GEN_2916 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2912; // @[ivncontrol4.scala 501:166 504:22]
  wire [31:0] _GEN_2917 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2913; // @[ivncontrol4.scala 501:166 505:22]
  wire [31:0] _GEN_2918 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2914; // @[ivncontrol4.scala 501:166 506:22]
  wire [31:0] _GEN_2919 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2232; // @[ivncontrol4.scala 494:166 496:23]
  wire [31:0] _GEN_2920 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2915; // @[ivncontrol4.scala 494:166 497:22]
  wire [31:0] _GEN_2921 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2916; // @[ivncontrol4.scala 494:166 498:22]
  wire [31:0] _GEN_2922 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2917; // @[ivncontrol4.scala 494:166 499:22]
  wire [31:0] _GEN_2923 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2918; // @[ivncontrol4.scala 494:166 500:22]
  wire [31:0] _GEN_2924 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2231; // @[ivncontrol4.scala 486:166 488:22]
  wire [31:0] _GEN_2925 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2919; // @[ivncontrol4.scala 486:166 489:21]
  wire [31:0] _GEN_2926 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2920; // @[ivncontrol4.scala 486:166 490:22]
  wire [31:0] _GEN_2927 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2921; // @[ivncontrol4.scala 486:166 491:22]
  wire [31:0] _GEN_2928 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2922; // @[ivncontrol4.scala 486:166 492:22]
  wire [31:0] _GEN_2929 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2923; // @[ivncontrol4.scala 486:166 493:22]
  wire [31:0] _GEN_2930 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2230; // @[ivncontrol4.scala 477:162 478:22]
  wire [31:0] _GEN_2931 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2924; // @[ivncontrol4.scala 477:162 479:21]
  wire [31:0] _GEN_2932 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2925; // @[ivncontrol4.scala 477:162 480:21]
  wire [31:0] _GEN_2933 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2926; // @[ivncontrol4.scala 477:162 481:22]
  wire [31:0] _GEN_2934 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2927; // @[ivncontrol4.scala 477:162 482:22]
  wire [31:0] _GEN_2935 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2928; // @[ivncontrol4.scala 477:162 483:22]
  wire [31:0] _GEN_2936 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2929; // @[ivncontrol4.scala 477:162 484:22]
  wire [31:0] _GEN_3034 = 4'h1 == _i_vn_1_T_25[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3035 = 4'h2 == _i_vn_1_T_25[3:0] ? rowcount_2 : _GEN_3034; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3036 = 4'h3 == _i_vn_1_T_25[3:0] ? rowcount_3 : _GEN_3035; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3037 = 4'h4 == _i_vn_1_T_25[3:0] ? rowcount_4 : _GEN_3036; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3038 = 4'h5 == _i_vn_1_T_25[3:0] ? rowcount_5 : _GEN_3037; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3039 = 4'h6 == _i_vn_1_T_25[3:0] ? rowcount_6 : _GEN_3038; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3040 = 4'h7 == _i_vn_1_T_25[3:0] ? rowcount_7 : _GEN_3039; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3041 = 4'h8 == _i_vn_1_T_25[3:0] ? rowcount_8 : _GEN_3040; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3042 = 4'h9 == _i_vn_1_T_25[3:0] ? rowcount_9 : _GEN_3041; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3043 = 4'ha == _i_vn_1_T_25[3:0] ? rowcount_10 : _GEN_3042; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3044 = 4'hb == _i_vn_1_T_25[3:0] ? rowcount_11 : _GEN_3043; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3045 = 4'hc == _i_vn_1_T_25[3:0] ? rowcount_12 : _GEN_3044; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3046 = 4'hd == _i_vn_1_T_25[3:0] ? rowcount_13 : _GEN_3045; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3047 = 4'he == _i_vn_1_T_25[3:0] ? rowcount_14 : _GEN_3046; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3048 = 4'hf == _i_vn_1_T_25[3:0] ? rowcount_15 : _GEN_3047; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _T_932 = _T_710 + _GEN_3048; // @[ivncontrol4.scala 528:152]
  wire [31:0] _T_934 = 32'h8 - _T_932; // @[ivncontrol4.scala 528:19]
  wire [31:0] _i_vn_1_T_27 = 32'h7 + pin; // @[ivncontrol4.scala 529:29]
  wire [31:0] _GEN_3721 = _T_934 == 32'h1 ? _i_vn_1_T_27 : _GEN_2936; // @[ivncontrol4.scala 571:188 574:22]
  wire [31:0] _GEN_3722 = _T_934 == 32'h2 ? _i_vn_1_T_27 : _GEN_2935; // @[ivncontrol4.scala 565:188 568:22]
  wire [31:0] _GEN_3723 = _T_934 == 32'h2 ? _i_vn_1_T_27 : _GEN_3721; // @[ivncontrol4.scala 565:188 569:22]
  wire [31:0] _GEN_3724 = _T_934 == 32'h3 ? _i_vn_1_T_27 : _GEN_2934; // @[ivncontrol4.scala 558:190 560:23]
  wire [31:0] _GEN_3725 = _T_934 == 32'h3 ? _i_vn_1_T_27 : _GEN_3722; // @[ivncontrol4.scala 558:190 561:22]
  wire [31:0] _GEN_3726 = _T_934 == 32'h3 ? _i_vn_1_T_27 : _GEN_3723; // @[ivncontrol4.scala 558:190 562:22]
  wire [31:0] _GEN_3727 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_2933; // @[ivncontrol4.scala 552:188 554:22]
  wire [31:0] _GEN_3728 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_3724; // @[ivncontrol4.scala 552:188 555:22]
  wire [31:0] _GEN_3729 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_3725; // @[ivncontrol4.scala 552:188 556:22]
  wire [31:0] _GEN_3730 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_3726; // @[ivncontrol4.scala 552:188 557:22]
  wire [31:0] _GEN_3731 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_2932; // @[ivncontrol4.scala 545:188 547:23]
  wire [31:0] _GEN_3732 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3727; // @[ivncontrol4.scala 545:188 548:22]
  wire [31:0] _GEN_3733 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3728; // @[ivncontrol4.scala 545:188 549:22]
  wire [31:0] _GEN_3734 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3729; // @[ivncontrol4.scala 545:188 550:22]
  wire [31:0] _GEN_3735 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3730; // @[ivncontrol4.scala 545:188 551:22]
  wire [31:0] _GEN_3736 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_2931; // @[ivncontrol4.scala 537:188 539:22]
  wire [31:0] _GEN_3737 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3731; // @[ivncontrol4.scala 537:188 540:21]
  wire [31:0] _GEN_3738 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3732; // @[ivncontrol4.scala 537:188 541:22]
  wire [31:0] _GEN_3739 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3733; // @[ivncontrol4.scala 537:188 542:22]
  wire [31:0] _GEN_3740 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3734; // @[ivncontrol4.scala 537:188 543:22]
  wire [31:0] _GEN_3741 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3735; // @[ivncontrol4.scala 537:188 544:22]
  wire [31:0] _GEN_3742 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_2930; // @[ivncontrol4.scala 528:184 529:22]
  wire [31:0] _GEN_3743 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3736; // @[ivncontrol4.scala 528:184 530:21]
  wire [31:0] _GEN_3744 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3737; // @[ivncontrol4.scala 528:184 531:21]
  wire [31:0] _GEN_3745 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3738; // @[ivncontrol4.scala 528:184 532:22]
  wire [31:0] _GEN_3746 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3739; // @[ivncontrol4.scala 528:184 533:22]
  wire [31:0] _GEN_3747 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3740; // @[ivncontrol4.scala 528:184 534:22]
  wire [31:0] _GEN_3748 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3741; // @[ivncontrol4.scala 528:184 535:22]
  wire [31:0] _GEN_3749 = _GEN_244 ? _GEN_409 : 32'h18; // @[ivncontrol4.scala 125:17 172:28]
  wire [31:0] _GEN_3750 = _GEN_244 ? _GEN_3742 : 32'h17; // @[ivncontrol4.scala 125:17 172:28]
  wire [31:0] _GEN_3751 = _GEN_244 ? _GEN_3743 : 32'h5; // @[ivncontrol4.scala 125:17 172:28]
  wire [31:0] _GEN_3752 = _GEN_244 ? _GEN_3744 : 32'h17; // @[ivncontrol4.scala 125:17 172:28]
  wire [31:0] _GEN_3753 = _GEN_244 ? _GEN_3745 : 32'h2; // @[ivncontrol4.scala 126:18 172:28]
  wire [31:0] _GEN_3754 = _GEN_244 ? _GEN_3746 : 32'h11; // @[ivncontrol4.scala 126:18 172:28]
  wire [31:0] _GEN_3755 = _GEN_244 ? _GEN_3747 : 32'h16; // @[ivncontrol4.scala 126:18 172:28]
  wire [31:0] _GEN_3756 = _GEN_244 ? _GEN_3748 : 32'h1d; // @[ivncontrol4.scala 126:18 172:28]
  wire [31:0] _GEN_4137 = reset ? 32'h0 : _GEN_3749; // @[ivncontrol4.scala 16:{23,23}]
  wire [31:0] _GEN_4138 = reset ? 32'h0 : _GEN_3750; // @[ivncontrol4.scala 16:{23,23}]
  wire [31:0] _GEN_4139 = reset ? 32'h0 : _GEN_3751; // @[ivncontrol4.scala 16:{23,23}]
  wire [31:0] _GEN_4140 = reset ? 32'h0 : _GEN_3752; // @[ivncontrol4.scala 16:{23,23}]
  wire [31:0] _GEN_4141 = reset ? 32'h0 : _GEN_3753; // @[ivncontrol4.scala 17:{24,24}]
  wire [31:0] _GEN_4142 = reset ? 32'h0 : _GEN_3754; // @[ivncontrol4.scala 17:{24,24}]
  wire [31:0] _GEN_4143 = reset ? 32'h0 : _GEN_3755; // @[ivncontrol4.scala 17:{24,24}]
  wire [31:0] _GEN_4144 = reset ? 32'h0 : _GEN_3756; // @[ivncontrol4.scala 17:{24,24}]
  assign io_o_vn_0 = i_vn_0; // @[ivncontrol4.scala 121:13]
  assign io_o_vn_1 = i_vn_1; // @[ivncontrol4.scala 121:13]
  assign io_o_vn_2 = i_vn_2; // @[ivncontrol4.scala 121:13]
  assign io_o_vn_3 = i_vn_3; // @[ivncontrol4.scala 121:13]
  assign io_o_vn2_0 = i_vn2_0; // @[ivncontrol4.scala 122:14]
  assign io_o_vn2_1 = i_vn2_1; // @[ivncontrol4.scala 122:14]
  assign io_o_vn2_2 = i_vn2_2; // @[ivncontrol4.scala 122:14]
  assign io_o_vn2_3 = i_vn2_3; // @[ivncontrol4.scala 122:14]
  assign io_ProcessValid = _k_T_2 & io_ProcessValid_REG; // @[ivncontrol4.scala 41:36 42:25 44:25]
  always @(posedge clock) begin
    i_vn_0 <= _GEN_4137[4:0]; // @[ivncontrol4.scala 16:{23,23}]
    i_vn_1 <= _GEN_4138[4:0]; // @[ivncontrol4.scala 16:{23,23}]
    i_vn_2 <= _GEN_4139[4:0]; // @[ivncontrol4.scala 16:{23,23}]
    i_vn_3 <= _GEN_4140[4:0]; // @[ivncontrol4.scala 16:{23,23}]
    i_vn2_0 <= _GEN_4141[4:0]; // @[ivncontrol4.scala 17:{24,24}]
    i_vn2_1 <= _GEN_4142[4:0]; // @[ivncontrol4.scala 17:{24,24}]
    i_vn2_2 <= _GEN_4143[4:0]; // @[ivncontrol4.scala 17:{24,24}]
    i_vn2_3 <= _GEN_4144[4:0]; // @[ivncontrol4.scala 17:{24,24}]
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_0 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_0 <= count_0; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_1 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_1 <= count_1; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_2 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_2 <= count_2; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_3 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_3 <= count_3; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_4 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_4 <= count_4; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_5 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_5 <= count_5; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_6 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_6 <= count_6; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_7 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_7 <= count_7; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_8 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_8 <= 32'h0; // @[ivncontrol4.scala 81:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_9 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_9 <= 32'h0; // @[ivncontrol4.scala 81:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_10 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_10 <= 32'h0; // @[ivncontrol4.scala 81:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_11 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_11 <= 32'h0; // @[ivncontrol4.scala 81:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_12 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_12 <= 32'h0; // @[ivncontrol4.scala 81:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_13 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_13 <= 32'h0; // @[ivncontrol4.scala 81:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_14 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_14 <= 32'h0; // @[ivncontrol4.scala 81:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_15 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end
    if (reset) begin // @[ivncontrol4.scala 31:22]
      pin <= 32'h0; // @[ivncontrol4.scala 31:22]
    end else if (_T_72 & rowcount_6 == 32'h0 & rowcount_7 != 32'h0) begin // @[ivncontrol4.scala 166:192]
      pin <= 32'h7; // @[ivncontrol4.scala 167:13]
    end else if (_T_59 & rowcount_5 == 32'h0 & rowcount_6 != 32'h0) begin // @[ivncontrol4.scala 163:169]
      pin <= 32'h6; // @[ivncontrol4.scala 164:13]
    end else if (_T_48 & rowcount_4 == 32'h0 & rowcount_5 != 32'h0) begin // @[ivncontrol4.scala 160:146]
      pin <= 32'h5; // @[ivncontrol4.scala 161:13]
    end else begin
      pin <= _GEN_249;
    end
    if (reset) begin // @[ivncontrol4.scala 35:20]
      i <= 32'h0; // @[ivncontrol4.scala 35:20]
    end else if (i < 32'h7 & _k_T_1) begin // @[ivncontrol4.scala 103:74]
      i <= _i_T_1; // @[ivncontrol4.scala 104:11]
    end
    if (reset) begin // @[ivncontrol4.scala 36:20]
      j <= 32'h0; // @[ivncontrol4.scala 36:20]
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 107:71]
      j <= _j_T_1; // @[ivncontrol4.scala 108:11]
    end else if (!(_k_T_2)) begin // @[ivncontrol4.scala 110:81]
      j <= 32'h0; // @[ivncontrol4.scala 114:11]
    end
    k <= i == 32'h7 & j == 32'h7; // @[ivncontrol4.scala 38:31]
    io_ProcessValid_REG <= k; // @[ivncontrol4.scala 42:35]
    if (3'h0 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h0 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h0 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h0 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h0 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h0 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h0 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h0 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h0 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_0 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h1 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_1 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h2 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_2 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h3 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_3 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h4 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_4 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h5 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_5 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h6 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_6 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h7 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_7 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  i_vn_0 = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  i_vn_1 = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  i_vn_2 = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  i_vn_3 = _RAND_3[4:0];
  _RAND_4 = {1{`RANDOM}};
  i_vn2_0 = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  i_vn2_1 = _RAND_5[4:0];
  _RAND_6 = {1{`RANDOM}};
  i_vn2_2 = _RAND_6[4:0];
  _RAND_7 = {1{`RANDOM}};
  i_vn2_3 = _RAND_7[4:0];
  _RAND_8 = {1{`RANDOM}};
  rowcount_0 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  rowcount_1 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  rowcount_2 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  rowcount_3 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  rowcount_4 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  rowcount_5 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  rowcount_6 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  rowcount_7 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  rowcount_8 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  rowcount_9 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  rowcount_10 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  rowcount_11 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  rowcount_12 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  rowcount_13 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  rowcount_14 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  rowcount_15 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  pin = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  i = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  j = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  k = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  io_ProcessValid_REG = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  mat_0_0 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  mat_0_1 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  mat_0_2 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  mat_0_3 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  mat_0_4 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  mat_0_5 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  mat_0_6 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  mat_0_7 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  mat_1_0 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  mat_1_1 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  mat_1_2 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  mat_1_3 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  mat_1_4 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  mat_1_5 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  mat_1_6 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  mat_1_7 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  mat_2_0 = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  mat_2_1 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  mat_2_2 = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  mat_2_3 = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  mat_2_4 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  mat_2_5 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  mat_2_6 = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  mat_2_7 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  mat_3_0 = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  mat_3_1 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  mat_3_2 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  mat_3_3 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  mat_3_4 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  mat_3_5 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  mat_3_6 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  mat_3_7 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  mat_4_0 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  mat_4_1 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  mat_4_2 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  mat_4_3 = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  mat_4_4 = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  mat_4_5 = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  mat_4_6 = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  mat_4_7 = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  mat_5_0 = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  mat_5_1 = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  mat_5_2 = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  mat_5_3 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  mat_5_4 = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  mat_5_5 = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  mat_5_6 = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  mat_5_7 = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  mat_6_0 = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  mat_6_1 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  mat_6_2 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  mat_6_3 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  mat_6_4 = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  mat_6_5 = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  mat_6_6 = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  mat_6_7 = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  mat_7_0 = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  mat_7_1 = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  mat_7_2 = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  mat_7_3 = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  mat_7_4 = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  mat_7_5 = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  mat_7_6 = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  mat_7_7 = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  count_0 = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  count_1 = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  count_2 = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  count_3 = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  count_4 = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  count_5 = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  count_6 = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  count_7 = _RAND_100[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ivncontrol4_1(
  input         clock,
  input         reset,
  input  [15:0] io_Stationary_matrix_0_0,
  input  [15:0] io_Stationary_matrix_0_1,
  input  [15:0] io_Stationary_matrix_0_2,
  input  [15:0] io_Stationary_matrix_0_3,
  input  [15:0] io_Stationary_matrix_0_4,
  input  [15:0] io_Stationary_matrix_0_5,
  input  [15:0] io_Stationary_matrix_0_6,
  input  [15:0] io_Stationary_matrix_0_7,
  input  [15:0] io_Stationary_matrix_1_0,
  input  [15:0] io_Stationary_matrix_1_1,
  input  [15:0] io_Stationary_matrix_1_2,
  input  [15:0] io_Stationary_matrix_1_3,
  input  [15:0] io_Stationary_matrix_1_4,
  input  [15:0] io_Stationary_matrix_1_5,
  input  [15:0] io_Stationary_matrix_1_6,
  input  [15:0] io_Stationary_matrix_1_7,
  input  [15:0] io_Stationary_matrix_2_0,
  input  [15:0] io_Stationary_matrix_2_1,
  input  [15:0] io_Stationary_matrix_2_2,
  input  [15:0] io_Stationary_matrix_2_3,
  input  [15:0] io_Stationary_matrix_2_4,
  input  [15:0] io_Stationary_matrix_2_5,
  input  [15:0] io_Stationary_matrix_2_6,
  input  [15:0] io_Stationary_matrix_2_7,
  input  [15:0] io_Stationary_matrix_3_0,
  input  [15:0] io_Stationary_matrix_3_1,
  input  [15:0] io_Stationary_matrix_3_2,
  input  [15:0] io_Stationary_matrix_3_3,
  input  [15:0] io_Stationary_matrix_3_4,
  input  [15:0] io_Stationary_matrix_3_5,
  input  [15:0] io_Stationary_matrix_3_6,
  input  [15:0] io_Stationary_matrix_3_7,
  input  [15:0] io_Stationary_matrix_4_0,
  input  [15:0] io_Stationary_matrix_4_1,
  input  [15:0] io_Stationary_matrix_4_2,
  input  [15:0] io_Stationary_matrix_4_3,
  input  [15:0] io_Stationary_matrix_4_4,
  input  [15:0] io_Stationary_matrix_4_5,
  input  [15:0] io_Stationary_matrix_4_6,
  input  [15:0] io_Stationary_matrix_4_7,
  input  [15:0] io_Stationary_matrix_5_0,
  input  [15:0] io_Stationary_matrix_5_1,
  input  [15:0] io_Stationary_matrix_5_2,
  input  [15:0] io_Stationary_matrix_5_3,
  input  [15:0] io_Stationary_matrix_5_4,
  input  [15:0] io_Stationary_matrix_5_5,
  input  [15:0] io_Stationary_matrix_5_6,
  input  [15:0] io_Stationary_matrix_5_7,
  input  [15:0] io_Stationary_matrix_6_0,
  input  [15:0] io_Stationary_matrix_6_1,
  input  [15:0] io_Stationary_matrix_6_2,
  input  [15:0] io_Stationary_matrix_6_3,
  input  [15:0] io_Stationary_matrix_6_4,
  input  [15:0] io_Stationary_matrix_6_5,
  input  [15:0] io_Stationary_matrix_6_6,
  input  [15:0] io_Stationary_matrix_6_7,
  input  [15:0] io_Stationary_matrix_7_0,
  input  [15:0] io_Stationary_matrix_7_1,
  input  [15:0] io_Stationary_matrix_7_2,
  input  [15:0] io_Stationary_matrix_7_3,
  input  [15:0] io_Stationary_matrix_7_4,
  input  [15:0] io_Stationary_matrix_7_5,
  input  [15:0] io_Stationary_matrix_7_6,
  input  [15:0] io_Stationary_matrix_7_7,
  output [4:0]  io_o_vn_0,
  output [4:0]  io_o_vn_1,
  output [4:0]  io_o_vn_2,
  output [4:0]  io_o_vn_3,
  output [4:0]  io_o_vn2_0,
  output [4:0]  io_o_vn2_1,
  output [4:0]  io_o_vn2_2,
  output [4:0]  io_o_vn2_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
`endif // RANDOMIZE_REG_INIT
  reg [4:0] i_vn_0; // @[ivncontrol4.scala 16:23]
  reg [4:0] i_vn_1; // @[ivncontrol4.scala 16:23]
  reg [4:0] i_vn_2; // @[ivncontrol4.scala 16:23]
  reg [4:0] i_vn_3; // @[ivncontrol4.scala 16:23]
  reg [4:0] i_vn2_0; // @[ivncontrol4.scala 17:24]
  reg [4:0] i_vn2_1; // @[ivncontrol4.scala 17:24]
  reg [4:0] i_vn2_2; // @[ivncontrol4.scala 17:24]
  reg [4:0] i_vn2_3; // @[ivncontrol4.scala 17:24]
  reg [31:0] rowcount_0; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_1; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_2; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_3; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_4; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_5; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_6; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_7; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_8; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_9; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_10; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_11; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_12; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_13; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_14; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_15; // @[ivncontrol4.scala 21:27]
  reg [31:0] pin; // @[ivncontrol4.scala 31:22]
  reg [31:0] i; // @[ivncontrol4.scala 35:20]
  reg [31:0] j; // @[ivncontrol4.scala 36:20]
  wire  _k_T_1 = j == 32'h7; // @[ivncontrol4.scala 38:37]
  wire  _k_T_2 = i == 32'h7 & j == 32'h7; // @[ivncontrol4.scala 38:31]
  reg [31:0] mat_0_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_0_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_0_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_0_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_0_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_0_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_0_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_0_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] count_0; // @[ivncontrol4.scala 52:20]
  reg [31:0] count_1; // @[ivncontrol4.scala 52:20]
  reg [31:0] count_2; // @[ivncontrol4.scala 52:20]
  reg [31:0] count_3; // @[ivncontrol4.scala 52:20]
  reg [31:0] count_4; // @[ivncontrol4.scala 52:20]
  reg [31:0] count_5; // @[ivncontrol4.scala 52:20]
  reg [31:0] count_6; // @[ivncontrol4.scala 52:20]
  reg [31:0] count_7; // @[ivncontrol4.scala 52:20]
  wire [15:0] _GEN_66 = 3'h0 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_0_1 : io_Stationary_matrix_0_0; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_67 = 3'h0 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_0_2 : _GEN_66; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_68 = 3'h0 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_0_3 : _GEN_67; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_69 = 3'h0 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_0_4 : _GEN_68; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_70 = 3'h0 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_0_5 : _GEN_69; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_71 = 3'h0 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_0_6 : _GEN_70; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_72 = 3'h0 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_0_7 : _GEN_71; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_73 = 3'h1 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_1_0 : _GEN_72; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_74 = 3'h1 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_1_1 : _GEN_73; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_75 = 3'h1 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_1_2 : _GEN_74; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_76 = 3'h1 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_1_3 : _GEN_75; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_77 = 3'h1 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_1_4 : _GEN_76; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_78 = 3'h1 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_1_5 : _GEN_77; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_79 = 3'h1 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_1_6 : _GEN_78; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_80 = 3'h1 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_1_7 : _GEN_79; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_81 = 3'h2 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_2_0 : _GEN_80; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_82 = 3'h2 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_2_1 : _GEN_81; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_83 = 3'h2 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_2_2 : _GEN_82; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_84 = 3'h2 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_2_3 : _GEN_83; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_85 = 3'h2 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_2_4 : _GEN_84; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_86 = 3'h2 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_2_5 : _GEN_85; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_87 = 3'h2 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_2_6 : _GEN_86; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_88 = 3'h2 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_2_7 : _GEN_87; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_89 = 3'h3 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_3_0 : _GEN_88; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_90 = 3'h3 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_3_1 : _GEN_89; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_91 = 3'h3 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_3_2 : _GEN_90; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_92 = 3'h3 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_3_3 : _GEN_91; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_93 = 3'h3 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_3_4 : _GEN_92; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_94 = 3'h3 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_3_5 : _GEN_93; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_95 = 3'h3 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_3_6 : _GEN_94; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_96 = 3'h3 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_3_7 : _GEN_95; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_97 = 3'h4 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_4_0 : _GEN_96; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_98 = 3'h4 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_4_1 : _GEN_97; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_99 = 3'h4 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_4_2 : _GEN_98; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_100 = 3'h4 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_4_3 : _GEN_99; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_101 = 3'h4 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_4_4 : _GEN_100; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_102 = 3'h4 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_4_5 : _GEN_101; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_103 = 3'h4 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_4_6 : _GEN_102; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_104 = 3'h4 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_4_7 : _GEN_103; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_105 = 3'h5 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_5_0 : _GEN_104; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_106 = 3'h5 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_5_1 : _GEN_105; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_107 = 3'h5 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_5_2 : _GEN_106; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_108 = 3'h5 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_5_3 : _GEN_107; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_109 = 3'h5 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_5_4 : _GEN_108; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_110 = 3'h5 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_5_5 : _GEN_109; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_111 = 3'h5 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_5_6 : _GEN_110; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_112 = 3'h5 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_5_7 : _GEN_111; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_113 = 3'h6 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_6_0 : _GEN_112; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_114 = 3'h6 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_6_1 : _GEN_113; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_115 = 3'h6 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_6_2 : _GEN_114; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_116 = 3'h6 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_6_3 : _GEN_115; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_117 = 3'h6 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_6_4 : _GEN_116; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_118 = 3'h6 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_6_5 : _GEN_117; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_119 = 3'h6 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_6_6 : _GEN_118; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_120 = 3'h6 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_6_7 : _GEN_119; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_121 = 3'h7 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_7_0 : _GEN_120; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_122 = 3'h7 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_7_1 : _GEN_121; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_123 = 3'h7 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_7_2 : _GEN_122; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_124 = 3'h7 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_7_3 : _GEN_123; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_125 = 3'h7 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_7_4 : _GEN_124; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_126 = 3'h7 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_7_5 : _GEN_125; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_127 = 3'h7 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_7_6 : _GEN_126; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_128 = 3'h7 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_7_7 : _GEN_127; // @[ivncontrol4.scala 57:{15,15}]
  wire [31:0] _mat_T_3_T_4 = {{16'd0}, _GEN_128}; // @[ivncontrol4.scala 57:{15,15}]
  wire  _GEN_225 = count_7 >= 32'h8; // @[ivncontrol4.scala 66:28 67:16]
  wire  valid1 = count_7 >= 32'h8; // @[ivncontrol4.scala 66:28 67:16]
  wire [31:0] _GEN_194 = 3'h1 == i[2:0] ? count_1 : count_0; // @[ivncontrol4.scala 60:{33,33}]
  wire [31:0] _GEN_195 = 3'h2 == i[2:0] ? count_2 : _GEN_194; // @[ivncontrol4.scala 60:{33,33}]
  wire [31:0] _GEN_196 = 3'h3 == i[2:0] ? count_3 : _GEN_195; // @[ivncontrol4.scala 60:{33,33}]
  wire [31:0] _GEN_197 = 3'h4 == i[2:0] ? count_4 : _GEN_196; // @[ivncontrol4.scala 60:{33,33}]
  wire [31:0] _GEN_198 = 3'h5 == i[2:0] ? count_5 : _GEN_197; // @[ivncontrol4.scala 60:{33,33}]
  wire [31:0] _GEN_199 = 3'h6 == i[2:0] ? count_6 : _GEN_198; // @[ivncontrol4.scala 60:{33,33}]
  wire [31:0] _GEN_200 = 3'h7 == i[2:0] ? count_7 : _GEN_199; // @[ivncontrol4.scala 60:{33,33}]
  wire [31:0] _count_T_2 = _GEN_200 + 32'h1; // @[ivncontrol4.scala 60:33]
  wire [31:0] _i_T_1 = i + 32'h1; // @[ivncontrol4.scala 104:16]
  wire [31:0] _j_T_1 = j + 32'h1; // @[ivncontrol4.scala 108:16]
  wire  _GEN_244 = _k_T_2; // @[ivncontrol4.scala 136:75 137:14 139:14]
  wire [31:0] _GEN_245 = rowcount_0 != 32'h0 ? 32'h0 : pin; // @[ivncontrol4.scala 145:30 146:13 31:22]
  wire  _T_27 = rowcount_0 == 32'h0; // @[ivncontrol4.scala 148:23]
  wire [31:0] _GEN_246 = rowcount_0 == 32'h0 & rowcount_1 != 32'h0 ? 32'h1 : _GEN_245; // @[ivncontrol4.scala 148:54 149:13]
  wire  _T_32 = _T_27 & rowcount_1 == 32'h0; // @[ivncontrol4.scala 151:31]
  wire [31:0] _GEN_247 = _T_27 & rowcount_1 == 32'h0 & rowcount_2 != 32'h0 ? 32'h2 : _GEN_246; // @[ivncontrol4.scala 151:77 152:13]
  wire  _T_39 = _T_32 & rowcount_2 == 32'h0; // @[ivncontrol4.scala 154:54]
  wire [31:0] _GEN_248 = _T_32 & rowcount_2 == 32'h0 & rowcount_3 != 32'h0 ? 32'h3 : _GEN_247; // @[ivncontrol4.scala 154:100 155:13]
  wire  _T_48 = _T_39 & rowcount_3 == 32'h0; // @[ivncontrol4.scala 157:77]
  wire [31:0] _GEN_249 = _T_39 & rowcount_3 == 32'h0 & rowcount_4 != 32'h0 ? 32'h4 : _GEN_248; // @[ivncontrol4.scala 157:123 158:13]
  wire  _T_59 = _T_48 & rowcount_4 == 32'h0; // @[ivncontrol4.scala 160:100]
  wire  _T_72 = _T_59 & rowcount_5 == 32'h0; // @[ivncontrol4.scala 163:123]
  wire  valid = _k_T_2; // @[ivncontrol4.scala 136:75 137:14 139:14]
  wire [32:0] _T_91 = {{1'd0}, pin}; // @[ivncontrol4.scala 174:27]
  wire [31:0] _GEN_254 = 4'h1 == _T_91[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_255 = 4'h2 == _T_91[3:0] ? rowcount_2 : _GEN_254; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_256 = 4'h3 == _T_91[3:0] ? rowcount_3 : _GEN_255; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_257 = 4'h4 == _T_91[3:0] ? rowcount_4 : _GEN_256; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_258 = 4'h5 == _T_91[3:0] ? rowcount_5 : _GEN_257; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_259 = 4'h6 == _T_91[3:0] ? rowcount_6 : _GEN_258; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_260 = 4'h7 == _T_91[3:0] ? rowcount_7 : _GEN_259; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_261 = 4'h8 == _T_91[3:0] ? rowcount_8 : _GEN_260; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_262 = 4'h9 == _T_91[3:0] ? rowcount_9 : _GEN_261; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_263 = 4'ha == _T_91[3:0] ? rowcount_10 : _GEN_262; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_264 = 4'hb == _T_91[3:0] ? rowcount_11 : _GEN_263; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_265 = 4'hc == _T_91[3:0] ? rowcount_12 : _GEN_264; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_266 = 4'hd == _T_91[3:0] ? rowcount_13 : _GEN_265; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_267 = 4'he == _T_91[3:0] ? rowcount_14 : _GEN_266; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_268 = 4'hf == _T_91[3:0] ? rowcount_15 : _GEN_267; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_381 = _GEN_268 == 32'h1 ? _T_91[31:0] : 32'h13; // @[ivncontrol4.scala 125:17 224:50 225:21]
  wire [31:0] _GEN_382 = _GEN_268 == 32'h2 ? _T_91[31:0] : _GEN_381; // @[ivncontrol4.scala 220:51 221:21]
  wire [31:0] _GEN_383 = _GEN_268 == 32'h2 ? _T_91[31:0] : 32'h2; // @[ivncontrol4.scala 125:17 220:51 222:21]
  wire [31:0] _GEN_384 = _GEN_268 == 32'h3 ? _T_91[31:0] : _GEN_382; // @[ivncontrol4.scala 215:50 216:21]
  wire [31:0] _GEN_385 = _GEN_268 == 32'h3 ? _T_91[31:0] : _GEN_383; // @[ivncontrol4.scala 215:50 217:21]
  wire [31:0] _GEN_386 = _GEN_268 == 32'h3 ? _T_91[31:0] : 32'h9; // @[ivncontrol4.scala 125:17 215:50 218:21]
  wire [31:0] _GEN_387 = _GEN_268 == 32'h4 ? _T_91[31:0] : _GEN_384; // @[ivncontrol4.scala 207:50 208:21]
  wire [31:0] _GEN_388 = _GEN_268 == 32'h4 ? _T_91[31:0] : _GEN_385; // @[ivncontrol4.scala 207:50 209:21]
  wire [31:0] _GEN_389 = _GEN_268 == 32'h4 ? _T_91[31:0] : _GEN_386; // @[ivncontrol4.scala 207:50 210:21]
  wire [31:0] _GEN_390 = _GEN_268 == 32'h4 ? _T_91[31:0] : 32'h8; // @[ivncontrol4.scala 125:17 207:50 211:21]
  wire [31:0] _GEN_391 = _GEN_268 == 32'h5 ? _T_91[31:0] : _GEN_387; // @[ivncontrol4.scala 200:50 201:21]
  wire [31:0] _GEN_392 = _GEN_268 == 32'h5 ? _T_91[31:0] : _GEN_388; // @[ivncontrol4.scala 200:50 202:21]
  wire [31:0] _GEN_393 = _GEN_268 == 32'h5 ? _T_91[31:0] : _GEN_389; // @[ivncontrol4.scala 200:50 203:21]
  wire [31:0] _GEN_394 = _GEN_268 == 32'h5 ? _T_91[31:0] : _GEN_390; // @[ivncontrol4.scala 200:50 204:21]
  wire [31:0] _GEN_395 = _GEN_268 == 32'h5 ? _T_91[31:0] : 32'h10; // @[ivncontrol4.scala 126:18 200:50 205:22]
  wire [31:0] _GEN_396 = _GEN_268 == 32'h6 ? _T_91[31:0] : _GEN_391; // @[ivncontrol4.scala 192:52 193:21]
  wire [31:0] _GEN_397 = _GEN_268 == 32'h6 ? _T_91[31:0] : _GEN_392; // @[ivncontrol4.scala 192:52 194:21]
  wire [31:0] _GEN_398 = _GEN_268 == 32'h6 ? _T_91[31:0] : _GEN_393; // @[ivncontrol4.scala 192:52 195:21]
  wire [31:0] _GEN_399 = _GEN_268 == 32'h6 ? _T_91[31:0] : _GEN_394; // @[ivncontrol4.scala 192:52 196:21]
  wire [31:0] _GEN_400 = _GEN_268 == 32'h6 ? _T_91[31:0] : _GEN_395; // @[ivncontrol4.scala 192:52 197:22]
  wire [31:0] _GEN_401 = _GEN_268 == 32'h6 ? _T_91[31:0] : 32'h6; // @[ivncontrol4.scala 126:18 192:52 198:22]
  wire [31:0] _GEN_402 = _GEN_268 == 32'h7 ? _T_91[31:0] : _GEN_396; // @[ivncontrol4.scala 184:52 185:21]
  wire [31:0] _GEN_403 = _GEN_268 == 32'h7 ? _T_91[31:0] : _GEN_397; // @[ivncontrol4.scala 184:52 186:21]
  wire [31:0] _GEN_404 = _GEN_268 == 32'h7 ? _T_91[31:0] : _GEN_398; // @[ivncontrol4.scala 184:52 187:21]
  wire [31:0] _GEN_405 = _GEN_268 == 32'h7 ? _T_91[31:0] : _GEN_399; // @[ivncontrol4.scala 184:52 188:21]
  wire [31:0] _GEN_406 = _GEN_268 == 32'h7 ? _T_91[31:0] : _GEN_400; // @[ivncontrol4.scala 184:52 189:22]
  wire [31:0] _GEN_407 = _GEN_268 == 32'h7 ? _T_91[31:0] : _GEN_401; // @[ivncontrol4.scala 184:52 190:22]
  wire [31:0] _GEN_408 = _GEN_268 == 32'h7 ? _T_91[31:0] : 32'h17; // @[ivncontrol4.scala 126:18 184:52 191:22]
  wire [31:0] _GEN_409 = _GEN_268 >= 32'h8 ? _T_91[31:0] : _GEN_402; // @[ivncontrol4.scala 174:42 175:21]
  wire [31:0] _GEN_410 = _GEN_268 >= 32'h8 ? _T_91[31:0] : _GEN_403; // @[ivncontrol4.scala 174:42 176:21]
  wire [31:0] _GEN_411 = _GEN_268 >= 32'h8 ? _T_91[31:0] : _GEN_404; // @[ivncontrol4.scala 174:42 177:21]
  wire [31:0] _GEN_412 = _GEN_268 >= 32'h8 ? _T_91[31:0] : _GEN_405; // @[ivncontrol4.scala 174:42 178:21]
  wire [31:0] _GEN_413 = _GEN_268 >= 32'h8 ? _T_91[31:0] : _GEN_406; // @[ivncontrol4.scala 174:42 179:22]
  wire [31:0] _GEN_414 = _GEN_268 >= 32'h8 ? _T_91[31:0] : _GEN_407; // @[ivncontrol4.scala 174:42 180:22]
  wire [31:0] _GEN_415 = _GEN_268 >= 32'h8 ? _T_91[31:0] : _GEN_408; // @[ivncontrol4.scala 174:42 181:22]
  wire [31:0] _GEN_416 = _GEN_268 >= 32'h8 ? _T_91[31:0] : 32'h15; // @[ivncontrol4.scala 126:18 174:42 182:22]
  wire [31:0] _T_127 = 32'h8 - _GEN_268; // @[ivncontrol4.scala 228:18]
  wire [31:0] _i_vn_1_T_15 = 32'h1 + pin; // @[ivncontrol4.scala 229:29]
  wire [31:0] _GEN_529 = _T_127 == 32'h1 ? _i_vn_1_T_15 : _GEN_416; // @[ivncontrol4.scala 269:54 272:22]
  wire [31:0] _GEN_530 = _T_127 == 32'h2 ? _i_vn_1_T_15 : _GEN_415; // @[ivncontrol4.scala 264:54 267:22]
  wire [31:0] _GEN_531 = _T_127 == 32'h2 ? _i_vn_1_T_15 : _GEN_529; // @[ivncontrol4.scala 264:54 268:22]
  wire [31:0] _GEN_532 = _T_127 == 32'h3 ? _i_vn_1_T_15 : _GEN_414; // @[ivncontrol4.scala 257:54 259:22]
  wire [31:0] _GEN_533 = _T_127 == 32'h3 ? _i_vn_1_T_15 : _GEN_530; // @[ivncontrol4.scala 257:54 260:22]
  wire [31:0] _GEN_534 = _T_127 == 32'h3 ? _i_vn_1_T_15 : _GEN_531; // @[ivncontrol4.scala 257:54 261:22]
  wire [31:0] _GEN_535 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_413; // @[ivncontrol4.scala 251:54 253:22]
  wire [31:0] _GEN_536 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_532; // @[ivncontrol4.scala 251:54 254:22]
  wire [31:0] _GEN_537 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_533; // @[ivncontrol4.scala 251:54 255:22]
  wire [31:0] _GEN_538 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_534; // @[ivncontrol4.scala 251:54 256:22]
  wire [31:0] _GEN_539 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_412; // @[ivncontrol4.scala 244:54 246:21]
  wire [31:0] _GEN_540 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_535; // @[ivncontrol4.scala 244:54 247:22]
  wire [31:0] _GEN_541 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_536; // @[ivncontrol4.scala 244:54 248:22]
  wire [31:0] _GEN_542 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_537; // @[ivncontrol4.scala 244:54 249:22]
  wire [31:0] _GEN_543 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_538; // @[ivncontrol4.scala 244:54 250:22]
  wire [31:0] _GEN_544 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_411; // @[ivncontrol4.scala 237:54 238:22]
  wire [31:0] _GEN_545 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_539; // @[ivncontrol4.scala 237:54 239:21]
  wire [31:0] _GEN_546 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_540; // @[ivncontrol4.scala 237:54 240:22]
  wire [31:0] _GEN_547 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_541; // @[ivncontrol4.scala 237:54 241:22]
  wire [31:0] _GEN_548 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_542; // @[ivncontrol4.scala 237:54 242:22]
  wire [31:0] _GEN_549 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_543; // @[ivncontrol4.scala 237:54 243:22]
  wire [31:0] _GEN_550 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_410; // @[ivncontrol4.scala 228:49 229:22]
  wire [31:0] _GEN_551 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_544; // @[ivncontrol4.scala 228:49 230:21]
  wire [31:0] _GEN_552 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_545; // @[ivncontrol4.scala 228:49 231:21]
  wire [31:0] _GEN_553 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_546; // @[ivncontrol4.scala 228:49 232:22]
  wire [31:0] _GEN_554 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_547; // @[ivncontrol4.scala 228:49 233:22]
  wire [31:0] _GEN_555 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_548; // @[ivncontrol4.scala 228:49 234:22]
  wire [31:0] _GEN_556 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_549; // @[ivncontrol4.scala 228:49 235:22]
  wire [31:0] _GEN_574 = 4'h1 == _i_vn_1_T_15[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_575 = 4'h2 == _i_vn_1_T_15[3:0] ? rowcount_2 : _GEN_574; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_576 = 4'h3 == _i_vn_1_T_15[3:0] ? rowcount_3 : _GEN_575; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_577 = 4'h4 == _i_vn_1_T_15[3:0] ? rowcount_4 : _GEN_576; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_578 = 4'h5 == _i_vn_1_T_15[3:0] ? rowcount_5 : _GEN_577; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_579 = 4'h6 == _i_vn_1_T_15[3:0] ? rowcount_6 : _GEN_578; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_580 = 4'h7 == _i_vn_1_T_15[3:0] ? rowcount_7 : _GEN_579; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_581 = 4'h8 == _i_vn_1_T_15[3:0] ? rowcount_8 : _GEN_580; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_582 = 4'h9 == _i_vn_1_T_15[3:0] ? rowcount_9 : _GEN_581; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_583 = 4'ha == _i_vn_1_T_15[3:0] ? rowcount_10 : _GEN_582; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_584 = 4'hb == _i_vn_1_T_15[3:0] ? rowcount_11 : _GEN_583; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_585 = 4'hc == _i_vn_1_T_15[3:0] ? rowcount_12 : _GEN_584; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_586 = 4'hd == _i_vn_1_T_15[3:0] ? rowcount_13 : _GEN_585; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_587 = 4'he == _i_vn_1_T_15[3:0] ? rowcount_14 : _GEN_586; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_588 = 4'hf == _i_vn_1_T_15[3:0] ? rowcount_15 : _GEN_587; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _T_172 = _GEN_268 + _GEN_588; // @[ivncontrol4.scala 275:41]
  wire [31:0] _T_174 = 32'h8 - _T_172; // @[ivncontrol4.scala 275:18]
  wire [31:0] _i_vn_1_T_17 = 32'h2 + pin; // @[ivncontrol4.scala 276:29]
  wire [31:0] _GEN_781 = _T_174 == 32'h1 ? _i_vn_1_T_17 : _GEN_556; // @[ivncontrol4.scala 318:78 321:22]
  wire [31:0] _GEN_782 = _T_174 == 32'h2 ? _i_vn_1_T_17 : _GEN_555; // @[ivncontrol4.scala 312:76 315:22]
  wire [31:0] _GEN_783 = _T_174 == 32'h2 ? _i_vn_1_T_17 : _GEN_781; // @[ivncontrol4.scala 312:76 316:22]
  wire [31:0] _GEN_784 = _T_174 == 32'h3 ? _i_vn_1_T_17 : _GEN_554; // @[ivncontrol4.scala 305:78 307:23]
  wire [31:0] _GEN_785 = _T_174 == 32'h3 ? _i_vn_1_T_17 : _GEN_782; // @[ivncontrol4.scala 305:78 308:22]
  wire [31:0] _GEN_786 = _T_174 == 32'h3 ? _i_vn_1_T_17 : _GEN_783; // @[ivncontrol4.scala 305:78 309:22]
  wire [31:0] _GEN_787 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_553; // @[ivncontrol4.scala 299:78 301:22]
  wire [31:0] _GEN_788 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_784; // @[ivncontrol4.scala 299:78 302:22]
  wire [31:0] _GEN_789 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_785; // @[ivncontrol4.scala 299:78 303:22]
  wire [31:0] _GEN_790 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_786; // @[ivncontrol4.scala 299:78 304:22]
  wire [31:0] _GEN_791 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_552; // @[ivncontrol4.scala 292:76 294:23]
  wire [31:0] _GEN_792 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_787; // @[ivncontrol4.scala 292:76 295:22]
  wire [31:0] _GEN_793 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_788; // @[ivncontrol4.scala 292:76 296:22]
  wire [31:0] _GEN_794 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_789; // @[ivncontrol4.scala 292:76 297:22]
  wire [31:0] _GEN_795 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_790; // @[ivncontrol4.scala 292:76 298:22]
  wire [31:0] _GEN_796 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_551; // @[ivncontrol4.scala 284:77 286:22]
  wire [31:0] _GEN_797 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_791; // @[ivncontrol4.scala 284:77 287:21]
  wire [31:0] _GEN_798 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_792; // @[ivncontrol4.scala 284:77 288:22]
  wire [31:0] _GEN_799 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_793; // @[ivncontrol4.scala 284:77 289:22]
  wire [31:0] _GEN_800 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_794; // @[ivncontrol4.scala 284:77 290:22]
  wire [31:0] _GEN_801 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_795; // @[ivncontrol4.scala 284:77 291:22]
  wire [31:0] _GEN_802 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_550; // @[ivncontrol4.scala 275:73 276:22]
  wire [31:0] _GEN_803 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_796; // @[ivncontrol4.scala 275:73 277:21]
  wire [31:0] _GEN_804 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_797; // @[ivncontrol4.scala 275:73 278:21]
  wire [31:0] _GEN_805 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_798; // @[ivncontrol4.scala 275:73 279:22]
  wire [31:0] _GEN_806 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_799; // @[ivncontrol4.scala 275:73 280:22]
  wire [31:0] _GEN_807 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_800; // @[ivncontrol4.scala 275:73 281:22]
  wire [31:0] _GEN_808 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_801; // @[ivncontrol4.scala 275:73 282:22]
  wire [31:0] _GEN_842 = 4'h1 == _i_vn_1_T_17[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_843 = 4'h2 == _i_vn_1_T_17[3:0] ? rowcount_2 : _GEN_842; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_844 = 4'h3 == _i_vn_1_T_17[3:0] ? rowcount_3 : _GEN_843; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_845 = 4'h4 == _i_vn_1_T_17[3:0] ? rowcount_4 : _GEN_844; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_846 = 4'h5 == _i_vn_1_T_17[3:0] ? rowcount_5 : _GEN_845; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_847 = 4'h6 == _i_vn_1_T_17[3:0] ? rowcount_6 : _GEN_846; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_848 = 4'h7 == _i_vn_1_T_17[3:0] ? rowcount_7 : _GEN_847; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_849 = 4'h8 == _i_vn_1_T_17[3:0] ? rowcount_8 : _GEN_848; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_850 = 4'h9 == _i_vn_1_T_17[3:0] ? rowcount_9 : _GEN_849; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_851 = 4'ha == _i_vn_1_T_17[3:0] ? rowcount_10 : _GEN_850; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_852 = 4'hb == _i_vn_1_T_17[3:0] ? rowcount_11 : _GEN_851; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_853 = 4'hc == _i_vn_1_T_17[3:0] ? rowcount_12 : _GEN_852; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_854 = 4'hd == _i_vn_1_T_17[3:0] ? rowcount_13 : _GEN_853; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_855 = 4'he == _i_vn_1_T_17[3:0] ? rowcount_14 : _GEN_854; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_856 = 4'hf == _i_vn_1_T_17[3:0] ? rowcount_15 : _GEN_855; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _T_254 = _T_172 + _GEN_856; // @[ivncontrol4.scala 326:62]
  wire [31:0] _T_256 = 32'h8 - _T_254; // @[ivncontrol4.scala 326:17]
  wire [31:0] _i_vn_1_T_19 = 32'h3 + pin; // @[ivncontrol4.scala 327:29]
  wire [31:0] _GEN_1145 = _T_256 == 32'h1 ? _i_vn_1_T_19 : _GEN_808; // @[ivncontrol4.scala 369:100 372:22]
  wire [31:0] _GEN_1146 = _T_256 == 32'h2 ? _i_vn_1_T_19 : _GEN_807; // @[ivncontrol4.scala 363:98 366:22]
  wire [31:0] _GEN_1147 = _T_256 == 32'h2 ? _i_vn_1_T_19 : _GEN_1145; // @[ivncontrol4.scala 363:98 367:22]
  wire [31:0] _GEN_1148 = _T_256 == 32'h3 ? _i_vn_1_T_19 : _GEN_806; // @[ivncontrol4.scala 356:100 358:23]
  wire [31:0] _GEN_1149 = _T_256 == 32'h3 ? _i_vn_1_T_19 : _GEN_1146; // @[ivncontrol4.scala 356:100 359:22]
  wire [31:0] _GEN_1150 = _T_256 == 32'h3 ? _i_vn_1_T_19 : _GEN_1147; // @[ivncontrol4.scala 356:100 360:22]
  wire [31:0] _GEN_1151 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_805; // @[ivncontrol4.scala 350:100 352:22]
  wire [31:0] _GEN_1152 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_1148; // @[ivncontrol4.scala 350:100 353:22]
  wire [31:0] _GEN_1153 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_1149; // @[ivncontrol4.scala 350:100 354:22]
  wire [31:0] _GEN_1154 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_1150; // @[ivncontrol4.scala 350:100 355:22]
  wire [31:0] _GEN_1155 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_804; // @[ivncontrol4.scala 343:98 345:23]
  wire [31:0] _GEN_1156 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1151; // @[ivncontrol4.scala 343:98 346:22]
  wire [31:0] _GEN_1157 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1152; // @[ivncontrol4.scala 343:98 347:22]
  wire [31:0] _GEN_1158 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1153; // @[ivncontrol4.scala 343:98 348:22]
  wire [31:0] _GEN_1159 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1154; // @[ivncontrol4.scala 343:98 349:22]
  wire [31:0] _GEN_1160 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_803; // @[ivncontrol4.scala 335:99 337:22]
  wire [31:0] _GEN_1161 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1155; // @[ivncontrol4.scala 335:99 338:21]
  wire [31:0] _GEN_1162 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1156; // @[ivncontrol4.scala 335:99 339:22]
  wire [31:0] _GEN_1163 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1157; // @[ivncontrol4.scala 335:99 340:22]
  wire [31:0] _GEN_1164 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1158; // @[ivncontrol4.scala 335:99 341:22]
  wire [31:0] _GEN_1165 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1159; // @[ivncontrol4.scala 335:99 342:22]
  wire [31:0] _GEN_1166 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_802; // @[ivncontrol4.scala 326:94 327:22]
  wire [31:0] _GEN_1167 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1160; // @[ivncontrol4.scala 326:94 328:21]
  wire [31:0] _GEN_1168 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1161; // @[ivncontrol4.scala 326:94 329:21]
  wire [31:0] _GEN_1169 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1162; // @[ivncontrol4.scala 326:94 330:22]
  wire [31:0] _GEN_1170 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1163; // @[ivncontrol4.scala 326:94 331:22]
  wire [31:0] _GEN_1171 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1164; // @[ivncontrol4.scala 326:94 332:22]
  wire [31:0] _GEN_1172 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1165; // @[ivncontrol4.scala 326:94 333:22]
  wire [31:0] _GEN_1222 = 4'h1 == _i_vn_1_T_19[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1223 = 4'h2 == _i_vn_1_T_19[3:0] ? rowcount_2 : _GEN_1222; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1224 = 4'h3 == _i_vn_1_T_19[3:0] ? rowcount_3 : _GEN_1223; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1225 = 4'h4 == _i_vn_1_T_19[3:0] ? rowcount_4 : _GEN_1224; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1226 = 4'h5 == _i_vn_1_T_19[3:0] ? rowcount_5 : _GEN_1225; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1227 = 4'h6 == _i_vn_1_T_19[3:0] ? rowcount_6 : _GEN_1226; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1228 = 4'h7 == _i_vn_1_T_19[3:0] ? rowcount_7 : _GEN_1227; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1229 = 4'h8 == _i_vn_1_T_19[3:0] ? rowcount_8 : _GEN_1228; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1230 = 4'h9 == _i_vn_1_T_19[3:0] ? rowcount_9 : _GEN_1229; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1231 = 4'ha == _i_vn_1_T_19[3:0] ? rowcount_10 : _GEN_1230; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1232 = 4'hb == _i_vn_1_T_19[3:0] ? rowcount_11 : _GEN_1231; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1233 = 4'hc == _i_vn_1_T_19[3:0] ? rowcount_12 : _GEN_1232; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1234 = 4'hd == _i_vn_1_T_19[3:0] ? rowcount_13 : _GEN_1233; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1235 = 4'he == _i_vn_1_T_19[3:0] ? rowcount_14 : _GEN_1234; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1236 = 4'hf == _i_vn_1_T_19[3:0] ? rowcount_15 : _GEN_1235; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _T_371 = _T_254 + _GEN_1236; // @[ivncontrol4.scala 376:86]
  wire [31:0] _T_373 = 32'h8 - _T_371; // @[ivncontrol4.scala 376:19]
  wire [31:0] _i_vn_1_T_21 = 32'h4 + pin; // @[ivncontrol4.scala 377:29]
  wire [31:0] _GEN_1621 = _T_373 == 32'h1 ? _i_vn_1_T_21 : _GEN_1172; // @[ivncontrol4.scala 419:122 422:22]
  wire [31:0] _GEN_1622 = _T_373 == 32'h2 ? _i_vn_1_T_21 : _GEN_1171; // @[ivncontrol4.scala 413:121 416:22]
  wire [31:0] _GEN_1623 = _T_373 == 32'h2 ? _i_vn_1_T_21 : _GEN_1621; // @[ivncontrol4.scala 413:121 417:22]
  wire [31:0] _GEN_1624 = _T_373 == 32'h3 ? _i_vn_1_T_21 : _GEN_1170; // @[ivncontrol4.scala 406:123 408:23]
  wire [31:0] _GEN_1625 = _T_373 == 32'h3 ? _i_vn_1_T_21 : _GEN_1622; // @[ivncontrol4.scala 406:123 409:22]
  wire [31:0] _GEN_1626 = _T_373 == 32'h3 ? _i_vn_1_T_21 : _GEN_1623; // @[ivncontrol4.scala 406:123 410:22]
  wire [31:0] _GEN_1627 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1169; // @[ivncontrol4.scala 400:122 402:22]
  wire [31:0] _GEN_1628 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1624; // @[ivncontrol4.scala 400:122 403:22]
  wire [31:0] _GEN_1629 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1625; // @[ivncontrol4.scala 400:122 404:22]
  wire [31:0] _GEN_1630 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1626; // @[ivncontrol4.scala 400:122 405:22]
  wire [31:0] _GEN_1631 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1168; // @[ivncontrol4.scala 393:121 395:23]
  wire [31:0] _GEN_1632 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1627; // @[ivncontrol4.scala 393:121 396:22]
  wire [31:0] _GEN_1633 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1628; // @[ivncontrol4.scala 393:121 397:22]
  wire [31:0] _GEN_1634 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1629; // @[ivncontrol4.scala 393:121 398:22]
  wire [31:0] _GEN_1635 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1630; // @[ivncontrol4.scala 393:121 399:22]
  wire [31:0] _GEN_1636 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1167; // @[ivncontrol4.scala 385:121 387:22]
  wire [31:0] _GEN_1637 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1631; // @[ivncontrol4.scala 385:121 388:21]
  wire [31:0] _GEN_1638 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1632; // @[ivncontrol4.scala 385:121 389:22]
  wire [31:0] _GEN_1639 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1633; // @[ivncontrol4.scala 385:121 390:22]
  wire [31:0] _GEN_1640 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1634; // @[ivncontrol4.scala 385:121 391:22]
  wire [31:0] _GEN_1641 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1635; // @[ivncontrol4.scala 385:121 392:22]
  wire [31:0] _GEN_1642 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1166; // @[ivncontrol4.scala 376:118 377:22]
  wire [31:0] _GEN_1643 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1636; // @[ivncontrol4.scala 376:118 378:21]
  wire [31:0] _GEN_1644 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1637; // @[ivncontrol4.scala 376:118 379:21]
  wire [31:0] _GEN_1645 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1638; // @[ivncontrol4.scala 376:118 380:22]
  wire [31:0] _GEN_1646 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1639; // @[ivncontrol4.scala 376:118 381:22]
  wire [31:0] _GEN_1647 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1640; // @[ivncontrol4.scala 376:118 382:22]
  wire [31:0] _GEN_1648 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1641; // @[ivncontrol4.scala 376:118 383:22]
  wire [31:0] _GEN_1714 = 4'h1 == _i_vn_1_T_21[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1715 = 4'h2 == _i_vn_1_T_21[3:0] ? rowcount_2 : _GEN_1714; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1716 = 4'h3 == _i_vn_1_T_21[3:0] ? rowcount_3 : _GEN_1715; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1717 = 4'h4 == _i_vn_1_T_21[3:0] ? rowcount_4 : _GEN_1716; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1718 = 4'h5 == _i_vn_1_T_21[3:0] ? rowcount_5 : _GEN_1717; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1719 = 4'h6 == _i_vn_1_T_21[3:0] ? rowcount_6 : _GEN_1718; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1720 = 4'h7 == _i_vn_1_T_21[3:0] ? rowcount_7 : _GEN_1719; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1721 = 4'h8 == _i_vn_1_T_21[3:0] ? rowcount_8 : _GEN_1720; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1722 = 4'h9 == _i_vn_1_T_21[3:0] ? rowcount_9 : _GEN_1721; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1723 = 4'ha == _i_vn_1_T_21[3:0] ? rowcount_10 : _GEN_1722; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1724 = 4'hb == _i_vn_1_T_21[3:0] ? rowcount_11 : _GEN_1723; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1725 = 4'hc == _i_vn_1_T_21[3:0] ? rowcount_12 : _GEN_1724; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1726 = 4'hd == _i_vn_1_T_21[3:0] ? rowcount_13 : _GEN_1725; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1727 = 4'he == _i_vn_1_T_21[3:0] ? rowcount_14 : _GEN_1726; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1728 = 4'hf == _i_vn_1_T_21[3:0] ? rowcount_15 : _GEN_1727; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _T_523 = _T_371 + _GEN_1728; // @[ivncontrol4.scala 426:108]
  wire [31:0] _T_525 = 32'h8 - _T_523; // @[ivncontrol4.scala 426:19]
  wire [31:0] _i_vn_1_T_23 = 32'h5 + pin; // @[ivncontrol4.scala 427:29]
  wire [31:0] _GEN_2209 = _T_525 == 32'h1 ? _i_vn_1_T_23 : _GEN_1648; // @[ivncontrol4.scala 469:144 472:22]
  wire [31:0] _GEN_2210 = _T_525 == 32'h2 ? _i_vn_1_T_23 : _GEN_1647; // @[ivncontrol4.scala 463:143 466:22]
  wire [31:0] _GEN_2211 = _T_525 == 32'h2 ? _i_vn_1_T_23 : _GEN_2209; // @[ivncontrol4.scala 463:143 467:22]
  wire [31:0] _GEN_2212 = _T_525 == 32'h3 ? _i_vn_1_T_23 : _GEN_1646; // @[ivncontrol4.scala 456:145 458:23]
  wire [31:0] _GEN_2213 = _T_525 == 32'h3 ? _i_vn_1_T_23 : _GEN_2210; // @[ivncontrol4.scala 456:145 459:22]
  wire [31:0] _GEN_2214 = _T_525 == 32'h3 ? _i_vn_1_T_23 : _GEN_2211; // @[ivncontrol4.scala 456:145 460:22]
  wire [31:0] _GEN_2215 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_1645; // @[ivncontrol4.scala 450:143 452:22]
  wire [31:0] _GEN_2216 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_2212; // @[ivncontrol4.scala 450:143 453:22]
  wire [31:0] _GEN_2217 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_2213; // @[ivncontrol4.scala 450:143 454:22]
  wire [31:0] _GEN_2218 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_2214; // @[ivncontrol4.scala 450:143 455:22]
  wire [31:0] _GEN_2219 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_1644; // @[ivncontrol4.scala 443:143 445:23]
  wire [31:0] _GEN_2220 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2215; // @[ivncontrol4.scala 443:143 446:22]
  wire [31:0] _GEN_2221 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2216; // @[ivncontrol4.scala 443:143 447:22]
  wire [31:0] _GEN_2222 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2217; // @[ivncontrol4.scala 443:143 448:22]
  wire [31:0] _GEN_2223 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2218; // @[ivncontrol4.scala 443:143 449:22]
  wire [31:0] _GEN_2224 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_1643; // @[ivncontrol4.scala 435:143 437:22]
  wire [31:0] _GEN_2225 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2219; // @[ivncontrol4.scala 435:143 438:21]
  wire [31:0] _GEN_2226 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2220; // @[ivncontrol4.scala 435:143 439:22]
  wire [31:0] _GEN_2227 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2221; // @[ivncontrol4.scala 435:143 440:22]
  wire [31:0] _GEN_2228 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2222; // @[ivncontrol4.scala 435:143 441:22]
  wire [31:0] _GEN_2229 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2223; // @[ivncontrol4.scala 435:143 442:22]
  wire [31:0] _GEN_2230 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_1642; // @[ivncontrol4.scala 426:140 427:22]
  wire [31:0] _GEN_2231 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2224; // @[ivncontrol4.scala 426:140 428:21]
  wire [31:0] _GEN_2232 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2225; // @[ivncontrol4.scala 426:140 429:21]
  wire [31:0] _GEN_2233 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2226; // @[ivncontrol4.scala 426:140 430:22]
  wire [31:0] _GEN_2234 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2227; // @[ivncontrol4.scala 426:140 431:22]
  wire [31:0] _GEN_2235 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2228; // @[ivncontrol4.scala 426:140 432:22]
  wire [31:0] _GEN_2236 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2229; // @[ivncontrol4.scala 426:140 433:22]
  wire [31:0] _GEN_2318 = 4'h1 == _i_vn_1_T_23[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2319 = 4'h2 == _i_vn_1_T_23[3:0] ? rowcount_2 : _GEN_2318; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2320 = 4'h3 == _i_vn_1_T_23[3:0] ? rowcount_3 : _GEN_2319; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2321 = 4'h4 == _i_vn_1_T_23[3:0] ? rowcount_4 : _GEN_2320; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2322 = 4'h5 == _i_vn_1_T_23[3:0] ? rowcount_5 : _GEN_2321; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2323 = 4'h6 == _i_vn_1_T_23[3:0] ? rowcount_6 : _GEN_2322; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2324 = 4'h7 == _i_vn_1_T_23[3:0] ? rowcount_7 : _GEN_2323; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2325 = 4'h8 == _i_vn_1_T_23[3:0] ? rowcount_8 : _GEN_2324; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2326 = 4'h9 == _i_vn_1_T_23[3:0] ? rowcount_9 : _GEN_2325; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2327 = 4'ha == _i_vn_1_T_23[3:0] ? rowcount_10 : _GEN_2326; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2328 = 4'hb == _i_vn_1_T_23[3:0] ? rowcount_11 : _GEN_2327; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2329 = 4'hc == _i_vn_1_T_23[3:0] ? rowcount_12 : _GEN_2328; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2330 = 4'hd == _i_vn_1_T_23[3:0] ? rowcount_13 : _GEN_2329; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2331 = 4'he == _i_vn_1_T_23[3:0] ? rowcount_14 : _GEN_2330; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2332 = 4'hf == _i_vn_1_T_23[3:0] ? rowcount_15 : _GEN_2331; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _T_710 = _T_523 + _GEN_2332; // @[ivncontrol4.scala 477:130]
  wire [31:0] _T_712 = 32'h8 - _T_710; // @[ivncontrol4.scala 477:19]
  wire [31:0] _i_vn_1_T_25 = 32'h6 + pin; // @[ivncontrol4.scala 478:29]
  wire [31:0] _GEN_2909 = _T_712 == 32'h1 ? _i_vn_1_T_25 : _GEN_2236; // @[ivncontrol4.scala 520:166 523:22]
  wire [31:0] _GEN_2910 = _T_712 == 32'h2 ? _i_vn_1_T_25 : _GEN_2235; // @[ivncontrol4.scala 514:166 517:22]
  wire [31:0] _GEN_2911 = _T_712 == 32'h2 ? _i_vn_1_T_25 : _GEN_2909; // @[ivncontrol4.scala 514:166 518:22]
  wire [31:0] _GEN_2912 = _T_712 == 32'h3 ? _i_vn_1_T_25 : _GEN_2234; // @[ivncontrol4.scala 507:168 509:23]
  wire [31:0] _GEN_2913 = _T_712 == 32'h3 ? _i_vn_1_T_25 : _GEN_2910; // @[ivncontrol4.scala 507:168 510:22]
  wire [31:0] _GEN_2914 = _T_712 == 32'h3 ? _i_vn_1_T_25 : _GEN_2911; // @[ivncontrol4.scala 507:168 511:22]
  wire [31:0] _GEN_2915 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2233; // @[ivncontrol4.scala 501:166 503:22]
  wire [31:0] _GEN_2916 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2912; // @[ivncontrol4.scala 501:166 504:22]
  wire [31:0] _GEN_2917 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2913; // @[ivncontrol4.scala 501:166 505:22]
  wire [31:0] _GEN_2918 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2914; // @[ivncontrol4.scala 501:166 506:22]
  wire [31:0] _GEN_2919 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2232; // @[ivncontrol4.scala 494:166 496:23]
  wire [31:0] _GEN_2920 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2915; // @[ivncontrol4.scala 494:166 497:22]
  wire [31:0] _GEN_2921 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2916; // @[ivncontrol4.scala 494:166 498:22]
  wire [31:0] _GEN_2922 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2917; // @[ivncontrol4.scala 494:166 499:22]
  wire [31:0] _GEN_2923 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2918; // @[ivncontrol4.scala 494:166 500:22]
  wire [31:0] _GEN_2924 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2231; // @[ivncontrol4.scala 486:166 488:22]
  wire [31:0] _GEN_2925 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2919; // @[ivncontrol4.scala 486:166 489:21]
  wire [31:0] _GEN_2926 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2920; // @[ivncontrol4.scala 486:166 490:22]
  wire [31:0] _GEN_2927 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2921; // @[ivncontrol4.scala 486:166 491:22]
  wire [31:0] _GEN_2928 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2922; // @[ivncontrol4.scala 486:166 492:22]
  wire [31:0] _GEN_2929 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2923; // @[ivncontrol4.scala 486:166 493:22]
  wire [31:0] _GEN_2930 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2230; // @[ivncontrol4.scala 477:162 478:22]
  wire [31:0] _GEN_2931 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2924; // @[ivncontrol4.scala 477:162 479:21]
  wire [31:0] _GEN_2932 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2925; // @[ivncontrol4.scala 477:162 480:21]
  wire [31:0] _GEN_2933 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2926; // @[ivncontrol4.scala 477:162 481:22]
  wire [31:0] _GEN_2934 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2927; // @[ivncontrol4.scala 477:162 482:22]
  wire [31:0] _GEN_2935 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2928; // @[ivncontrol4.scala 477:162 483:22]
  wire [31:0] _GEN_2936 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2929; // @[ivncontrol4.scala 477:162 484:22]
  wire [31:0] _GEN_3034 = 4'h1 == _i_vn_1_T_25[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3035 = 4'h2 == _i_vn_1_T_25[3:0] ? rowcount_2 : _GEN_3034; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3036 = 4'h3 == _i_vn_1_T_25[3:0] ? rowcount_3 : _GEN_3035; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3037 = 4'h4 == _i_vn_1_T_25[3:0] ? rowcount_4 : _GEN_3036; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3038 = 4'h5 == _i_vn_1_T_25[3:0] ? rowcount_5 : _GEN_3037; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3039 = 4'h6 == _i_vn_1_T_25[3:0] ? rowcount_6 : _GEN_3038; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3040 = 4'h7 == _i_vn_1_T_25[3:0] ? rowcount_7 : _GEN_3039; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3041 = 4'h8 == _i_vn_1_T_25[3:0] ? rowcount_8 : _GEN_3040; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3042 = 4'h9 == _i_vn_1_T_25[3:0] ? rowcount_9 : _GEN_3041; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3043 = 4'ha == _i_vn_1_T_25[3:0] ? rowcount_10 : _GEN_3042; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3044 = 4'hb == _i_vn_1_T_25[3:0] ? rowcount_11 : _GEN_3043; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3045 = 4'hc == _i_vn_1_T_25[3:0] ? rowcount_12 : _GEN_3044; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3046 = 4'hd == _i_vn_1_T_25[3:0] ? rowcount_13 : _GEN_3045; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3047 = 4'he == _i_vn_1_T_25[3:0] ? rowcount_14 : _GEN_3046; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3048 = 4'hf == _i_vn_1_T_25[3:0] ? rowcount_15 : _GEN_3047; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _T_932 = _T_710 + _GEN_3048; // @[ivncontrol4.scala 528:152]
  wire [31:0] _T_934 = 32'h8 - _T_932; // @[ivncontrol4.scala 528:19]
  wire [31:0] _i_vn_1_T_27 = 32'h7 + pin; // @[ivncontrol4.scala 529:29]
  wire [31:0] _GEN_3721 = _T_934 == 32'h1 ? _i_vn_1_T_27 : _GEN_2936; // @[ivncontrol4.scala 571:188 574:22]
  wire [31:0] _GEN_3722 = _T_934 == 32'h2 ? _i_vn_1_T_27 : _GEN_2935; // @[ivncontrol4.scala 565:188 568:22]
  wire [31:0] _GEN_3723 = _T_934 == 32'h2 ? _i_vn_1_T_27 : _GEN_3721; // @[ivncontrol4.scala 565:188 569:22]
  wire [31:0] _GEN_3724 = _T_934 == 32'h3 ? _i_vn_1_T_27 : _GEN_2934; // @[ivncontrol4.scala 558:190 560:23]
  wire [31:0] _GEN_3725 = _T_934 == 32'h3 ? _i_vn_1_T_27 : _GEN_3722; // @[ivncontrol4.scala 558:190 561:22]
  wire [31:0] _GEN_3726 = _T_934 == 32'h3 ? _i_vn_1_T_27 : _GEN_3723; // @[ivncontrol4.scala 558:190 562:22]
  wire [31:0] _GEN_3727 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_2933; // @[ivncontrol4.scala 552:188 554:22]
  wire [31:0] _GEN_3728 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_3724; // @[ivncontrol4.scala 552:188 555:22]
  wire [31:0] _GEN_3729 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_3725; // @[ivncontrol4.scala 552:188 556:22]
  wire [31:0] _GEN_3730 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_3726; // @[ivncontrol4.scala 552:188 557:22]
  wire [31:0] _GEN_3731 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_2932; // @[ivncontrol4.scala 545:188 547:23]
  wire [31:0] _GEN_3732 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3727; // @[ivncontrol4.scala 545:188 548:22]
  wire [31:0] _GEN_3733 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3728; // @[ivncontrol4.scala 545:188 549:22]
  wire [31:0] _GEN_3734 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3729; // @[ivncontrol4.scala 545:188 550:22]
  wire [31:0] _GEN_3735 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3730; // @[ivncontrol4.scala 545:188 551:22]
  wire [31:0] _GEN_3736 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_2931; // @[ivncontrol4.scala 537:188 539:22]
  wire [31:0] _GEN_3737 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3731; // @[ivncontrol4.scala 537:188 540:21]
  wire [31:0] _GEN_3738 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3732; // @[ivncontrol4.scala 537:188 541:22]
  wire [31:0] _GEN_3739 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3733; // @[ivncontrol4.scala 537:188 542:22]
  wire [31:0] _GEN_3740 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3734; // @[ivncontrol4.scala 537:188 543:22]
  wire [31:0] _GEN_3741 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3735; // @[ivncontrol4.scala 537:188 544:22]
  wire [31:0] _GEN_3742 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_2930; // @[ivncontrol4.scala 528:184 529:22]
  wire [31:0] _GEN_3743 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3736; // @[ivncontrol4.scala 528:184 530:21]
  wire [31:0] _GEN_3744 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3737; // @[ivncontrol4.scala 528:184 531:21]
  wire [31:0] _GEN_3745 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3738; // @[ivncontrol4.scala 528:184 532:22]
  wire [31:0] _GEN_3746 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3739; // @[ivncontrol4.scala 528:184 533:22]
  wire [31:0] _GEN_3747 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3740; // @[ivncontrol4.scala 528:184 534:22]
  wire [31:0] _GEN_3748 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3741; // @[ivncontrol4.scala 528:184 535:22]
  wire [31:0] _GEN_3749 = _GEN_244 ? _GEN_409 : 32'h13; // @[ivncontrol4.scala 125:17 172:28]
  wire [31:0] _GEN_3750 = _GEN_244 ? _GEN_3742 : 32'h2; // @[ivncontrol4.scala 125:17 172:28]
  wire [31:0] _GEN_3751 = _GEN_244 ? _GEN_3743 : 32'h9; // @[ivncontrol4.scala 125:17 172:28]
  wire [31:0] _GEN_3752 = _GEN_244 ? _GEN_3744 : 32'h8; // @[ivncontrol4.scala 125:17 172:28]
  wire [31:0] _GEN_3753 = _GEN_244 ? _GEN_3745 : 32'h10; // @[ivncontrol4.scala 126:18 172:28]
  wire [31:0] _GEN_3754 = _GEN_244 ? _GEN_3746 : 32'h6; // @[ivncontrol4.scala 126:18 172:28]
  wire [31:0] _GEN_3755 = _GEN_244 ? _GEN_3747 : 32'h17; // @[ivncontrol4.scala 126:18 172:28]
  wire [31:0] _GEN_3756 = _GEN_244 ? _GEN_3748 : 32'h15; // @[ivncontrol4.scala 126:18 172:28]
  wire [31:0] _GEN_4137 = reset ? 32'h0 : _GEN_3749; // @[ivncontrol4.scala 16:{23,23}]
  wire [31:0] _GEN_4138 = reset ? 32'h0 : _GEN_3750; // @[ivncontrol4.scala 16:{23,23}]
  wire [31:0] _GEN_4139 = reset ? 32'h0 : _GEN_3751; // @[ivncontrol4.scala 16:{23,23}]
  wire [31:0] _GEN_4140 = reset ? 32'h0 : _GEN_3752; // @[ivncontrol4.scala 16:{23,23}]
  wire [31:0] _GEN_4141 = reset ? 32'h0 : _GEN_3753; // @[ivncontrol4.scala 17:{24,24}]
  wire [31:0] _GEN_4142 = reset ? 32'h0 : _GEN_3754; // @[ivncontrol4.scala 17:{24,24}]
  wire [31:0] _GEN_4143 = reset ? 32'h0 : _GEN_3755; // @[ivncontrol4.scala 17:{24,24}]
  wire [31:0] _GEN_4144 = reset ? 32'h0 : _GEN_3756; // @[ivncontrol4.scala 17:{24,24}]
  assign io_o_vn_0 = i_vn_0; // @[ivncontrol4.scala 121:13]
  assign io_o_vn_1 = i_vn_1; // @[ivncontrol4.scala 121:13]
  assign io_o_vn_2 = i_vn_2; // @[ivncontrol4.scala 121:13]
  assign io_o_vn_3 = i_vn_3; // @[ivncontrol4.scala 121:13]
  assign io_o_vn2_0 = i_vn2_0; // @[ivncontrol4.scala 122:14]
  assign io_o_vn2_1 = i_vn2_1; // @[ivncontrol4.scala 122:14]
  assign io_o_vn2_2 = i_vn2_2; // @[ivncontrol4.scala 122:14]
  assign io_o_vn2_3 = i_vn2_3; // @[ivncontrol4.scala 122:14]
  always @(posedge clock) begin
    i_vn_0 <= _GEN_4137[4:0]; // @[ivncontrol4.scala 16:{23,23}]
    i_vn_1 <= _GEN_4138[4:0]; // @[ivncontrol4.scala 16:{23,23}]
    i_vn_2 <= _GEN_4139[4:0]; // @[ivncontrol4.scala 16:{23,23}]
    i_vn_3 <= _GEN_4140[4:0]; // @[ivncontrol4.scala 16:{23,23}]
    i_vn2_0 <= _GEN_4141[4:0]; // @[ivncontrol4.scala 17:{24,24}]
    i_vn2_1 <= _GEN_4142[4:0]; // @[ivncontrol4.scala 17:{24,24}]
    i_vn2_2 <= _GEN_4143[4:0]; // @[ivncontrol4.scala 17:{24,24}]
    i_vn2_3 <= _GEN_4144[4:0]; // @[ivncontrol4.scala 17:{24,24}]
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_0 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_0 <= count_0; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_1 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_1 <= count_1; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_2 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_2 <= count_2; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_3 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_3 <= count_3; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_4 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_4 <= count_4; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_5 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_5 <= count_5; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_6 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_6 <= count_6; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_7 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_7 <= count_7; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_8 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_8 <= 32'h0; // @[ivncontrol4.scala 81:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_9 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_9 <= 32'h0; // @[ivncontrol4.scala 81:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_10 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_10 <= 32'h0; // @[ivncontrol4.scala 81:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_11 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_11 <= 32'h0; // @[ivncontrol4.scala 81:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_12 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_12 <= 32'h0; // @[ivncontrol4.scala 81:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_13 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_13 <= 32'h0; // @[ivncontrol4.scala 81:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_14 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_14 <= 32'h0; // @[ivncontrol4.scala 81:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_15 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end
    if (reset) begin // @[ivncontrol4.scala 31:22]
      pin <= 32'h0; // @[ivncontrol4.scala 31:22]
    end else if (_T_72 & rowcount_6 == 32'h0 & rowcount_7 != 32'h0) begin // @[ivncontrol4.scala 166:192]
      pin <= 32'h7; // @[ivncontrol4.scala 167:13]
    end else if (_T_59 & rowcount_5 == 32'h0 & rowcount_6 != 32'h0) begin // @[ivncontrol4.scala 163:169]
      pin <= 32'h6; // @[ivncontrol4.scala 164:13]
    end else if (_T_48 & rowcount_4 == 32'h0 & rowcount_5 != 32'h0) begin // @[ivncontrol4.scala 160:146]
      pin <= 32'h5; // @[ivncontrol4.scala 161:13]
    end else begin
      pin <= _GEN_249;
    end
    if (reset) begin // @[ivncontrol4.scala 35:20]
      i <= 32'h0; // @[ivncontrol4.scala 35:20]
    end else if (i < 32'h7 & _k_T_1) begin // @[ivncontrol4.scala 103:74]
      i <= _i_T_1; // @[ivncontrol4.scala 104:11]
    end
    if (reset) begin // @[ivncontrol4.scala 36:20]
      j <= 32'h0; // @[ivncontrol4.scala 36:20]
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 107:71]
      j <= _j_T_1; // @[ivncontrol4.scala 108:11]
    end else if (!(_k_T_2)) begin // @[ivncontrol4.scala 110:81]
      j <= 32'h0; // @[ivncontrol4.scala 114:11]
    end
    if (3'h0 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h0 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h0 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h0 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h0 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h0 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h0 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h0 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h0 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_0 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h1 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_1 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h2 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_2 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h3 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_3 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h4 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_4 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h5 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_5 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h6 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_6 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h7 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_7 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  i_vn_0 = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  i_vn_1 = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  i_vn_2 = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  i_vn_3 = _RAND_3[4:0];
  _RAND_4 = {1{`RANDOM}};
  i_vn2_0 = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  i_vn2_1 = _RAND_5[4:0];
  _RAND_6 = {1{`RANDOM}};
  i_vn2_2 = _RAND_6[4:0];
  _RAND_7 = {1{`RANDOM}};
  i_vn2_3 = _RAND_7[4:0];
  _RAND_8 = {1{`RANDOM}};
  rowcount_0 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  rowcount_1 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  rowcount_2 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  rowcount_3 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  rowcount_4 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  rowcount_5 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  rowcount_6 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  rowcount_7 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  rowcount_8 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  rowcount_9 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  rowcount_10 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  rowcount_11 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  rowcount_12 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  rowcount_13 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  rowcount_14 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  rowcount_15 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  pin = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  i = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  j = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  mat_0_0 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  mat_0_1 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  mat_0_2 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  mat_0_3 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  mat_0_4 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  mat_0_5 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  mat_0_6 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  mat_0_7 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  mat_1_0 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  mat_1_1 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  mat_1_2 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  mat_1_3 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  mat_1_4 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  mat_1_5 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  mat_1_6 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  mat_1_7 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  mat_2_0 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  mat_2_1 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  mat_2_2 = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  mat_2_3 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  mat_2_4 = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  mat_2_5 = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  mat_2_6 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  mat_2_7 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  mat_3_0 = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  mat_3_1 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  mat_3_2 = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  mat_3_3 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  mat_3_4 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  mat_3_5 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  mat_3_6 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  mat_3_7 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  mat_4_0 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  mat_4_1 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  mat_4_2 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  mat_4_3 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  mat_4_4 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  mat_4_5 = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  mat_4_6 = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  mat_4_7 = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  mat_5_0 = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  mat_5_1 = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  mat_5_2 = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  mat_5_3 = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  mat_5_4 = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  mat_5_5 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  mat_5_6 = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  mat_5_7 = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  mat_6_0 = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  mat_6_1 = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  mat_6_2 = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  mat_6_3 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  mat_6_4 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  mat_6_5 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  mat_6_6 = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  mat_6_7 = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  mat_7_0 = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  mat_7_1 = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  mat_7_2 = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  mat_7_3 = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  mat_7_4 = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  mat_7_5 = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  mat_7_6 = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  mat_7_7 = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  count_0 = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  count_1 = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  count_2 = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  count_3 = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  count_4 = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  count_5 = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  count_6 = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  count_7 = _RAND_98[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ivncontrol4_2(
  input         clock,
  input         reset,
  input  [15:0] io_Stationary_matrix_0_0,
  input  [15:0] io_Stationary_matrix_0_1,
  input  [15:0] io_Stationary_matrix_0_2,
  input  [15:0] io_Stationary_matrix_0_3,
  input  [15:0] io_Stationary_matrix_0_4,
  input  [15:0] io_Stationary_matrix_0_5,
  input  [15:0] io_Stationary_matrix_0_6,
  input  [15:0] io_Stationary_matrix_0_7,
  input  [15:0] io_Stationary_matrix_1_0,
  input  [15:0] io_Stationary_matrix_1_1,
  input  [15:0] io_Stationary_matrix_1_2,
  input  [15:0] io_Stationary_matrix_1_3,
  input  [15:0] io_Stationary_matrix_1_4,
  input  [15:0] io_Stationary_matrix_1_5,
  input  [15:0] io_Stationary_matrix_1_6,
  input  [15:0] io_Stationary_matrix_1_7,
  input  [15:0] io_Stationary_matrix_2_0,
  input  [15:0] io_Stationary_matrix_2_1,
  input  [15:0] io_Stationary_matrix_2_2,
  input  [15:0] io_Stationary_matrix_2_3,
  input  [15:0] io_Stationary_matrix_2_4,
  input  [15:0] io_Stationary_matrix_2_5,
  input  [15:0] io_Stationary_matrix_2_6,
  input  [15:0] io_Stationary_matrix_2_7,
  input  [15:0] io_Stationary_matrix_3_0,
  input  [15:0] io_Stationary_matrix_3_1,
  input  [15:0] io_Stationary_matrix_3_2,
  input  [15:0] io_Stationary_matrix_3_3,
  input  [15:0] io_Stationary_matrix_3_4,
  input  [15:0] io_Stationary_matrix_3_5,
  input  [15:0] io_Stationary_matrix_3_6,
  input  [15:0] io_Stationary_matrix_3_7,
  input  [15:0] io_Stationary_matrix_4_0,
  input  [15:0] io_Stationary_matrix_4_1,
  input  [15:0] io_Stationary_matrix_4_2,
  input  [15:0] io_Stationary_matrix_4_3,
  input  [15:0] io_Stationary_matrix_4_4,
  input  [15:0] io_Stationary_matrix_4_5,
  input  [15:0] io_Stationary_matrix_4_6,
  input  [15:0] io_Stationary_matrix_4_7,
  input  [15:0] io_Stationary_matrix_5_0,
  input  [15:0] io_Stationary_matrix_5_1,
  input  [15:0] io_Stationary_matrix_5_2,
  input  [15:0] io_Stationary_matrix_5_3,
  input  [15:0] io_Stationary_matrix_5_4,
  input  [15:0] io_Stationary_matrix_5_5,
  input  [15:0] io_Stationary_matrix_5_6,
  input  [15:0] io_Stationary_matrix_5_7,
  input  [15:0] io_Stationary_matrix_6_0,
  input  [15:0] io_Stationary_matrix_6_1,
  input  [15:0] io_Stationary_matrix_6_2,
  input  [15:0] io_Stationary_matrix_6_3,
  input  [15:0] io_Stationary_matrix_6_4,
  input  [15:0] io_Stationary_matrix_6_5,
  input  [15:0] io_Stationary_matrix_6_6,
  input  [15:0] io_Stationary_matrix_6_7,
  input  [15:0] io_Stationary_matrix_7_0,
  input  [15:0] io_Stationary_matrix_7_1,
  input  [15:0] io_Stationary_matrix_7_2,
  input  [15:0] io_Stationary_matrix_7_3,
  input  [15:0] io_Stationary_matrix_7_4,
  input  [15:0] io_Stationary_matrix_7_5,
  input  [15:0] io_Stationary_matrix_7_6,
  input  [15:0] io_Stationary_matrix_7_7,
  output [4:0]  io_o_vn_0,
  output [4:0]  io_o_vn_1,
  output [4:0]  io_o_vn_2,
  output [4:0]  io_o_vn_3,
  output [4:0]  io_o_vn2_0,
  output [4:0]  io_o_vn2_1,
  output [4:0]  io_o_vn2_2,
  output [4:0]  io_o_vn2_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
`endif // RANDOMIZE_REG_INIT
  reg [4:0] i_vn_0; // @[ivncontrol4.scala 16:23]
  reg [4:0] i_vn_1; // @[ivncontrol4.scala 16:23]
  reg [4:0] i_vn_2; // @[ivncontrol4.scala 16:23]
  reg [4:0] i_vn_3; // @[ivncontrol4.scala 16:23]
  reg [4:0] i_vn2_0; // @[ivncontrol4.scala 17:24]
  reg [4:0] i_vn2_1; // @[ivncontrol4.scala 17:24]
  reg [4:0] i_vn2_2; // @[ivncontrol4.scala 17:24]
  reg [4:0] i_vn2_3; // @[ivncontrol4.scala 17:24]
  reg [31:0] rowcount_0; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_1; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_2; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_3; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_4; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_5; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_6; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_7; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_8; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_9; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_10; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_11; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_12; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_13; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_14; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_15; // @[ivncontrol4.scala 21:27]
  reg [31:0] pin; // @[ivncontrol4.scala 31:22]
  reg [31:0] i; // @[ivncontrol4.scala 35:20]
  reg [31:0] j; // @[ivncontrol4.scala 36:20]
  wire  _k_T_1 = j == 32'h7; // @[ivncontrol4.scala 38:37]
  wire  _k_T_2 = i == 32'h7 & j == 32'h7; // @[ivncontrol4.scala 38:31]
  reg [31:0] mat_0_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_0_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_0_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_0_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_0_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_0_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_0_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_0_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] count_0; // @[ivncontrol4.scala 52:20]
  reg [31:0] count_1; // @[ivncontrol4.scala 52:20]
  reg [31:0] count_2; // @[ivncontrol4.scala 52:20]
  reg [31:0] count_3; // @[ivncontrol4.scala 52:20]
  reg [31:0] count_4; // @[ivncontrol4.scala 52:20]
  reg [31:0] count_5; // @[ivncontrol4.scala 52:20]
  reg [31:0] count_6; // @[ivncontrol4.scala 52:20]
  reg [31:0] count_7; // @[ivncontrol4.scala 52:20]
  wire [15:0] _GEN_66 = 3'h0 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_0_1 : io_Stationary_matrix_0_0; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_67 = 3'h0 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_0_2 : _GEN_66; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_68 = 3'h0 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_0_3 : _GEN_67; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_69 = 3'h0 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_0_4 : _GEN_68; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_70 = 3'h0 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_0_5 : _GEN_69; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_71 = 3'h0 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_0_6 : _GEN_70; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_72 = 3'h0 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_0_7 : _GEN_71; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_73 = 3'h1 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_1_0 : _GEN_72; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_74 = 3'h1 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_1_1 : _GEN_73; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_75 = 3'h1 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_1_2 : _GEN_74; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_76 = 3'h1 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_1_3 : _GEN_75; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_77 = 3'h1 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_1_4 : _GEN_76; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_78 = 3'h1 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_1_5 : _GEN_77; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_79 = 3'h1 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_1_6 : _GEN_78; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_80 = 3'h1 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_1_7 : _GEN_79; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_81 = 3'h2 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_2_0 : _GEN_80; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_82 = 3'h2 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_2_1 : _GEN_81; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_83 = 3'h2 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_2_2 : _GEN_82; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_84 = 3'h2 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_2_3 : _GEN_83; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_85 = 3'h2 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_2_4 : _GEN_84; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_86 = 3'h2 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_2_5 : _GEN_85; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_87 = 3'h2 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_2_6 : _GEN_86; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_88 = 3'h2 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_2_7 : _GEN_87; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_89 = 3'h3 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_3_0 : _GEN_88; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_90 = 3'h3 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_3_1 : _GEN_89; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_91 = 3'h3 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_3_2 : _GEN_90; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_92 = 3'h3 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_3_3 : _GEN_91; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_93 = 3'h3 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_3_4 : _GEN_92; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_94 = 3'h3 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_3_5 : _GEN_93; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_95 = 3'h3 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_3_6 : _GEN_94; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_96 = 3'h3 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_3_7 : _GEN_95; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_97 = 3'h4 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_4_0 : _GEN_96; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_98 = 3'h4 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_4_1 : _GEN_97; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_99 = 3'h4 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_4_2 : _GEN_98; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_100 = 3'h4 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_4_3 : _GEN_99; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_101 = 3'h4 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_4_4 : _GEN_100; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_102 = 3'h4 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_4_5 : _GEN_101; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_103 = 3'h4 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_4_6 : _GEN_102; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_104 = 3'h4 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_4_7 : _GEN_103; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_105 = 3'h5 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_5_0 : _GEN_104; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_106 = 3'h5 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_5_1 : _GEN_105; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_107 = 3'h5 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_5_2 : _GEN_106; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_108 = 3'h5 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_5_3 : _GEN_107; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_109 = 3'h5 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_5_4 : _GEN_108; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_110 = 3'h5 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_5_5 : _GEN_109; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_111 = 3'h5 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_5_6 : _GEN_110; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_112 = 3'h5 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_5_7 : _GEN_111; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_113 = 3'h6 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_6_0 : _GEN_112; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_114 = 3'h6 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_6_1 : _GEN_113; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_115 = 3'h6 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_6_2 : _GEN_114; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_116 = 3'h6 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_6_3 : _GEN_115; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_117 = 3'h6 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_6_4 : _GEN_116; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_118 = 3'h6 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_6_5 : _GEN_117; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_119 = 3'h6 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_6_6 : _GEN_118; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_120 = 3'h6 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_6_7 : _GEN_119; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_121 = 3'h7 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_7_0 : _GEN_120; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_122 = 3'h7 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_7_1 : _GEN_121; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_123 = 3'h7 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_7_2 : _GEN_122; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_124 = 3'h7 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_7_3 : _GEN_123; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_125 = 3'h7 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_7_4 : _GEN_124; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_126 = 3'h7 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_7_5 : _GEN_125; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_127 = 3'h7 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_7_6 : _GEN_126; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_128 = 3'h7 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_7_7 : _GEN_127; // @[ivncontrol4.scala 57:{15,15}]
  wire [31:0] _mat_T_3_T_4 = {{16'd0}, _GEN_128}; // @[ivncontrol4.scala 57:{15,15}]
  wire  _GEN_225 = count_7 >= 32'h8; // @[ivncontrol4.scala 66:28 67:16]
  wire  valid1 = count_7 >= 32'h8; // @[ivncontrol4.scala 66:28 67:16]
  wire [31:0] _GEN_194 = 3'h1 == i[2:0] ? count_1 : count_0; // @[ivncontrol4.scala 60:{33,33}]
  wire [31:0] _GEN_195 = 3'h2 == i[2:0] ? count_2 : _GEN_194; // @[ivncontrol4.scala 60:{33,33}]
  wire [31:0] _GEN_196 = 3'h3 == i[2:0] ? count_3 : _GEN_195; // @[ivncontrol4.scala 60:{33,33}]
  wire [31:0] _GEN_197 = 3'h4 == i[2:0] ? count_4 : _GEN_196; // @[ivncontrol4.scala 60:{33,33}]
  wire [31:0] _GEN_198 = 3'h5 == i[2:0] ? count_5 : _GEN_197; // @[ivncontrol4.scala 60:{33,33}]
  wire [31:0] _GEN_199 = 3'h6 == i[2:0] ? count_6 : _GEN_198; // @[ivncontrol4.scala 60:{33,33}]
  wire [31:0] _GEN_200 = 3'h7 == i[2:0] ? count_7 : _GEN_199; // @[ivncontrol4.scala 60:{33,33}]
  wire [31:0] _count_T_2 = _GEN_200 + 32'h1; // @[ivncontrol4.scala 60:33]
  wire [31:0] _i_T_1 = i + 32'h1; // @[ivncontrol4.scala 104:16]
  wire [31:0] _j_T_1 = j + 32'h1; // @[ivncontrol4.scala 108:16]
  wire  _GEN_244 = _k_T_2; // @[ivncontrol4.scala 136:75 137:14 139:14]
  wire [31:0] _GEN_245 = rowcount_0 != 32'h0 ? 32'h0 : pin; // @[ivncontrol4.scala 145:30 146:13 31:22]
  wire  _T_27 = rowcount_0 == 32'h0; // @[ivncontrol4.scala 148:23]
  wire [31:0] _GEN_246 = rowcount_0 == 32'h0 & rowcount_1 != 32'h0 ? 32'h1 : _GEN_245; // @[ivncontrol4.scala 148:54 149:13]
  wire  _T_32 = _T_27 & rowcount_1 == 32'h0; // @[ivncontrol4.scala 151:31]
  wire [31:0] _GEN_247 = _T_27 & rowcount_1 == 32'h0 & rowcount_2 != 32'h0 ? 32'h2 : _GEN_246; // @[ivncontrol4.scala 151:77 152:13]
  wire  _T_39 = _T_32 & rowcount_2 == 32'h0; // @[ivncontrol4.scala 154:54]
  wire [31:0] _GEN_248 = _T_32 & rowcount_2 == 32'h0 & rowcount_3 != 32'h0 ? 32'h3 : _GEN_247; // @[ivncontrol4.scala 154:100 155:13]
  wire  _T_48 = _T_39 & rowcount_3 == 32'h0; // @[ivncontrol4.scala 157:77]
  wire [31:0] _GEN_249 = _T_39 & rowcount_3 == 32'h0 & rowcount_4 != 32'h0 ? 32'h4 : _GEN_248; // @[ivncontrol4.scala 157:123 158:13]
  wire  _T_59 = _T_48 & rowcount_4 == 32'h0; // @[ivncontrol4.scala 160:100]
  wire  _T_72 = _T_59 & rowcount_5 == 32'h0; // @[ivncontrol4.scala 163:123]
  wire  valid = _k_T_2; // @[ivncontrol4.scala 136:75 137:14 139:14]
  wire [32:0] _T_91 = {{1'd0}, pin}; // @[ivncontrol4.scala 174:27]
  wire [31:0] _GEN_254 = 4'h1 == _T_91[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_255 = 4'h2 == _T_91[3:0] ? rowcount_2 : _GEN_254; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_256 = 4'h3 == _T_91[3:0] ? rowcount_3 : _GEN_255; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_257 = 4'h4 == _T_91[3:0] ? rowcount_4 : _GEN_256; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_258 = 4'h5 == _T_91[3:0] ? rowcount_5 : _GEN_257; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_259 = 4'h6 == _T_91[3:0] ? rowcount_6 : _GEN_258; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_260 = 4'h7 == _T_91[3:0] ? rowcount_7 : _GEN_259; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_261 = 4'h8 == _T_91[3:0] ? rowcount_8 : _GEN_260; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_262 = 4'h9 == _T_91[3:0] ? rowcount_9 : _GEN_261; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_263 = 4'ha == _T_91[3:0] ? rowcount_10 : _GEN_262; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_264 = 4'hb == _T_91[3:0] ? rowcount_11 : _GEN_263; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_265 = 4'hc == _T_91[3:0] ? rowcount_12 : _GEN_264; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_266 = 4'hd == _T_91[3:0] ? rowcount_13 : _GEN_265; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_267 = 4'he == _T_91[3:0] ? rowcount_14 : _GEN_266; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_268 = 4'hf == _T_91[3:0] ? rowcount_15 : _GEN_267; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_381 = _GEN_268 == 32'h1 ? _T_91[31:0] : 32'h18; // @[ivncontrol4.scala 125:17 224:50 225:21]
  wire [31:0] _GEN_382 = _GEN_268 == 32'h2 ? _T_91[31:0] : _GEN_381; // @[ivncontrol4.scala 220:51 221:21]
  wire [31:0] _GEN_383 = _GEN_268 == 32'h2 ? _T_91[31:0] : 32'h1e; // @[ivncontrol4.scala 125:17 220:51 222:21]
  wire [31:0] _GEN_384 = _GEN_268 == 32'h3 ? _T_91[31:0] : _GEN_382; // @[ivncontrol4.scala 215:50 216:21]
  wire [31:0] _GEN_385 = _GEN_268 == 32'h3 ? _T_91[31:0] : _GEN_383; // @[ivncontrol4.scala 215:50 217:21]
  wire [31:0] _GEN_386 = _GEN_268 == 32'h3 ? _T_91[31:0] : 32'h1e; // @[ivncontrol4.scala 125:17 215:50 218:21]
  wire [31:0] _GEN_387 = _GEN_268 == 32'h4 ? _T_91[31:0] : _GEN_384; // @[ivncontrol4.scala 207:50 208:21]
  wire [31:0] _GEN_388 = _GEN_268 == 32'h4 ? _T_91[31:0] : _GEN_385; // @[ivncontrol4.scala 207:50 209:21]
  wire [31:0] _GEN_389 = _GEN_268 == 32'h4 ? _T_91[31:0] : _GEN_386; // @[ivncontrol4.scala 207:50 210:21]
  wire [31:0] _GEN_390 = _GEN_268 == 32'h4 ? _T_91[31:0] : 32'h14; // @[ivncontrol4.scala 125:17 207:50 211:21]
  wire [31:0] _GEN_391 = _GEN_268 == 32'h5 ? _T_91[31:0] : _GEN_387; // @[ivncontrol4.scala 200:50 201:21]
  wire [31:0] _GEN_392 = _GEN_268 == 32'h5 ? _T_91[31:0] : _GEN_388; // @[ivncontrol4.scala 200:50 202:21]
  wire [31:0] _GEN_393 = _GEN_268 == 32'h5 ? _T_91[31:0] : _GEN_389; // @[ivncontrol4.scala 200:50 203:21]
  wire [31:0] _GEN_394 = _GEN_268 == 32'h5 ? _T_91[31:0] : _GEN_390; // @[ivncontrol4.scala 200:50 204:21]
  wire [31:0] _GEN_395 = _GEN_268 == 32'h5 ? _T_91[31:0] : 32'h9; // @[ivncontrol4.scala 126:18 200:50 205:22]
  wire [31:0] _GEN_396 = _GEN_268 == 32'h6 ? _T_91[31:0] : _GEN_391; // @[ivncontrol4.scala 192:52 193:21]
  wire [31:0] _GEN_397 = _GEN_268 == 32'h6 ? _T_91[31:0] : _GEN_392; // @[ivncontrol4.scala 192:52 194:21]
  wire [31:0] _GEN_398 = _GEN_268 == 32'h6 ? _T_91[31:0] : _GEN_393; // @[ivncontrol4.scala 192:52 195:21]
  wire [31:0] _GEN_399 = _GEN_268 == 32'h6 ? _T_91[31:0] : _GEN_394; // @[ivncontrol4.scala 192:52 196:21]
  wire [31:0] _GEN_400 = _GEN_268 == 32'h6 ? _T_91[31:0] : _GEN_395; // @[ivncontrol4.scala 192:52 197:22]
  wire [31:0] _GEN_401 = _GEN_268 == 32'h6 ? _T_91[31:0] : 32'hc; // @[ivncontrol4.scala 126:18 192:52 198:22]
  wire [31:0] _GEN_402 = _GEN_268 == 32'h7 ? _T_91[31:0] : _GEN_396; // @[ivncontrol4.scala 184:52 185:21]
  wire [31:0] _GEN_403 = _GEN_268 == 32'h7 ? _T_91[31:0] : _GEN_397; // @[ivncontrol4.scala 184:52 186:21]
  wire [31:0] _GEN_404 = _GEN_268 == 32'h7 ? _T_91[31:0] : _GEN_398; // @[ivncontrol4.scala 184:52 187:21]
  wire [31:0] _GEN_405 = _GEN_268 == 32'h7 ? _T_91[31:0] : _GEN_399; // @[ivncontrol4.scala 184:52 188:21]
  wire [31:0] _GEN_406 = _GEN_268 == 32'h7 ? _T_91[31:0] : _GEN_400; // @[ivncontrol4.scala 184:52 189:22]
  wire [31:0] _GEN_407 = _GEN_268 == 32'h7 ? _T_91[31:0] : _GEN_401; // @[ivncontrol4.scala 184:52 190:22]
  wire [31:0] _GEN_408 = _GEN_268 == 32'h7 ? _T_91[31:0] : 32'hb; // @[ivncontrol4.scala 126:18 184:52 191:22]
  wire [31:0] _GEN_409 = _GEN_268 >= 32'h8 ? _T_91[31:0] : _GEN_402; // @[ivncontrol4.scala 174:42 175:21]
  wire [31:0] _GEN_410 = _GEN_268 >= 32'h8 ? _T_91[31:0] : _GEN_403; // @[ivncontrol4.scala 174:42 176:21]
  wire [31:0] _GEN_411 = _GEN_268 >= 32'h8 ? _T_91[31:0] : _GEN_404; // @[ivncontrol4.scala 174:42 177:21]
  wire [31:0] _GEN_412 = _GEN_268 >= 32'h8 ? _T_91[31:0] : _GEN_405; // @[ivncontrol4.scala 174:42 178:21]
  wire [31:0] _GEN_413 = _GEN_268 >= 32'h8 ? _T_91[31:0] : _GEN_406; // @[ivncontrol4.scala 174:42 179:22]
  wire [31:0] _GEN_414 = _GEN_268 >= 32'h8 ? _T_91[31:0] : _GEN_407; // @[ivncontrol4.scala 174:42 180:22]
  wire [31:0] _GEN_415 = _GEN_268 >= 32'h8 ? _T_91[31:0] : _GEN_408; // @[ivncontrol4.scala 174:42 181:22]
  wire [31:0] _GEN_416 = _GEN_268 >= 32'h8 ? _T_91[31:0] : 32'h19; // @[ivncontrol4.scala 126:18 174:42 182:22]
  wire [31:0] _T_127 = 32'h8 - _GEN_268; // @[ivncontrol4.scala 228:18]
  wire [31:0] _i_vn_1_T_15 = 32'h1 + pin; // @[ivncontrol4.scala 229:29]
  wire [31:0] _GEN_529 = _T_127 == 32'h1 ? _i_vn_1_T_15 : _GEN_416; // @[ivncontrol4.scala 269:54 272:22]
  wire [31:0] _GEN_530 = _T_127 == 32'h2 ? _i_vn_1_T_15 : _GEN_415; // @[ivncontrol4.scala 264:54 267:22]
  wire [31:0] _GEN_531 = _T_127 == 32'h2 ? _i_vn_1_T_15 : _GEN_529; // @[ivncontrol4.scala 264:54 268:22]
  wire [31:0] _GEN_532 = _T_127 == 32'h3 ? _i_vn_1_T_15 : _GEN_414; // @[ivncontrol4.scala 257:54 259:22]
  wire [31:0] _GEN_533 = _T_127 == 32'h3 ? _i_vn_1_T_15 : _GEN_530; // @[ivncontrol4.scala 257:54 260:22]
  wire [31:0] _GEN_534 = _T_127 == 32'h3 ? _i_vn_1_T_15 : _GEN_531; // @[ivncontrol4.scala 257:54 261:22]
  wire [31:0] _GEN_535 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_413; // @[ivncontrol4.scala 251:54 253:22]
  wire [31:0] _GEN_536 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_532; // @[ivncontrol4.scala 251:54 254:22]
  wire [31:0] _GEN_537 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_533; // @[ivncontrol4.scala 251:54 255:22]
  wire [31:0] _GEN_538 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_534; // @[ivncontrol4.scala 251:54 256:22]
  wire [31:0] _GEN_539 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_412; // @[ivncontrol4.scala 244:54 246:21]
  wire [31:0] _GEN_540 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_535; // @[ivncontrol4.scala 244:54 247:22]
  wire [31:0] _GEN_541 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_536; // @[ivncontrol4.scala 244:54 248:22]
  wire [31:0] _GEN_542 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_537; // @[ivncontrol4.scala 244:54 249:22]
  wire [31:0] _GEN_543 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_538; // @[ivncontrol4.scala 244:54 250:22]
  wire [31:0] _GEN_544 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_411; // @[ivncontrol4.scala 237:54 238:22]
  wire [31:0] _GEN_545 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_539; // @[ivncontrol4.scala 237:54 239:21]
  wire [31:0] _GEN_546 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_540; // @[ivncontrol4.scala 237:54 240:22]
  wire [31:0] _GEN_547 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_541; // @[ivncontrol4.scala 237:54 241:22]
  wire [31:0] _GEN_548 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_542; // @[ivncontrol4.scala 237:54 242:22]
  wire [31:0] _GEN_549 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_543; // @[ivncontrol4.scala 237:54 243:22]
  wire [31:0] _GEN_550 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_410; // @[ivncontrol4.scala 228:49 229:22]
  wire [31:0] _GEN_551 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_544; // @[ivncontrol4.scala 228:49 230:21]
  wire [31:0] _GEN_552 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_545; // @[ivncontrol4.scala 228:49 231:21]
  wire [31:0] _GEN_553 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_546; // @[ivncontrol4.scala 228:49 232:22]
  wire [31:0] _GEN_554 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_547; // @[ivncontrol4.scala 228:49 233:22]
  wire [31:0] _GEN_555 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_548; // @[ivncontrol4.scala 228:49 234:22]
  wire [31:0] _GEN_556 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_549; // @[ivncontrol4.scala 228:49 235:22]
  wire [31:0] _GEN_574 = 4'h1 == _i_vn_1_T_15[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_575 = 4'h2 == _i_vn_1_T_15[3:0] ? rowcount_2 : _GEN_574; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_576 = 4'h3 == _i_vn_1_T_15[3:0] ? rowcount_3 : _GEN_575; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_577 = 4'h4 == _i_vn_1_T_15[3:0] ? rowcount_4 : _GEN_576; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_578 = 4'h5 == _i_vn_1_T_15[3:0] ? rowcount_5 : _GEN_577; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_579 = 4'h6 == _i_vn_1_T_15[3:0] ? rowcount_6 : _GEN_578; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_580 = 4'h7 == _i_vn_1_T_15[3:0] ? rowcount_7 : _GEN_579; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_581 = 4'h8 == _i_vn_1_T_15[3:0] ? rowcount_8 : _GEN_580; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_582 = 4'h9 == _i_vn_1_T_15[3:0] ? rowcount_9 : _GEN_581; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_583 = 4'ha == _i_vn_1_T_15[3:0] ? rowcount_10 : _GEN_582; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_584 = 4'hb == _i_vn_1_T_15[3:0] ? rowcount_11 : _GEN_583; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_585 = 4'hc == _i_vn_1_T_15[3:0] ? rowcount_12 : _GEN_584; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_586 = 4'hd == _i_vn_1_T_15[3:0] ? rowcount_13 : _GEN_585; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_587 = 4'he == _i_vn_1_T_15[3:0] ? rowcount_14 : _GEN_586; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_588 = 4'hf == _i_vn_1_T_15[3:0] ? rowcount_15 : _GEN_587; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _T_172 = _GEN_268 + _GEN_588; // @[ivncontrol4.scala 275:41]
  wire [31:0] _T_174 = 32'h8 - _T_172; // @[ivncontrol4.scala 275:18]
  wire [31:0] _i_vn_1_T_17 = 32'h2 + pin; // @[ivncontrol4.scala 276:29]
  wire [31:0] _GEN_781 = _T_174 == 32'h1 ? _i_vn_1_T_17 : _GEN_556; // @[ivncontrol4.scala 318:78 321:22]
  wire [31:0] _GEN_782 = _T_174 == 32'h2 ? _i_vn_1_T_17 : _GEN_555; // @[ivncontrol4.scala 312:76 315:22]
  wire [31:0] _GEN_783 = _T_174 == 32'h2 ? _i_vn_1_T_17 : _GEN_781; // @[ivncontrol4.scala 312:76 316:22]
  wire [31:0] _GEN_784 = _T_174 == 32'h3 ? _i_vn_1_T_17 : _GEN_554; // @[ivncontrol4.scala 305:78 307:23]
  wire [31:0] _GEN_785 = _T_174 == 32'h3 ? _i_vn_1_T_17 : _GEN_782; // @[ivncontrol4.scala 305:78 308:22]
  wire [31:0] _GEN_786 = _T_174 == 32'h3 ? _i_vn_1_T_17 : _GEN_783; // @[ivncontrol4.scala 305:78 309:22]
  wire [31:0] _GEN_787 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_553; // @[ivncontrol4.scala 299:78 301:22]
  wire [31:0] _GEN_788 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_784; // @[ivncontrol4.scala 299:78 302:22]
  wire [31:0] _GEN_789 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_785; // @[ivncontrol4.scala 299:78 303:22]
  wire [31:0] _GEN_790 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_786; // @[ivncontrol4.scala 299:78 304:22]
  wire [31:0] _GEN_791 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_552; // @[ivncontrol4.scala 292:76 294:23]
  wire [31:0] _GEN_792 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_787; // @[ivncontrol4.scala 292:76 295:22]
  wire [31:0] _GEN_793 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_788; // @[ivncontrol4.scala 292:76 296:22]
  wire [31:0] _GEN_794 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_789; // @[ivncontrol4.scala 292:76 297:22]
  wire [31:0] _GEN_795 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_790; // @[ivncontrol4.scala 292:76 298:22]
  wire [31:0] _GEN_796 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_551; // @[ivncontrol4.scala 284:77 286:22]
  wire [31:0] _GEN_797 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_791; // @[ivncontrol4.scala 284:77 287:21]
  wire [31:0] _GEN_798 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_792; // @[ivncontrol4.scala 284:77 288:22]
  wire [31:0] _GEN_799 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_793; // @[ivncontrol4.scala 284:77 289:22]
  wire [31:0] _GEN_800 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_794; // @[ivncontrol4.scala 284:77 290:22]
  wire [31:0] _GEN_801 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_795; // @[ivncontrol4.scala 284:77 291:22]
  wire [31:0] _GEN_802 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_550; // @[ivncontrol4.scala 275:73 276:22]
  wire [31:0] _GEN_803 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_796; // @[ivncontrol4.scala 275:73 277:21]
  wire [31:0] _GEN_804 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_797; // @[ivncontrol4.scala 275:73 278:21]
  wire [31:0] _GEN_805 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_798; // @[ivncontrol4.scala 275:73 279:22]
  wire [31:0] _GEN_806 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_799; // @[ivncontrol4.scala 275:73 280:22]
  wire [31:0] _GEN_807 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_800; // @[ivncontrol4.scala 275:73 281:22]
  wire [31:0] _GEN_808 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_801; // @[ivncontrol4.scala 275:73 282:22]
  wire [31:0] _GEN_842 = 4'h1 == _i_vn_1_T_17[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_843 = 4'h2 == _i_vn_1_T_17[3:0] ? rowcount_2 : _GEN_842; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_844 = 4'h3 == _i_vn_1_T_17[3:0] ? rowcount_3 : _GEN_843; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_845 = 4'h4 == _i_vn_1_T_17[3:0] ? rowcount_4 : _GEN_844; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_846 = 4'h5 == _i_vn_1_T_17[3:0] ? rowcount_5 : _GEN_845; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_847 = 4'h6 == _i_vn_1_T_17[3:0] ? rowcount_6 : _GEN_846; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_848 = 4'h7 == _i_vn_1_T_17[3:0] ? rowcount_7 : _GEN_847; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_849 = 4'h8 == _i_vn_1_T_17[3:0] ? rowcount_8 : _GEN_848; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_850 = 4'h9 == _i_vn_1_T_17[3:0] ? rowcount_9 : _GEN_849; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_851 = 4'ha == _i_vn_1_T_17[3:0] ? rowcount_10 : _GEN_850; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_852 = 4'hb == _i_vn_1_T_17[3:0] ? rowcount_11 : _GEN_851; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_853 = 4'hc == _i_vn_1_T_17[3:0] ? rowcount_12 : _GEN_852; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_854 = 4'hd == _i_vn_1_T_17[3:0] ? rowcount_13 : _GEN_853; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_855 = 4'he == _i_vn_1_T_17[3:0] ? rowcount_14 : _GEN_854; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_856 = 4'hf == _i_vn_1_T_17[3:0] ? rowcount_15 : _GEN_855; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _T_254 = _T_172 + _GEN_856; // @[ivncontrol4.scala 326:62]
  wire [31:0] _T_256 = 32'h8 - _T_254; // @[ivncontrol4.scala 326:17]
  wire [31:0] _i_vn_1_T_19 = 32'h3 + pin; // @[ivncontrol4.scala 327:29]
  wire [31:0] _GEN_1145 = _T_256 == 32'h1 ? _i_vn_1_T_19 : _GEN_808; // @[ivncontrol4.scala 369:100 372:22]
  wire [31:0] _GEN_1146 = _T_256 == 32'h2 ? _i_vn_1_T_19 : _GEN_807; // @[ivncontrol4.scala 363:98 366:22]
  wire [31:0] _GEN_1147 = _T_256 == 32'h2 ? _i_vn_1_T_19 : _GEN_1145; // @[ivncontrol4.scala 363:98 367:22]
  wire [31:0] _GEN_1148 = _T_256 == 32'h3 ? _i_vn_1_T_19 : _GEN_806; // @[ivncontrol4.scala 356:100 358:23]
  wire [31:0] _GEN_1149 = _T_256 == 32'h3 ? _i_vn_1_T_19 : _GEN_1146; // @[ivncontrol4.scala 356:100 359:22]
  wire [31:0] _GEN_1150 = _T_256 == 32'h3 ? _i_vn_1_T_19 : _GEN_1147; // @[ivncontrol4.scala 356:100 360:22]
  wire [31:0] _GEN_1151 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_805; // @[ivncontrol4.scala 350:100 352:22]
  wire [31:0] _GEN_1152 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_1148; // @[ivncontrol4.scala 350:100 353:22]
  wire [31:0] _GEN_1153 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_1149; // @[ivncontrol4.scala 350:100 354:22]
  wire [31:0] _GEN_1154 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_1150; // @[ivncontrol4.scala 350:100 355:22]
  wire [31:0] _GEN_1155 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_804; // @[ivncontrol4.scala 343:98 345:23]
  wire [31:0] _GEN_1156 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1151; // @[ivncontrol4.scala 343:98 346:22]
  wire [31:0] _GEN_1157 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1152; // @[ivncontrol4.scala 343:98 347:22]
  wire [31:0] _GEN_1158 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1153; // @[ivncontrol4.scala 343:98 348:22]
  wire [31:0] _GEN_1159 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1154; // @[ivncontrol4.scala 343:98 349:22]
  wire [31:0] _GEN_1160 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_803; // @[ivncontrol4.scala 335:99 337:22]
  wire [31:0] _GEN_1161 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1155; // @[ivncontrol4.scala 335:99 338:21]
  wire [31:0] _GEN_1162 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1156; // @[ivncontrol4.scala 335:99 339:22]
  wire [31:0] _GEN_1163 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1157; // @[ivncontrol4.scala 335:99 340:22]
  wire [31:0] _GEN_1164 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1158; // @[ivncontrol4.scala 335:99 341:22]
  wire [31:0] _GEN_1165 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1159; // @[ivncontrol4.scala 335:99 342:22]
  wire [31:0] _GEN_1166 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_802; // @[ivncontrol4.scala 326:94 327:22]
  wire [31:0] _GEN_1167 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1160; // @[ivncontrol4.scala 326:94 328:21]
  wire [31:0] _GEN_1168 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1161; // @[ivncontrol4.scala 326:94 329:21]
  wire [31:0] _GEN_1169 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1162; // @[ivncontrol4.scala 326:94 330:22]
  wire [31:0] _GEN_1170 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1163; // @[ivncontrol4.scala 326:94 331:22]
  wire [31:0] _GEN_1171 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1164; // @[ivncontrol4.scala 326:94 332:22]
  wire [31:0] _GEN_1172 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1165; // @[ivncontrol4.scala 326:94 333:22]
  wire [31:0] _GEN_1222 = 4'h1 == _i_vn_1_T_19[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1223 = 4'h2 == _i_vn_1_T_19[3:0] ? rowcount_2 : _GEN_1222; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1224 = 4'h3 == _i_vn_1_T_19[3:0] ? rowcount_3 : _GEN_1223; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1225 = 4'h4 == _i_vn_1_T_19[3:0] ? rowcount_4 : _GEN_1224; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1226 = 4'h5 == _i_vn_1_T_19[3:0] ? rowcount_5 : _GEN_1225; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1227 = 4'h6 == _i_vn_1_T_19[3:0] ? rowcount_6 : _GEN_1226; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1228 = 4'h7 == _i_vn_1_T_19[3:0] ? rowcount_7 : _GEN_1227; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1229 = 4'h8 == _i_vn_1_T_19[3:0] ? rowcount_8 : _GEN_1228; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1230 = 4'h9 == _i_vn_1_T_19[3:0] ? rowcount_9 : _GEN_1229; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1231 = 4'ha == _i_vn_1_T_19[3:0] ? rowcount_10 : _GEN_1230; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1232 = 4'hb == _i_vn_1_T_19[3:0] ? rowcount_11 : _GEN_1231; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1233 = 4'hc == _i_vn_1_T_19[3:0] ? rowcount_12 : _GEN_1232; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1234 = 4'hd == _i_vn_1_T_19[3:0] ? rowcount_13 : _GEN_1233; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1235 = 4'he == _i_vn_1_T_19[3:0] ? rowcount_14 : _GEN_1234; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1236 = 4'hf == _i_vn_1_T_19[3:0] ? rowcount_15 : _GEN_1235; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _T_371 = _T_254 + _GEN_1236; // @[ivncontrol4.scala 376:86]
  wire [31:0] _T_373 = 32'h8 - _T_371; // @[ivncontrol4.scala 376:19]
  wire [31:0] _i_vn_1_T_21 = 32'h4 + pin; // @[ivncontrol4.scala 377:29]
  wire [31:0] _GEN_1621 = _T_373 == 32'h1 ? _i_vn_1_T_21 : _GEN_1172; // @[ivncontrol4.scala 419:122 422:22]
  wire [31:0] _GEN_1622 = _T_373 == 32'h2 ? _i_vn_1_T_21 : _GEN_1171; // @[ivncontrol4.scala 413:121 416:22]
  wire [31:0] _GEN_1623 = _T_373 == 32'h2 ? _i_vn_1_T_21 : _GEN_1621; // @[ivncontrol4.scala 413:121 417:22]
  wire [31:0] _GEN_1624 = _T_373 == 32'h3 ? _i_vn_1_T_21 : _GEN_1170; // @[ivncontrol4.scala 406:123 408:23]
  wire [31:0] _GEN_1625 = _T_373 == 32'h3 ? _i_vn_1_T_21 : _GEN_1622; // @[ivncontrol4.scala 406:123 409:22]
  wire [31:0] _GEN_1626 = _T_373 == 32'h3 ? _i_vn_1_T_21 : _GEN_1623; // @[ivncontrol4.scala 406:123 410:22]
  wire [31:0] _GEN_1627 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1169; // @[ivncontrol4.scala 400:122 402:22]
  wire [31:0] _GEN_1628 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1624; // @[ivncontrol4.scala 400:122 403:22]
  wire [31:0] _GEN_1629 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1625; // @[ivncontrol4.scala 400:122 404:22]
  wire [31:0] _GEN_1630 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1626; // @[ivncontrol4.scala 400:122 405:22]
  wire [31:0] _GEN_1631 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1168; // @[ivncontrol4.scala 393:121 395:23]
  wire [31:0] _GEN_1632 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1627; // @[ivncontrol4.scala 393:121 396:22]
  wire [31:0] _GEN_1633 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1628; // @[ivncontrol4.scala 393:121 397:22]
  wire [31:0] _GEN_1634 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1629; // @[ivncontrol4.scala 393:121 398:22]
  wire [31:0] _GEN_1635 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1630; // @[ivncontrol4.scala 393:121 399:22]
  wire [31:0] _GEN_1636 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1167; // @[ivncontrol4.scala 385:121 387:22]
  wire [31:0] _GEN_1637 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1631; // @[ivncontrol4.scala 385:121 388:21]
  wire [31:0] _GEN_1638 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1632; // @[ivncontrol4.scala 385:121 389:22]
  wire [31:0] _GEN_1639 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1633; // @[ivncontrol4.scala 385:121 390:22]
  wire [31:0] _GEN_1640 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1634; // @[ivncontrol4.scala 385:121 391:22]
  wire [31:0] _GEN_1641 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1635; // @[ivncontrol4.scala 385:121 392:22]
  wire [31:0] _GEN_1642 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1166; // @[ivncontrol4.scala 376:118 377:22]
  wire [31:0] _GEN_1643 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1636; // @[ivncontrol4.scala 376:118 378:21]
  wire [31:0] _GEN_1644 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1637; // @[ivncontrol4.scala 376:118 379:21]
  wire [31:0] _GEN_1645 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1638; // @[ivncontrol4.scala 376:118 380:22]
  wire [31:0] _GEN_1646 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1639; // @[ivncontrol4.scala 376:118 381:22]
  wire [31:0] _GEN_1647 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1640; // @[ivncontrol4.scala 376:118 382:22]
  wire [31:0] _GEN_1648 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1641; // @[ivncontrol4.scala 376:118 383:22]
  wire [31:0] _GEN_1714 = 4'h1 == _i_vn_1_T_21[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1715 = 4'h2 == _i_vn_1_T_21[3:0] ? rowcount_2 : _GEN_1714; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1716 = 4'h3 == _i_vn_1_T_21[3:0] ? rowcount_3 : _GEN_1715; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1717 = 4'h4 == _i_vn_1_T_21[3:0] ? rowcount_4 : _GEN_1716; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1718 = 4'h5 == _i_vn_1_T_21[3:0] ? rowcount_5 : _GEN_1717; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1719 = 4'h6 == _i_vn_1_T_21[3:0] ? rowcount_6 : _GEN_1718; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1720 = 4'h7 == _i_vn_1_T_21[3:0] ? rowcount_7 : _GEN_1719; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1721 = 4'h8 == _i_vn_1_T_21[3:0] ? rowcount_8 : _GEN_1720; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1722 = 4'h9 == _i_vn_1_T_21[3:0] ? rowcount_9 : _GEN_1721; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1723 = 4'ha == _i_vn_1_T_21[3:0] ? rowcount_10 : _GEN_1722; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1724 = 4'hb == _i_vn_1_T_21[3:0] ? rowcount_11 : _GEN_1723; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1725 = 4'hc == _i_vn_1_T_21[3:0] ? rowcount_12 : _GEN_1724; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1726 = 4'hd == _i_vn_1_T_21[3:0] ? rowcount_13 : _GEN_1725; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1727 = 4'he == _i_vn_1_T_21[3:0] ? rowcount_14 : _GEN_1726; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1728 = 4'hf == _i_vn_1_T_21[3:0] ? rowcount_15 : _GEN_1727; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _T_523 = _T_371 + _GEN_1728; // @[ivncontrol4.scala 426:108]
  wire [31:0] _T_525 = 32'h8 - _T_523; // @[ivncontrol4.scala 426:19]
  wire [31:0] _i_vn_1_T_23 = 32'h5 + pin; // @[ivncontrol4.scala 427:29]
  wire [31:0] _GEN_2209 = _T_525 == 32'h1 ? _i_vn_1_T_23 : _GEN_1648; // @[ivncontrol4.scala 469:144 472:22]
  wire [31:0] _GEN_2210 = _T_525 == 32'h2 ? _i_vn_1_T_23 : _GEN_1647; // @[ivncontrol4.scala 463:143 466:22]
  wire [31:0] _GEN_2211 = _T_525 == 32'h2 ? _i_vn_1_T_23 : _GEN_2209; // @[ivncontrol4.scala 463:143 467:22]
  wire [31:0] _GEN_2212 = _T_525 == 32'h3 ? _i_vn_1_T_23 : _GEN_1646; // @[ivncontrol4.scala 456:145 458:23]
  wire [31:0] _GEN_2213 = _T_525 == 32'h3 ? _i_vn_1_T_23 : _GEN_2210; // @[ivncontrol4.scala 456:145 459:22]
  wire [31:0] _GEN_2214 = _T_525 == 32'h3 ? _i_vn_1_T_23 : _GEN_2211; // @[ivncontrol4.scala 456:145 460:22]
  wire [31:0] _GEN_2215 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_1645; // @[ivncontrol4.scala 450:143 452:22]
  wire [31:0] _GEN_2216 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_2212; // @[ivncontrol4.scala 450:143 453:22]
  wire [31:0] _GEN_2217 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_2213; // @[ivncontrol4.scala 450:143 454:22]
  wire [31:0] _GEN_2218 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_2214; // @[ivncontrol4.scala 450:143 455:22]
  wire [31:0] _GEN_2219 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_1644; // @[ivncontrol4.scala 443:143 445:23]
  wire [31:0] _GEN_2220 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2215; // @[ivncontrol4.scala 443:143 446:22]
  wire [31:0] _GEN_2221 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2216; // @[ivncontrol4.scala 443:143 447:22]
  wire [31:0] _GEN_2222 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2217; // @[ivncontrol4.scala 443:143 448:22]
  wire [31:0] _GEN_2223 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2218; // @[ivncontrol4.scala 443:143 449:22]
  wire [31:0] _GEN_2224 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_1643; // @[ivncontrol4.scala 435:143 437:22]
  wire [31:0] _GEN_2225 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2219; // @[ivncontrol4.scala 435:143 438:21]
  wire [31:0] _GEN_2226 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2220; // @[ivncontrol4.scala 435:143 439:22]
  wire [31:0] _GEN_2227 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2221; // @[ivncontrol4.scala 435:143 440:22]
  wire [31:0] _GEN_2228 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2222; // @[ivncontrol4.scala 435:143 441:22]
  wire [31:0] _GEN_2229 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2223; // @[ivncontrol4.scala 435:143 442:22]
  wire [31:0] _GEN_2230 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_1642; // @[ivncontrol4.scala 426:140 427:22]
  wire [31:0] _GEN_2231 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2224; // @[ivncontrol4.scala 426:140 428:21]
  wire [31:0] _GEN_2232 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2225; // @[ivncontrol4.scala 426:140 429:21]
  wire [31:0] _GEN_2233 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2226; // @[ivncontrol4.scala 426:140 430:22]
  wire [31:0] _GEN_2234 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2227; // @[ivncontrol4.scala 426:140 431:22]
  wire [31:0] _GEN_2235 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2228; // @[ivncontrol4.scala 426:140 432:22]
  wire [31:0] _GEN_2236 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2229; // @[ivncontrol4.scala 426:140 433:22]
  wire [31:0] _GEN_2318 = 4'h1 == _i_vn_1_T_23[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2319 = 4'h2 == _i_vn_1_T_23[3:0] ? rowcount_2 : _GEN_2318; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2320 = 4'h3 == _i_vn_1_T_23[3:0] ? rowcount_3 : _GEN_2319; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2321 = 4'h4 == _i_vn_1_T_23[3:0] ? rowcount_4 : _GEN_2320; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2322 = 4'h5 == _i_vn_1_T_23[3:0] ? rowcount_5 : _GEN_2321; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2323 = 4'h6 == _i_vn_1_T_23[3:0] ? rowcount_6 : _GEN_2322; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2324 = 4'h7 == _i_vn_1_T_23[3:0] ? rowcount_7 : _GEN_2323; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2325 = 4'h8 == _i_vn_1_T_23[3:0] ? rowcount_8 : _GEN_2324; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2326 = 4'h9 == _i_vn_1_T_23[3:0] ? rowcount_9 : _GEN_2325; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2327 = 4'ha == _i_vn_1_T_23[3:0] ? rowcount_10 : _GEN_2326; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2328 = 4'hb == _i_vn_1_T_23[3:0] ? rowcount_11 : _GEN_2327; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2329 = 4'hc == _i_vn_1_T_23[3:0] ? rowcount_12 : _GEN_2328; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2330 = 4'hd == _i_vn_1_T_23[3:0] ? rowcount_13 : _GEN_2329; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2331 = 4'he == _i_vn_1_T_23[3:0] ? rowcount_14 : _GEN_2330; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2332 = 4'hf == _i_vn_1_T_23[3:0] ? rowcount_15 : _GEN_2331; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _T_710 = _T_523 + _GEN_2332; // @[ivncontrol4.scala 477:130]
  wire [31:0] _T_712 = 32'h8 - _T_710; // @[ivncontrol4.scala 477:19]
  wire [31:0] _i_vn_1_T_25 = 32'h6 + pin; // @[ivncontrol4.scala 478:29]
  wire [31:0] _GEN_2909 = _T_712 == 32'h1 ? _i_vn_1_T_25 : _GEN_2236; // @[ivncontrol4.scala 520:166 523:22]
  wire [31:0] _GEN_2910 = _T_712 == 32'h2 ? _i_vn_1_T_25 : _GEN_2235; // @[ivncontrol4.scala 514:166 517:22]
  wire [31:0] _GEN_2911 = _T_712 == 32'h2 ? _i_vn_1_T_25 : _GEN_2909; // @[ivncontrol4.scala 514:166 518:22]
  wire [31:0] _GEN_2912 = _T_712 == 32'h3 ? _i_vn_1_T_25 : _GEN_2234; // @[ivncontrol4.scala 507:168 509:23]
  wire [31:0] _GEN_2913 = _T_712 == 32'h3 ? _i_vn_1_T_25 : _GEN_2910; // @[ivncontrol4.scala 507:168 510:22]
  wire [31:0] _GEN_2914 = _T_712 == 32'h3 ? _i_vn_1_T_25 : _GEN_2911; // @[ivncontrol4.scala 507:168 511:22]
  wire [31:0] _GEN_2915 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2233; // @[ivncontrol4.scala 501:166 503:22]
  wire [31:0] _GEN_2916 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2912; // @[ivncontrol4.scala 501:166 504:22]
  wire [31:0] _GEN_2917 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2913; // @[ivncontrol4.scala 501:166 505:22]
  wire [31:0] _GEN_2918 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2914; // @[ivncontrol4.scala 501:166 506:22]
  wire [31:0] _GEN_2919 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2232; // @[ivncontrol4.scala 494:166 496:23]
  wire [31:0] _GEN_2920 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2915; // @[ivncontrol4.scala 494:166 497:22]
  wire [31:0] _GEN_2921 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2916; // @[ivncontrol4.scala 494:166 498:22]
  wire [31:0] _GEN_2922 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2917; // @[ivncontrol4.scala 494:166 499:22]
  wire [31:0] _GEN_2923 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2918; // @[ivncontrol4.scala 494:166 500:22]
  wire [31:0] _GEN_2924 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2231; // @[ivncontrol4.scala 486:166 488:22]
  wire [31:0] _GEN_2925 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2919; // @[ivncontrol4.scala 486:166 489:21]
  wire [31:0] _GEN_2926 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2920; // @[ivncontrol4.scala 486:166 490:22]
  wire [31:0] _GEN_2927 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2921; // @[ivncontrol4.scala 486:166 491:22]
  wire [31:0] _GEN_2928 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2922; // @[ivncontrol4.scala 486:166 492:22]
  wire [31:0] _GEN_2929 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2923; // @[ivncontrol4.scala 486:166 493:22]
  wire [31:0] _GEN_2930 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2230; // @[ivncontrol4.scala 477:162 478:22]
  wire [31:0] _GEN_2931 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2924; // @[ivncontrol4.scala 477:162 479:21]
  wire [31:0] _GEN_2932 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2925; // @[ivncontrol4.scala 477:162 480:21]
  wire [31:0] _GEN_2933 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2926; // @[ivncontrol4.scala 477:162 481:22]
  wire [31:0] _GEN_2934 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2927; // @[ivncontrol4.scala 477:162 482:22]
  wire [31:0] _GEN_2935 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2928; // @[ivncontrol4.scala 477:162 483:22]
  wire [31:0] _GEN_2936 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2929; // @[ivncontrol4.scala 477:162 484:22]
  wire [31:0] _GEN_3034 = 4'h1 == _i_vn_1_T_25[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3035 = 4'h2 == _i_vn_1_T_25[3:0] ? rowcount_2 : _GEN_3034; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3036 = 4'h3 == _i_vn_1_T_25[3:0] ? rowcount_3 : _GEN_3035; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3037 = 4'h4 == _i_vn_1_T_25[3:0] ? rowcount_4 : _GEN_3036; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3038 = 4'h5 == _i_vn_1_T_25[3:0] ? rowcount_5 : _GEN_3037; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3039 = 4'h6 == _i_vn_1_T_25[3:0] ? rowcount_6 : _GEN_3038; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3040 = 4'h7 == _i_vn_1_T_25[3:0] ? rowcount_7 : _GEN_3039; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3041 = 4'h8 == _i_vn_1_T_25[3:0] ? rowcount_8 : _GEN_3040; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3042 = 4'h9 == _i_vn_1_T_25[3:0] ? rowcount_9 : _GEN_3041; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3043 = 4'ha == _i_vn_1_T_25[3:0] ? rowcount_10 : _GEN_3042; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3044 = 4'hb == _i_vn_1_T_25[3:0] ? rowcount_11 : _GEN_3043; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3045 = 4'hc == _i_vn_1_T_25[3:0] ? rowcount_12 : _GEN_3044; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3046 = 4'hd == _i_vn_1_T_25[3:0] ? rowcount_13 : _GEN_3045; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3047 = 4'he == _i_vn_1_T_25[3:0] ? rowcount_14 : _GEN_3046; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3048 = 4'hf == _i_vn_1_T_25[3:0] ? rowcount_15 : _GEN_3047; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _T_932 = _T_710 + _GEN_3048; // @[ivncontrol4.scala 528:152]
  wire [31:0] _T_934 = 32'h8 - _T_932; // @[ivncontrol4.scala 528:19]
  wire [31:0] _i_vn_1_T_27 = 32'h7 + pin; // @[ivncontrol4.scala 529:29]
  wire [31:0] _GEN_3721 = _T_934 == 32'h1 ? _i_vn_1_T_27 : _GEN_2936; // @[ivncontrol4.scala 571:188 574:22]
  wire [31:0] _GEN_3722 = _T_934 == 32'h2 ? _i_vn_1_T_27 : _GEN_2935; // @[ivncontrol4.scala 565:188 568:22]
  wire [31:0] _GEN_3723 = _T_934 == 32'h2 ? _i_vn_1_T_27 : _GEN_3721; // @[ivncontrol4.scala 565:188 569:22]
  wire [31:0] _GEN_3724 = _T_934 == 32'h3 ? _i_vn_1_T_27 : _GEN_2934; // @[ivncontrol4.scala 558:190 560:23]
  wire [31:0] _GEN_3725 = _T_934 == 32'h3 ? _i_vn_1_T_27 : _GEN_3722; // @[ivncontrol4.scala 558:190 561:22]
  wire [31:0] _GEN_3726 = _T_934 == 32'h3 ? _i_vn_1_T_27 : _GEN_3723; // @[ivncontrol4.scala 558:190 562:22]
  wire [31:0] _GEN_3727 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_2933; // @[ivncontrol4.scala 552:188 554:22]
  wire [31:0] _GEN_3728 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_3724; // @[ivncontrol4.scala 552:188 555:22]
  wire [31:0] _GEN_3729 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_3725; // @[ivncontrol4.scala 552:188 556:22]
  wire [31:0] _GEN_3730 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_3726; // @[ivncontrol4.scala 552:188 557:22]
  wire [31:0] _GEN_3731 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_2932; // @[ivncontrol4.scala 545:188 547:23]
  wire [31:0] _GEN_3732 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3727; // @[ivncontrol4.scala 545:188 548:22]
  wire [31:0] _GEN_3733 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3728; // @[ivncontrol4.scala 545:188 549:22]
  wire [31:0] _GEN_3734 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3729; // @[ivncontrol4.scala 545:188 550:22]
  wire [31:0] _GEN_3735 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3730; // @[ivncontrol4.scala 545:188 551:22]
  wire [31:0] _GEN_3736 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_2931; // @[ivncontrol4.scala 537:188 539:22]
  wire [31:0] _GEN_3737 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3731; // @[ivncontrol4.scala 537:188 540:21]
  wire [31:0] _GEN_3738 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3732; // @[ivncontrol4.scala 537:188 541:22]
  wire [31:0] _GEN_3739 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3733; // @[ivncontrol4.scala 537:188 542:22]
  wire [31:0] _GEN_3740 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3734; // @[ivncontrol4.scala 537:188 543:22]
  wire [31:0] _GEN_3741 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3735; // @[ivncontrol4.scala 537:188 544:22]
  wire [31:0] _GEN_3742 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_2930; // @[ivncontrol4.scala 528:184 529:22]
  wire [31:0] _GEN_3743 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3736; // @[ivncontrol4.scala 528:184 530:21]
  wire [31:0] _GEN_3744 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3737; // @[ivncontrol4.scala 528:184 531:21]
  wire [31:0] _GEN_3745 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3738; // @[ivncontrol4.scala 528:184 532:22]
  wire [31:0] _GEN_3746 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3739; // @[ivncontrol4.scala 528:184 533:22]
  wire [31:0] _GEN_3747 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3740; // @[ivncontrol4.scala 528:184 534:22]
  wire [31:0] _GEN_3748 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3741; // @[ivncontrol4.scala 528:184 535:22]
  wire [31:0] _GEN_3749 = _GEN_244 ? _GEN_409 : 32'h18; // @[ivncontrol4.scala 125:17 172:28]
  wire [31:0] _GEN_3750 = _GEN_244 ? _GEN_3742 : 32'h1e; // @[ivncontrol4.scala 125:17 172:28]
  wire [31:0] _GEN_3751 = _GEN_244 ? _GEN_3743 : 32'h1e; // @[ivncontrol4.scala 125:17 172:28]
  wire [31:0] _GEN_3752 = _GEN_244 ? _GEN_3744 : 32'h14; // @[ivncontrol4.scala 125:17 172:28]
  wire [31:0] _GEN_3753 = _GEN_244 ? _GEN_3745 : 32'h9; // @[ivncontrol4.scala 126:18 172:28]
  wire [31:0] _GEN_3754 = _GEN_244 ? _GEN_3746 : 32'hc; // @[ivncontrol4.scala 126:18 172:28]
  wire [31:0] _GEN_3755 = _GEN_244 ? _GEN_3747 : 32'hb; // @[ivncontrol4.scala 126:18 172:28]
  wire [31:0] _GEN_3756 = _GEN_244 ? _GEN_3748 : 32'h19; // @[ivncontrol4.scala 126:18 172:28]
  wire [31:0] _GEN_4137 = reset ? 32'h0 : _GEN_3749; // @[ivncontrol4.scala 16:{23,23}]
  wire [31:0] _GEN_4138 = reset ? 32'h0 : _GEN_3750; // @[ivncontrol4.scala 16:{23,23}]
  wire [31:0] _GEN_4139 = reset ? 32'h0 : _GEN_3751; // @[ivncontrol4.scala 16:{23,23}]
  wire [31:0] _GEN_4140 = reset ? 32'h0 : _GEN_3752; // @[ivncontrol4.scala 16:{23,23}]
  wire [31:0] _GEN_4141 = reset ? 32'h0 : _GEN_3753; // @[ivncontrol4.scala 17:{24,24}]
  wire [31:0] _GEN_4142 = reset ? 32'h0 : _GEN_3754; // @[ivncontrol4.scala 17:{24,24}]
  wire [31:0] _GEN_4143 = reset ? 32'h0 : _GEN_3755; // @[ivncontrol4.scala 17:{24,24}]
  wire [31:0] _GEN_4144 = reset ? 32'h0 : _GEN_3756; // @[ivncontrol4.scala 17:{24,24}]
  assign io_o_vn_0 = i_vn_0; // @[ivncontrol4.scala 121:13]
  assign io_o_vn_1 = i_vn_1; // @[ivncontrol4.scala 121:13]
  assign io_o_vn_2 = i_vn_2; // @[ivncontrol4.scala 121:13]
  assign io_o_vn_3 = i_vn_3; // @[ivncontrol4.scala 121:13]
  assign io_o_vn2_0 = i_vn2_0; // @[ivncontrol4.scala 122:14]
  assign io_o_vn2_1 = i_vn2_1; // @[ivncontrol4.scala 122:14]
  assign io_o_vn2_2 = i_vn2_2; // @[ivncontrol4.scala 122:14]
  assign io_o_vn2_3 = i_vn2_3; // @[ivncontrol4.scala 122:14]
  always @(posedge clock) begin
    i_vn_0 <= _GEN_4137[4:0]; // @[ivncontrol4.scala 16:{23,23}]
    i_vn_1 <= _GEN_4138[4:0]; // @[ivncontrol4.scala 16:{23,23}]
    i_vn_2 <= _GEN_4139[4:0]; // @[ivncontrol4.scala 16:{23,23}]
    i_vn_3 <= _GEN_4140[4:0]; // @[ivncontrol4.scala 16:{23,23}]
    i_vn2_0 <= _GEN_4141[4:0]; // @[ivncontrol4.scala 17:{24,24}]
    i_vn2_1 <= _GEN_4142[4:0]; // @[ivncontrol4.scala 17:{24,24}]
    i_vn2_2 <= _GEN_4143[4:0]; // @[ivncontrol4.scala 17:{24,24}]
    i_vn2_3 <= _GEN_4144[4:0]; // @[ivncontrol4.scala 17:{24,24}]
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_0 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_0 <= count_0; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_1 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_1 <= count_1; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_2 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_2 <= count_2; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_3 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_3 <= count_3; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_4 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_4 <= count_4; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_5 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_5 <= count_5; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_6 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_6 <= count_6; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_7 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_7 <= count_7; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_8 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_8 <= 32'h0; // @[ivncontrol4.scala 81:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_9 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_9 <= 32'h0; // @[ivncontrol4.scala 81:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_10 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_10 <= 32'h0; // @[ivncontrol4.scala 81:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_11 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_11 <= 32'h0; // @[ivncontrol4.scala 81:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_12 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_12 <= 32'h0; // @[ivncontrol4.scala 81:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_13 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_13 <= 32'h0; // @[ivncontrol4.scala 81:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_14 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_14 <= 32'h0; // @[ivncontrol4.scala 81:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_15 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end
    if (reset) begin // @[ivncontrol4.scala 31:22]
      pin <= 32'h0; // @[ivncontrol4.scala 31:22]
    end else if (_T_72 & rowcount_6 == 32'h0 & rowcount_7 != 32'h0) begin // @[ivncontrol4.scala 166:192]
      pin <= 32'h7; // @[ivncontrol4.scala 167:13]
    end else if (_T_59 & rowcount_5 == 32'h0 & rowcount_6 != 32'h0) begin // @[ivncontrol4.scala 163:169]
      pin <= 32'h6; // @[ivncontrol4.scala 164:13]
    end else if (_T_48 & rowcount_4 == 32'h0 & rowcount_5 != 32'h0) begin // @[ivncontrol4.scala 160:146]
      pin <= 32'h5; // @[ivncontrol4.scala 161:13]
    end else begin
      pin <= _GEN_249;
    end
    if (reset) begin // @[ivncontrol4.scala 35:20]
      i <= 32'h0; // @[ivncontrol4.scala 35:20]
    end else if (i < 32'h7 & _k_T_1) begin // @[ivncontrol4.scala 103:74]
      i <= _i_T_1; // @[ivncontrol4.scala 104:11]
    end
    if (reset) begin // @[ivncontrol4.scala 36:20]
      j <= 32'h0; // @[ivncontrol4.scala 36:20]
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 107:71]
      j <= _j_T_1; // @[ivncontrol4.scala 108:11]
    end else if (!(_k_T_2)) begin // @[ivncontrol4.scala 110:81]
      j <= 32'h0; // @[ivncontrol4.scala 114:11]
    end
    if (3'h0 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h0 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h0 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h0 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h0 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h0 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h0 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h0 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h0 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_0 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h1 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_1 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h2 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_2 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h3 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_3 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h4 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_4 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h5 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_5 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h6 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_6 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h7 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_7 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  i_vn_0 = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  i_vn_1 = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  i_vn_2 = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  i_vn_3 = _RAND_3[4:0];
  _RAND_4 = {1{`RANDOM}};
  i_vn2_0 = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  i_vn2_1 = _RAND_5[4:0];
  _RAND_6 = {1{`RANDOM}};
  i_vn2_2 = _RAND_6[4:0];
  _RAND_7 = {1{`RANDOM}};
  i_vn2_3 = _RAND_7[4:0];
  _RAND_8 = {1{`RANDOM}};
  rowcount_0 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  rowcount_1 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  rowcount_2 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  rowcount_3 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  rowcount_4 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  rowcount_5 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  rowcount_6 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  rowcount_7 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  rowcount_8 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  rowcount_9 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  rowcount_10 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  rowcount_11 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  rowcount_12 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  rowcount_13 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  rowcount_14 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  rowcount_15 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  pin = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  i = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  j = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  mat_0_0 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  mat_0_1 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  mat_0_2 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  mat_0_3 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  mat_0_4 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  mat_0_5 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  mat_0_6 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  mat_0_7 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  mat_1_0 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  mat_1_1 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  mat_1_2 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  mat_1_3 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  mat_1_4 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  mat_1_5 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  mat_1_6 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  mat_1_7 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  mat_2_0 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  mat_2_1 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  mat_2_2 = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  mat_2_3 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  mat_2_4 = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  mat_2_5 = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  mat_2_6 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  mat_2_7 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  mat_3_0 = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  mat_3_1 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  mat_3_2 = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  mat_3_3 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  mat_3_4 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  mat_3_5 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  mat_3_6 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  mat_3_7 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  mat_4_0 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  mat_4_1 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  mat_4_2 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  mat_4_3 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  mat_4_4 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  mat_4_5 = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  mat_4_6 = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  mat_4_7 = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  mat_5_0 = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  mat_5_1 = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  mat_5_2 = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  mat_5_3 = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  mat_5_4 = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  mat_5_5 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  mat_5_6 = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  mat_5_7 = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  mat_6_0 = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  mat_6_1 = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  mat_6_2 = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  mat_6_3 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  mat_6_4 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  mat_6_5 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  mat_6_6 = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  mat_6_7 = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  mat_7_0 = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  mat_7_1 = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  mat_7_2 = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  mat_7_3 = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  mat_7_4 = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  mat_7_5 = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  mat_7_6 = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  mat_7_7 = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  count_0 = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  count_1 = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  count_2 = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  count_3 = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  count_4 = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  count_5 = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  count_6 = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  count_7 = _RAND_98[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ivncontrol4_3(
  input         clock,
  input         reset,
  input  [15:0] io_Stationary_matrix_0_0,
  input  [15:0] io_Stationary_matrix_0_1,
  input  [15:0] io_Stationary_matrix_0_2,
  input  [15:0] io_Stationary_matrix_0_3,
  input  [15:0] io_Stationary_matrix_0_4,
  input  [15:0] io_Stationary_matrix_0_5,
  input  [15:0] io_Stationary_matrix_0_6,
  input  [15:0] io_Stationary_matrix_0_7,
  input  [15:0] io_Stationary_matrix_1_0,
  input  [15:0] io_Stationary_matrix_1_1,
  input  [15:0] io_Stationary_matrix_1_2,
  input  [15:0] io_Stationary_matrix_1_3,
  input  [15:0] io_Stationary_matrix_1_4,
  input  [15:0] io_Stationary_matrix_1_5,
  input  [15:0] io_Stationary_matrix_1_6,
  input  [15:0] io_Stationary_matrix_1_7,
  input  [15:0] io_Stationary_matrix_2_0,
  input  [15:0] io_Stationary_matrix_2_1,
  input  [15:0] io_Stationary_matrix_2_2,
  input  [15:0] io_Stationary_matrix_2_3,
  input  [15:0] io_Stationary_matrix_2_4,
  input  [15:0] io_Stationary_matrix_2_5,
  input  [15:0] io_Stationary_matrix_2_6,
  input  [15:0] io_Stationary_matrix_2_7,
  input  [15:0] io_Stationary_matrix_3_0,
  input  [15:0] io_Stationary_matrix_3_1,
  input  [15:0] io_Stationary_matrix_3_2,
  input  [15:0] io_Stationary_matrix_3_3,
  input  [15:0] io_Stationary_matrix_3_4,
  input  [15:0] io_Stationary_matrix_3_5,
  input  [15:0] io_Stationary_matrix_3_6,
  input  [15:0] io_Stationary_matrix_3_7,
  input  [15:0] io_Stationary_matrix_4_0,
  input  [15:0] io_Stationary_matrix_4_1,
  input  [15:0] io_Stationary_matrix_4_2,
  input  [15:0] io_Stationary_matrix_4_3,
  input  [15:0] io_Stationary_matrix_4_4,
  input  [15:0] io_Stationary_matrix_4_5,
  input  [15:0] io_Stationary_matrix_4_6,
  input  [15:0] io_Stationary_matrix_4_7,
  input  [15:0] io_Stationary_matrix_5_0,
  input  [15:0] io_Stationary_matrix_5_1,
  input  [15:0] io_Stationary_matrix_5_2,
  input  [15:0] io_Stationary_matrix_5_3,
  input  [15:0] io_Stationary_matrix_5_4,
  input  [15:0] io_Stationary_matrix_5_5,
  input  [15:0] io_Stationary_matrix_5_6,
  input  [15:0] io_Stationary_matrix_5_7,
  input  [15:0] io_Stationary_matrix_6_0,
  input  [15:0] io_Stationary_matrix_6_1,
  input  [15:0] io_Stationary_matrix_6_2,
  input  [15:0] io_Stationary_matrix_6_3,
  input  [15:0] io_Stationary_matrix_6_4,
  input  [15:0] io_Stationary_matrix_6_5,
  input  [15:0] io_Stationary_matrix_6_6,
  input  [15:0] io_Stationary_matrix_6_7,
  input  [15:0] io_Stationary_matrix_7_0,
  input  [15:0] io_Stationary_matrix_7_1,
  input  [15:0] io_Stationary_matrix_7_2,
  input  [15:0] io_Stationary_matrix_7_3,
  input  [15:0] io_Stationary_matrix_7_4,
  input  [15:0] io_Stationary_matrix_7_5,
  input  [15:0] io_Stationary_matrix_7_6,
  input  [15:0] io_Stationary_matrix_7_7,
  output [4:0]  io_o_vn_0,
  output [4:0]  io_o_vn_1,
  output [4:0]  io_o_vn_2,
  output [4:0]  io_o_vn_3,
  output [4:0]  io_o_vn2_0,
  output [4:0]  io_o_vn2_1,
  output [4:0]  io_o_vn2_2,
  output [4:0]  io_o_vn2_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
`endif // RANDOMIZE_REG_INIT
  reg [4:0] i_vn_0; // @[ivncontrol4.scala 16:23]
  reg [4:0] i_vn_1; // @[ivncontrol4.scala 16:23]
  reg [4:0] i_vn_2; // @[ivncontrol4.scala 16:23]
  reg [4:0] i_vn_3; // @[ivncontrol4.scala 16:23]
  reg [4:0] i_vn2_0; // @[ivncontrol4.scala 17:24]
  reg [4:0] i_vn2_1; // @[ivncontrol4.scala 17:24]
  reg [4:0] i_vn2_2; // @[ivncontrol4.scala 17:24]
  reg [4:0] i_vn2_3; // @[ivncontrol4.scala 17:24]
  reg [31:0] rowcount_0; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_1; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_2; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_3; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_4; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_5; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_6; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_7; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_8; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_9; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_10; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_11; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_12; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_13; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_14; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_15; // @[ivncontrol4.scala 21:27]
  reg [31:0] pin; // @[ivncontrol4.scala 31:22]
  reg [31:0] i; // @[ivncontrol4.scala 35:20]
  reg [31:0] j; // @[ivncontrol4.scala 36:20]
  wire  _k_T_1 = j == 32'h7; // @[ivncontrol4.scala 38:37]
  wire  _k_T_2 = i == 32'h7 & j == 32'h7; // @[ivncontrol4.scala 38:31]
  reg [31:0] mat_0_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_0_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_0_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_0_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_0_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_0_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_0_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_0_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] count_0; // @[ivncontrol4.scala 52:20]
  reg [31:0] count_1; // @[ivncontrol4.scala 52:20]
  reg [31:0] count_2; // @[ivncontrol4.scala 52:20]
  reg [31:0] count_3; // @[ivncontrol4.scala 52:20]
  reg [31:0] count_4; // @[ivncontrol4.scala 52:20]
  reg [31:0] count_5; // @[ivncontrol4.scala 52:20]
  reg [31:0] count_6; // @[ivncontrol4.scala 52:20]
  reg [31:0] count_7; // @[ivncontrol4.scala 52:20]
  wire [15:0] _GEN_66 = 3'h0 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_0_1 : io_Stationary_matrix_0_0; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_67 = 3'h0 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_0_2 : _GEN_66; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_68 = 3'h0 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_0_3 : _GEN_67; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_69 = 3'h0 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_0_4 : _GEN_68; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_70 = 3'h0 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_0_5 : _GEN_69; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_71 = 3'h0 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_0_6 : _GEN_70; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_72 = 3'h0 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_0_7 : _GEN_71; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_73 = 3'h1 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_1_0 : _GEN_72; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_74 = 3'h1 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_1_1 : _GEN_73; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_75 = 3'h1 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_1_2 : _GEN_74; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_76 = 3'h1 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_1_3 : _GEN_75; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_77 = 3'h1 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_1_4 : _GEN_76; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_78 = 3'h1 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_1_5 : _GEN_77; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_79 = 3'h1 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_1_6 : _GEN_78; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_80 = 3'h1 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_1_7 : _GEN_79; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_81 = 3'h2 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_2_0 : _GEN_80; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_82 = 3'h2 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_2_1 : _GEN_81; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_83 = 3'h2 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_2_2 : _GEN_82; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_84 = 3'h2 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_2_3 : _GEN_83; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_85 = 3'h2 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_2_4 : _GEN_84; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_86 = 3'h2 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_2_5 : _GEN_85; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_87 = 3'h2 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_2_6 : _GEN_86; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_88 = 3'h2 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_2_7 : _GEN_87; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_89 = 3'h3 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_3_0 : _GEN_88; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_90 = 3'h3 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_3_1 : _GEN_89; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_91 = 3'h3 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_3_2 : _GEN_90; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_92 = 3'h3 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_3_3 : _GEN_91; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_93 = 3'h3 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_3_4 : _GEN_92; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_94 = 3'h3 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_3_5 : _GEN_93; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_95 = 3'h3 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_3_6 : _GEN_94; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_96 = 3'h3 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_3_7 : _GEN_95; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_97 = 3'h4 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_4_0 : _GEN_96; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_98 = 3'h4 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_4_1 : _GEN_97; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_99 = 3'h4 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_4_2 : _GEN_98; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_100 = 3'h4 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_4_3 : _GEN_99; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_101 = 3'h4 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_4_4 : _GEN_100; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_102 = 3'h4 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_4_5 : _GEN_101; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_103 = 3'h4 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_4_6 : _GEN_102; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_104 = 3'h4 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_4_7 : _GEN_103; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_105 = 3'h5 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_5_0 : _GEN_104; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_106 = 3'h5 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_5_1 : _GEN_105; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_107 = 3'h5 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_5_2 : _GEN_106; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_108 = 3'h5 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_5_3 : _GEN_107; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_109 = 3'h5 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_5_4 : _GEN_108; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_110 = 3'h5 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_5_5 : _GEN_109; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_111 = 3'h5 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_5_6 : _GEN_110; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_112 = 3'h5 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_5_7 : _GEN_111; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_113 = 3'h6 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_6_0 : _GEN_112; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_114 = 3'h6 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_6_1 : _GEN_113; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_115 = 3'h6 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_6_2 : _GEN_114; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_116 = 3'h6 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_6_3 : _GEN_115; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_117 = 3'h6 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_6_4 : _GEN_116; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_118 = 3'h6 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_6_5 : _GEN_117; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_119 = 3'h6 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_6_6 : _GEN_118; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_120 = 3'h6 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_6_7 : _GEN_119; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_121 = 3'h7 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_7_0 : _GEN_120; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_122 = 3'h7 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_7_1 : _GEN_121; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_123 = 3'h7 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_7_2 : _GEN_122; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_124 = 3'h7 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_7_3 : _GEN_123; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_125 = 3'h7 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_7_4 : _GEN_124; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_126 = 3'h7 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_7_5 : _GEN_125; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_127 = 3'h7 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_7_6 : _GEN_126; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_128 = 3'h7 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_7_7 : _GEN_127; // @[ivncontrol4.scala 57:{15,15}]
  wire [31:0] _mat_T_3_T_4 = {{16'd0}, _GEN_128}; // @[ivncontrol4.scala 57:{15,15}]
  wire  _GEN_225 = count_7 >= 32'h8; // @[ivncontrol4.scala 66:28 67:16]
  wire  valid1 = count_7 >= 32'h8; // @[ivncontrol4.scala 66:28 67:16]
  wire [31:0] _GEN_194 = 3'h1 == i[2:0] ? count_1 : count_0; // @[ivncontrol4.scala 60:{33,33}]
  wire [31:0] _GEN_195 = 3'h2 == i[2:0] ? count_2 : _GEN_194; // @[ivncontrol4.scala 60:{33,33}]
  wire [31:0] _GEN_196 = 3'h3 == i[2:0] ? count_3 : _GEN_195; // @[ivncontrol4.scala 60:{33,33}]
  wire [31:0] _GEN_197 = 3'h4 == i[2:0] ? count_4 : _GEN_196; // @[ivncontrol4.scala 60:{33,33}]
  wire [31:0] _GEN_198 = 3'h5 == i[2:0] ? count_5 : _GEN_197; // @[ivncontrol4.scala 60:{33,33}]
  wire [31:0] _GEN_199 = 3'h6 == i[2:0] ? count_6 : _GEN_198; // @[ivncontrol4.scala 60:{33,33}]
  wire [31:0] _GEN_200 = 3'h7 == i[2:0] ? count_7 : _GEN_199; // @[ivncontrol4.scala 60:{33,33}]
  wire [31:0] _count_T_2 = _GEN_200 + 32'h1; // @[ivncontrol4.scala 60:33]
  wire [31:0] _i_T_1 = i + 32'h1; // @[ivncontrol4.scala 104:16]
  wire [31:0] _j_T_1 = j + 32'h1; // @[ivncontrol4.scala 108:16]
  wire  _GEN_244 = _k_T_2; // @[ivncontrol4.scala 136:75 137:14 139:14]
  wire [31:0] _GEN_245 = rowcount_0 != 32'h0 ? 32'h0 : pin; // @[ivncontrol4.scala 145:30 146:13 31:22]
  wire  _T_27 = rowcount_0 == 32'h0; // @[ivncontrol4.scala 148:23]
  wire [31:0] _GEN_246 = rowcount_0 == 32'h0 & rowcount_1 != 32'h0 ? 32'h1 : _GEN_245; // @[ivncontrol4.scala 148:54 149:13]
  wire  _T_32 = _T_27 & rowcount_1 == 32'h0; // @[ivncontrol4.scala 151:31]
  wire [31:0] _GEN_247 = _T_27 & rowcount_1 == 32'h0 & rowcount_2 != 32'h0 ? 32'h2 : _GEN_246; // @[ivncontrol4.scala 151:77 152:13]
  wire  _T_39 = _T_32 & rowcount_2 == 32'h0; // @[ivncontrol4.scala 154:54]
  wire [31:0] _GEN_248 = _T_32 & rowcount_2 == 32'h0 & rowcount_3 != 32'h0 ? 32'h3 : _GEN_247; // @[ivncontrol4.scala 154:100 155:13]
  wire  _T_48 = _T_39 & rowcount_3 == 32'h0; // @[ivncontrol4.scala 157:77]
  wire [31:0] _GEN_249 = _T_39 & rowcount_3 == 32'h0 & rowcount_4 != 32'h0 ? 32'h4 : _GEN_248; // @[ivncontrol4.scala 157:123 158:13]
  wire  _T_59 = _T_48 & rowcount_4 == 32'h0; // @[ivncontrol4.scala 160:100]
  wire  _T_72 = _T_59 & rowcount_5 == 32'h0; // @[ivncontrol4.scala 163:123]
  wire  valid = _k_T_2; // @[ivncontrol4.scala 136:75 137:14 139:14]
  wire [32:0] _T_91 = {{1'd0}, pin}; // @[ivncontrol4.scala 174:27]
  wire [31:0] _GEN_254 = 4'h1 == _T_91[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_255 = 4'h2 == _T_91[3:0] ? rowcount_2 : _GEN_254; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_256 = 4'h3 == _T_91[3:0] ? rowcount_3 : _GEN_255; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_257 = 4'h4 == _T_91[3:0] ? rowcount_4 : _GEN_256; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_258 = 4'h5 == _T_91[3:0] ? rowcount_5 : _GEN_257; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_259 = 4'h6 == _T_91[3:0] ? rowcount_6 : _GEN_258; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_260 = 4'h7 == _T_91[3:0] ? rowcount_7 : _GEN_259; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_261 = 4'h8 == _T_91[3:0] ? rowcount_8 : _GEN_260; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_262 = 4'h9 == _T_91[3:0] ? rowcount_9 : _GEN_261; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_263 = 4'ha == _T_91[3:0] ? rowcount_10 : _GEN_262; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_264 = 4'hb == _T_91[3:0] ? rowcount_11 : _GEN_263; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_265 = 4'hc == _T_91[3:0] ? rowcount_12 : _GEN_264; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_266 = 4'hd == _T_91[3:0] ? rowcount_13 : _GEN_265; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_267 = 4'he == _T_91[3:0] ? rowcount_14 : _GEN_266; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_268 = 4'hf == _T_91[3:0] ? rowcount_15 : _GEN_267; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_381 = _GEN_268 == 32'h1 ? _T_91[31:0] : 32'h1f; // @[ivncontrol4.scala 125:17 224:50 225:21]
  wire [31:0] _GEN_382 = _GEN_268 == 32'h2 ? _T_91[31:0] : _GEN_381; // @[ivncontrol4.scala 220:51 221:21]
  wire [31:0] _GEN_383 = _GEN_268 == 32'h2 ? _T_91[31:0] : 32'h16; // @[ivncontrol4.scala 125:17 220:51 222:21]
  wire [31:0] _GEN_384 = _GEN_268 == 32'h3 ? _T_91[31:0] : _GEN_382; // @[ivncontrol4.scala 215:50 216:21]
  wire [31:0] _GEN_385 = _GEN_268 == 32'h3 ? _T_91[31:0] : _GEN_383; // @[ivncontrol4.scala 215:50 217:21]
  wire [31:0] _GEN_386 = _GEN_268 == 32'h3 ? _T_91[31:0] : 32'h7; // @[ivncontrol4.scala 125:17 215:50 218:21]
  wire [31:0] _GEN_387 = _GEN_268 == 32'h4 ? _T_91[31:0] : _GEN_384; // @[ivncontrol4.scala 207:50 208:21]
  wire [31:0] _GEN_388 = _GEN_268 == 32'h4 ? _T_91[31:0] : _GEN_385; // @[ivncontrol4.scala 207:50 209:21]
  wire [31:0] _GEN_389 = _GEN_268 == 32'h4 ? _T_91[31:0] : _GEN_386; // @[ivncontrol4.scala 207:50 210:21]
  wire [31:0] _GEN_390 = _GEN_268 == 32'h4 ? _T_91[31:0] : 32'h7; // @[ivncontrol4.scala 125:17 207:50 211:21]
  wire [31:0] _GEN_391 = _GEN_268 == 32'h5 ? _T_91[31:0] : _GEN_387; // @[ivncontrol4.scala 200:50 201:21]
  wire [31:0] _GEN_392 = _GEN_268 == 32'h5 ? _T_91[31:0] : _GEN_388; // @[ivncontrol4.scala 200:50 202:21]
  wire [31:0] _GEN_393 = _GEN_268 == 32'h5 ? _T_91[31:0] : _GEN_389; // @[ivncontrol4.scala 200:50 203:21]
  wire [31:0] _GEN_394 = _GEN_268 == 32'h5 ? _T_91[31:0] : _GEN_390; // @[ivncontrol4.scala 200:50 204:21]
  wire [31:0] _GEN_395 = _GEN_268 == 32'h5 ? _T_91[31:0] : 32'h3; // @[ivncontrol4.scala 126:18 200:50 205:22]
  wire [31:0] _GEN_396 = _GEN_268 == 32'h6 ? _T_91[31:0] : _GEN_391; // @[ivncontrol4.scala 192:52 193:21]
  wire [31:0] _GEN_397 = _GEN_268 == 32'h6 ? _T_91[31:0] : _GEN_392; // @[ivncontrol4.scala 192:52 194:21]
  wire [31:0] _GEN_398 = _GEN_268 == 32'h6 ? _T_91[31:0] : _GEN_393; // @[ivncontrol4.scala 192:52 195:21]
  wire [31:0] _GEN_399 = _GEN_268 == 32'h6 ? _T_91[31:0] : _GEN_394; // @[ivncontrol4.scala 192:52 196:21]
  wire [31:0] _GEN_400 = _GEN_268 == 32'h6 ? _T_91[31:0] : _GEN_395; // @[ivncontrol4.scala 192:52 197:22]
  wire [31:0] _GEN_401 = _GEN_268 == 32'h6 ? _T_91[31:0] : 32'h19; // @[ivncontrol4.scala 126:18 192:52 198:22]
  wire [31:0] _GEN_402 = _GEN_268 == 32'h7 ? _T_91[31:0] : _GEN_396; // @[ivncontrol4.scala 184:52 185:21]
  wire [31:0] _GEN_403 = _GEN_268 == 32'h7 ? _T_91[31:0] : _GEN_397; // @[ivncontrol4.scala 184:52 186:21]
  wire [31:0] _GEN_404 = _GEN_268 == 32'h7 ? _T_91[31:0] : _GEN_398; // @[ivncontrol4.scala 184:52 187:21]
  wire [31:0] _GEN_405 = _GEN_268 == 32'h7 ? _T_91[31:0] : _GEN_399; // @[ivncontrol4.scala 184:52 188:21]
  wire [31:0] _GEN_406 = _GEN_268 == 32'h7 ? _T_91[31:0] : _GEN_400; // @[ivncontrol4.scala 184:52 189:22]
  wire [31:0] _GEN_407 = _GEN_268 == 32'h7 ? _T_91[31:0] : _GEN_401; // @[ivncontrol4.scala 184:52 190:22]
  wire [31:0] _GEN_408 = _GEN_268 == 32'h7 ? _T_91[31:0] : 32'hb; // @[ivncontrol4.scala 126:18 184:52 191:22]
  wire [31:0] _GEN_409 = _GEN_268 >= 32'h8 ? _T_91[31:0] : _GEN_402; // @[ivncontrol4.scala 174:42 175:21]
  wire [31:0] _GEN_410 = _GEN_268 >= 32'h8 ? _T_91[31:0] : _GEN_403; // @[ivncontrol4.scala 174:42 176:21]
  wire [31:0] _GEN_411 = _GEN_268 >= 32'h8 ? _T_91[31:0] : _GEN_404; // @[ivncontrol4.scala 174:42 177:21]
  wire [31:0] _GEN_412 = _GEN_268 >= 32'h8 ? _T_91[31:0] : _GEN_405; // @[ivncontrol4.scala 174:42 178:21]
  wire [31:0] _GEN_413 = _GEN_268 >= 32'h8 ? _T_91[31:0] : _GEN_406; // @[ivncontrol4.scala 174:42 179:22]
  wire [31:0] _GEN_414 = _GEN_268 >= 32'h8 ? _T_91[31:0] : _GEN_407; // @[ivncontrol4.scala 174:42 180:22]
  wire [31:0] _GEN_415 = _GEN_268 >= 32'h8 ? _T_91[31:0] : _GEN_408; // @[ivncontrol4.scala 174:42 181:22]
  wire [31:0] _GEN_416 = _GEN_268 >= 32'h8 ? _T_91[31:0] : 32'h1f; // @[ivncontrol4.scala 126:18 174:42 182:22]
  wire [31:0] _T_127 = 32'h8 - _GEN_268; // @[ivncontrol4.scala 228:18]
  wire [31:0] _i_vn_1_T_15 = 32'h1 + pin; // @[ivncontrol4.scala 229:29]
  wire [31:0] _GEN_529 = _T_127 == 32'h1 ? _i_vn_1_T_15 : _GEN_416; // @[ivncontrol4.scala 269:54 272:22]
  wire [31:0] _GEN_530 = _T_127 == 32'h2 ? _i_vn_1_T_15 : _GEN_415; // @[ivncontrol4.scala 264:54 267:22]
  wire [31:0] _GEN_531 = _T_127 == 32'h2 ? _i_vn_1_T_15 : _GEN_529; // @[ivncontrol4.scala 264:54 268:22]
  wire [31:0] _GEN_532 = _T_127 == 32'h3 ? _i_vn_1_T_15 : _GEN_414; // @[ivncontrol4.scala 257:54 259:22]
  wire [31:0] _GEN_533 = _T_127 == 32'h3 ? _i_vn_1_T_15 : _GEN_530; // @[ivncontrol4.scala 257:54 260:22]
  wire [31:0] _GEN_534 = _T_127 == 32'h3 ? _i_vn_1_T_15 : _GEN_531; // @[ivncontrol4.scala 257:54 261:22]
  wire [31:0] _GEN_535 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_413; // @[ivncontrol4.scala 251:54 253:22]
  wire [31:0] _GEN_536 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_532; // @[ivncontrol4.scala 251:54 254:22]
  wire [31:0] _GEN_537 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_533; // @[ivncontrol4.scala 251:54 255:22]
  wire [31:0] _GEN_538 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_534; // @[ivncontrol4.scala 251:54 256:22]
  wire [31:0] _GEN_539 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_412; // @[ivncontrol4.scala 244:54 246:21]
  wire [31:0] _GEN_540 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_535; // @[ivncontrol4.scala 244:54 247:22]
  wire [31:0] _GEN_541 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_536; // @[ivncontrol4.scala 244:54 248:22]
  wire [31:0] _GEN_542 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_537; // @[ivncontrol4.scala 244:54 249:22]
  wire [31:0] _GEN_543 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_538; // @[ivncontrol4.scala 244:54 250:22]
  wire [31:0] _GEN_544 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_411; // @[ivncontrol4.scala 237:54 238:22]
  wire [31:0] _GEN_545 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_539; // @[ivncontrol4.scala 237:54 239:21]
  wire [31:0] _GEN_546 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_540; // @[ivncontrol4.scala 237:54 240:22]
  wire [31:0] _GEN_547 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_541; // @[ivncontrol4.scala 237:54 241:22]
  wire [31:0] _GEN_548 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_542; // @[ivncontrol4.scala 237:54 242:22]
  wire [31:0] _GEN_549 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_543; // @[ivncontrol4.scala 237:54 243:22]
  wire [31:0] _GEN_550 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_410; // @[ivncontrol4.scala 228:49 229:22]
  wire [31:0] _GEN_551 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_544; // @[ivncontrol4.scala 228:49 230:21]
  wire [31:0] _GEN_552 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_545; // @[ivncontrol4.scala 228:49 231:21]
  wire [31:0] _GEN_553 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_546; // @[ivncontrol4.scala 228:49 232:22]
  wire [31:0] _GEN_554 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_547; // @[ivncontrol4.scala 228:49 233:22]
  wire [31:0] _GEN_555 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_548; // @[ivncontrol4.scala 228:49 234:22]
  wire [31:0] _GEN_556 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_549; // @[ivncontrol4.scala 228:49 235:22]
  wire [31:0] _GEN_574 = 4'h1 == _i_vn_1_T_15[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_575 = 4'h2 == _i_vn_1_T_15[3:0] ? rowcount_2 : _GEN_574; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_576 = 4'h3 == _i_vn_1_T_15[3:0] ? rowcount_3 : _GEN_575; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_577 = 4'h4 == _i_vn_1_T_15[3:0] ? rowcount_4 : _GEN_576; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_578 = 4'h5 == _i_vn_1_T_15[3:0] ? rowcount_5 : _GEN_577; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_579 = 4'h6 == _i_vn_1_T_15[3:0] ? rowcount_6 : _GEN_578; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_580 = 4'h7 == _i_vn_1_T_15[3:0] ? rowcount_7 : _GEN_579; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_581 = 4'h8 == _i_vn_1_T_15[3:0] ? rowcount_8 : _GEN_580; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_582 = 4'h9 == _i_vn_1_T_15[3:0] ? rowcount_9 : _GEN_581; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_583 = 4'ha == _i_vn_1_T_15[3:0] ? rowcount_10 : _GEN_582; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_584 = 4'hb == _i_vn_1_T_15[3:0] ? rowcount_11 : _GEN_583; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_585 = 4'hc == _i_vn_1_T_15[3:0] ? rowcount_12 : _GEN_584; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_586 = 4'hd == _i_vn_1_T_15[3:0] ? rowcount_13 : _GEN_585; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_587 = 4'he == _i_vn_1_T_15[3:0] ? rowcount_14 : _GEN_586; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_588 = 4'hf == _i_vn_1_T_15[3:0] ? rowcount_15 : _GEN_587; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _T_172 = _GEN_268 + _GEN_588; // @[ivncontrol4.scala 275:41]
  wire [31:0] _T_174 = 32'h8 - _T_172; // @[ivncontrol4.scala 275:18]
  wire [31:0] _i_vn_1_T_17 = 32'h2 + pin; // @[ivncontrol4.scala 276:29]
  wire [31:0] _GEN_781 = _T_174 == 32'h1 ? _i_vn_1_T_17 : _GEN_556; // @[ivncontrol4.scala 318:78 321:22]
  wire [31:0] _GEN_782 = _T_174 == 32'h2 ? _i_vn_1_T_17 : _GEN_555; // @[ivncontrol4.scala 312:76 315:22]
  wire [31:0] _GEN_783 = _T_174 == 32'h2 ? _i_vn_1_T_17 : _GEN_781; // @[ivncontrol4.scala 312:76 316:22]
  wire [31:0] _GEN_784 = _T_174 == 32'h3 ? _i_vn_1_T_17 : _GEN_554; // @[ivncontrol4.scala 305:78 307:23]
  wire [31:0] _GEN_785 = _T_174 == 32'h3 ? _i_vn_1_T_17 : _GEN_782; // @[ivncontrol4.scala 305:78 308:22]
  wire [31:0] _GEN_786 = _T_174 == 32'h3 ? _i_vn_1_T_17 : _GEN_783; // @[ivncontrol4.scala 305:78 309:22]
  wire [31:0] _GEN_787 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_553; // @[ivncontrol4.scala 299:78 301:22]
  wire [31:0] _GEN_788 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_784; // @[ivncontrol4.scala 299:78 302:22]
  wire [31:0] _GEN_789 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_785; // @[ivncontrol4.scala 299:78 303:22]
  wire [31:0] _GEN_790 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_786; // @[ivncontrol4.scala 299:78 304:22]
  wire [31:0] _GEN_791 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_552; // @[ivncontrol4.scala 292:76 294:23]
  wire [31:0] _GEN_792 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_787; // @[ivncontrol4.scala 292:76 295:22]
  wire [31:0] _GEN_793 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_788; // @[ivncontrol4.scala 292:76 296:22]
  wire [31:0] _GEN_794 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_789; // @[ivncontrol4.scala 292:76 297:22]
  wire [31:0] _GEN_795 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_790; // @[ivncontrol4.scala 292:76 298:22]
  wire [31:0] _GEN_796 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_551; // @[ivncontrol4.scala 284:77 286:22]
  wire [31:0] _GEN_797 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_791; // @[ivncontrol4.scala 284:77 287:21]
  wire [31:0] _GEN_798 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_792; // @[ivncontrol4.scala 284:77 288:22]
  wire [31:0] _GEN_799 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_793; // @[ivncontrol4.scala 284:77 289:22]
  wire [31:0] _GEN_800 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_794; // @[ivncontrol4.scala 284:77 290:22]
  wire [31:0] _GEN_801 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_795; // @[ivncontrol4.scala 284:77 291:22]
  wire [31:0] _GEN_802 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_550; // @[ivncontrol4.scala 275:73 276:22]
  wire [31:0] _GEN_803 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_796; // @[ivncontrol4.scala 275:73 277:21]
  wire [31:0] _GEN_804 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_797; // @[ivncontrol4.scala 275:73 278:21]
  wire [31:0] _GEN_805 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_798; // @[ivncontrol4.scala 275:73 279:22]
  wire [31:0] _GEN_806 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_799; // @[ivncontrol4.scala 275:73 280:22]
  wire [31:0] _GEN_807 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_800; // @[ivncontrol4.scala 275:73 281:22]
  wire [31:0] _GEN_808 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_801; // @[ivncontrol4.scala 275:73 282:22]
  wire [31:0] _GEN_842 = 4'h1 == _i_vn_1_T_17[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_843 = 4'h2 == _i_vn_1_T_17[3:0] ? rowcount_2 : _GEN_842; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_844 = 4'h3 == _i_vn_1_T_17[3:0] ? rowcount_3 : _GEN_843; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_845 = 4'h4 == _i_vn_1_T_17[3:0] ? rowcount_4 : _GEN_844; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_846 = 4'h5 == _i_vn_1_T_17[3:0] ? rowcount_5 : _GEN_845; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_847 = 4'h6 == _i_vn_1_T_17[3:0] ? rowcount_6 : _GEN_846; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_848 = 4'h7 == _i_vn_1_T_17[3:0] ? rowcount_7 : _GEN_847; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_849 = 4'h8 == _i_vn_1_T_17[3:0] ? rowcount_8 : _GEN_848; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_850 = 4'h9 == _i_vn_1_T_17[3:0] ? rowcount_9 : _GEN_849; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_851 = 4'ha == _i_vn_1_T_17[3:0] ? rowcount_10 : _GEN_850; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_852 = 4'hb == _i_vn_1_T_17[3:0] ? rowcount_11 : _GEN_851; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_853 = 4'hc == _i_vn_1_T_17[3:0] ? rowcount_12 : _GEN_852; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_854 = 4'hd == _i_vn_1_T_17[3:0] ? rowcount_13 : _GEN_853; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_855 = 4'he == _i_vn_1_T_17[3:0] ? rowcount_14 : _GEN_854; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_856 = 4'hf == _i_vn_1_T_17[3:0] ? rowcount_15 : _GEN_855; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _T_254 = _T_172 + _GEN_856; // @[ivncontrol4.scala 326:62]
  wire [31:0] _T_256 = 32'h8 - _T_254; // @[ivncontrol4.scala 326:17]
  wire [31:0] _i_vn_1_T_19 = 32'h3 + pin; // @[ivncontrol4.scala 327:29]
  wire [31:0] _GEN_1145 = _T_256 == 32'h1 ? _i_vn_1_T_19 : _GEN_808; // @[ivncontrol4.scala 369:100 372:22]
  wire [31:0] _GEN_1146 = _T_256 == 32'h2 ? _i_vn_1_T_19 : _GEN_807; // @[ivncontrol4.scala 363:98 366:22]
  wire [31:0] _GEN_1147 = _T_256 == 32'h2 ? _i_vn_1_T_19 : _GEN_1145; // @[ivncontrol4.scala 363:98 367:22]
  wire [31:0] _GEN_1148 = _T_256 == 32'h3 ? _i_vn_1_T_19 : _GEN_806; // @[ivncontrol4.scala 356:100 358:23]
  wire [31:0] _GEN_1149 = _T_256 == 32'h3 ? _i_vn_1_T_19 : _GEN_1146; // @[ivncontrol4.scala 356:100 359:22]
  wire [31:0] _GEN_1150 = _T_256 == 32'h3 ? _i_vn_1_T_19 : _GEN_1147; // @[ivncontrol4.scala 356:100 360:22]
  wire [31:0] _GEN_1151 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_805; // @[ivncontrol4.scala 350:100 352:22]
  wire [31:0] _GEN_1152 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_1148; // @[ivncontrol4.scala 350:100 353:22]
  wire [31:0] _GEN_1153 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_1149; // @[ivncontrol4.scala 350:100 354:22]
  wire [31:0] _GEN_1154 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_1150; // @[ivncontrol4.scala 350:100 355:22]
  wire [31:0] _GEN_1155 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_804; // @[ivncontrol4.scala 343:98 345:23]
  wire [31:0] _GEN_1156 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1151; // @[ivncontrol4.scala 343:98 346:22]
  wire [31:0] _GEN_1157 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1152; // @[ivncontrol4.scala 343:98 347:22]
  wire [31:0] _GEN_1158 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1153; // @[ivncontrol4.scala 343:98 348:22]
  wire [31:0] _GEN_1159 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1154; // @[ivncontrol4.scala 343:98 349:22]
  wire [31:0] _GEN_1160 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_803; // @[ivncontrol4.scala 335:99 337:22]
  wire [31:0] _GEN_1161 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1155; // @[ivncontrol4.scala 335:99 338:21]
  wire [31:0] _GEN_1162 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1156; // @[ivncontrol4.scala 335:99 339:22]
  wire [31:0] _GEN_1163 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1157; // @[ivncontrol4.scala 335:99 340:22]
  wire [31:0] _GEN_1164 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1158; // @[ivncontrol4.scala 335:99 341:22]
  wire [31:0] _GEN_1165 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1159; // @[ivncontrol4.scala 335:99 342:22]
  wire [31:0] _GEN_1166 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_802; // @[ivncontrol4.scala 326:94 327:22]
  wire [31:0] _GEN_1167 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1160; // @[ivncontrol4.scala 326:94 328:21]
  wire [31:0] _GEN_1168 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1161; // @[ivncontrol4.scala 326:94 329:21]
  wire [31:0] _GEN_1169 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1162; // @[ivncontrol4.scala 326:94 330:22]
  wire [31:0] _GEN_1170 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1163; // @[ivncontrol4.scala 326:94 331:22]
  wire [31:0] _GEN_1171 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1164; // @[ivncontrol4.scala 326:94 332:22]
  wire [31:0] _GEN_1172 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1165; // @[ivncontrol4.scala 326:94 333:22]
  wire [31:0] _GEN_1222 = 4'h1 == _i_vn_1_T_19[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1223 = 4'h2 == _i_vn_1_T_19[3:0] ? rowcount_2 : _GEN_1222; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1224 = 4'h3 == _i_vn_1_T_19[3:0] ? rowcount_3 : _GEN_1223; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1225 = 4'h4 == _i_vn_1_T_19[3:0] ? rowcount_4 : _GEN_1224; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1226 = 4'h5 == _i_vn_1_T_19[3:0] ? rowcount_5 : _GEN_1225; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1227 = 4'h6 == _i_vn_1_T_19[3:0] ? rowcount_6 : _GEN_1226; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1228 = 4'h7 == _i_vn_1_T_19[3:0] ? rowcount_7 : _GEN_1227; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1229 = 4'h8 == _i_vn_1_T_19[3:0] ? rowcount_8 : _GEN_1228; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1230 = 4'h9 == _i_vn_1_T_19[3:0] ? rowcount_9 : _GEN_1229; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1231 = 4'ha == _i_vn_1_T_19[3:0] ? rowcount_10 : _GEN_1230; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1232 = 4'hb == _i_vn_1_T_19[3:0] ? rowcount_11 : _GEN_1231; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1233 = 4'hc == _i_vn_1_T_19[3:0] ? rowcount_12 : _GEN_1232; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1234 = 4'hd == _i_vn_1_T_19[3:0] ? rowcount_13 : _GEN_1233; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1235 = 4'he == _i_vn_1_T_19[3:0] ? rowcount_14 : _GEN_1234; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1236 = 4'hf == _i_vn_1_T_19[3:0] ? rowcount_15 : _GEN_1235; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _T_371 = _T_254 + _GEN_1236; // @[ivncontrol4.scala 376:86]
  wire [31:0] _T_373 = 32'h8 - _T_371; // @[ivncontrol4.scala 376:19]
  wire [31:0] _i_vn_1_T_21 = 32'h4 + pin; // @[ivncontrol4.scala 377:29]
  wire [31:0] _GEN_1621 = _T_373 == 32'h1 ? _i_vn_1_T_21 : _GEN_1172; // @[ivncontrol4.scala 419:122 422:22]
  wire [31:0] _GEN_1622 = _T_373 == 32'h2 ? _i_vn_1_T_21 : _GEN_1171; // @[ivncontrol4.scala 413:121 416:22]
  wire [31:0] _GEN_1623 = _T_373 == 32'h2 ? _i_vn_1_T_21 : _GEN_1621; // @[ivncontrol4.scala 413:121 417:22]
  wire [31:0] _GEN_1624 = _T_373 == 32'h3 ? _i_vn_1_T_21 : _GEN_1170; // @[ivncontrol4.scala 406:123 408:23]
  wire [31:0] _GEN_1625 = _T_373 == 32'h3 ? _i_vn_1_T_21 : _GEN_1622; // @[ivncontrol4.scala 406:123 409:22]
  wire [31:0] _GEN_1626 = _T_373 == 32'h3 ? _i_vn_1_T_21 : _GEN_1623; // @[ivncontrol4.scala 406:123 410:22]
  wire [31:0] _GEN_1627 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1169; // @[ivncontrol4.scala 400:122 402:22]
  wire [31:0] _GEN_1628 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1624; // @[ivncontrol4.scala 400:122 403:22]
  wire [31:0] _GEN_1629 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1625; // @[ivncontrol4.scala 400:122 404:22]
  wire [31:0] _GEN_1630 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1626; // @[ivncontrol4.scala 400:122 405:22]
  wire [31:0] _GEN_1631 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1168; // @[ivncontrol4.scala 393:121 395:23]
  wire [31:0] _GEN_1632 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1627; // @[ivncontrol4.scala 393:121 396:22]
  wire [31:0] _GEN_1633 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1628; // @[ivncontrol4.scala 393:121 397:22]
  wire [31:0] _GEN_1634 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1629; // @[ivncontrol4.scala 393:121 398:22]
  wire [31:0] _GEN_1635 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1630; // @[ivncontrol4.scala 393:121 399:22]
  wire [31:0] _GEN_1636 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1167; // @[ivncontrol4.scala 385:121 387:22]
  wire [31:0] _GEN_1637 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1631; // @[ivncontrol4.scala 385:121 388:21]
  wire [31:0] _GEN_1638 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1632; // @[ivncontrol4.scala 385:121 389:22]
  wire [31:0] _GEN_1639 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1633; // @[ivncontrol4.scala 385:121 390:22]
  wire [31:0] _GEN_1640 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1634; // @[ivncontrol4.scala 385:121 391:22]
  wire [31:0] _GEN_1641 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1635; // @[ivncontrol4.scala 385:121 392:22]
  wire [31:0] _GEN_1642 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1166; // @[ivncontrol4.scala 376:118 377:22]
  wire [31:0] _GEN_1643 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1636; // @[ivncontrol4.scala 376:118 378:21]
  wire [31:0] _GEN_1644 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1637; // @[ivncontrol4.scala 376:118 379:21]
  wire [31:0] _GEN_1645 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1638; // @[ivncontrol4.scala 376:118 380:22]
  wire [31:0] _GEN_1646 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1639; // @[ivncontrol4.scala 376:118 381:22]
  wire [31:0] _GEN_1647 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1640; // @[ivncontrol4.scala 376:118 382:22]
  wire [31:0] _GEN_1648 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1641; // @[ivncontrol4.scala 376:118 383:22]
  wire [31:0] _GEN_1714 = 4'h1 == _i_vn_1_T_21[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1715 = 4'h2 == _i_vn_1_T_21[3:0] ? rowcount_2 : _GEN_1714; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1716 = 4'h3 == _i_vn_1_T_21[3:0] ? rowcount_3 : _GEN_1715; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1717 = 4'h4 == _i_vn_1_T_21[3:0] ? rowcount_4 : _GEN_1716; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1718 = 4'h5 == _i_vn_1_T_21[3:0] ? rowcount_5 : _GEN_1717; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1719 = 4'h6 == _i_vn_1_T_21[3:0] ? rowcount_6 : _GEN_1718; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1720 = 4'h7 == _i_vn_1_T_21[3:0] ? rowcount_7 : _GEN_1719; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1721 = 4'h8 == _i_vn_1_T_21[3:0] ? rowcount_8 : _GEN_1720; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1722 = 4'h9 == _i_vn_1_T_21[3:0] ? rowcount_9 : _GEN_1721; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1723 = 4'ha == _i_vn_1_T_21[3:0] ? rowcount_10 : _GEN_1722; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1724 = 4'hb == _i_vn_1_T_21[3:0] ? rowcount_11 : _GEN_1723; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1725 = 4'hc == _i_vn_1_T_21[3:0] ? rowcount_12 : _GEN_1724; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1726 = 4'hd == _i_vn_1_T_21[3:0] ? rowcount_13 : _GEN_1725; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1727 = 4'he == _i_vn_1_T_21[3:0] ? rowcount_14 : _GEN_1726; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1728 = 4'hf == _i_vn_1_T_21[3:0] ? rowcount_15 : _GEN_1727; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _T_523 = _T_371 + _GEN_1728; // @[ivncontrol4.scala 426:108]
  wire [31:0] _T_525 = 32'h8 - _T_523; // @[ivncontrol4.scala 426:19]
  wire [31:0] _i_vn_1_T_23 = 32'h5 + pin; // @[ivncontrol4.scala 427:29]
  wire [31:0] _GEN_2209 = _T_525 == 32'h1 ? _i_vn_1_T_23 : _GEN_1648; // @[ivncontrol4.scala 469:144 472:22]
  wire [31:0] _GEN_2210 = _T_525 == 32'h2 ? _i_vn_1_T_23 : _GEN_1647; // @[ivncontrol4.scala 463:143 466:22]
  wire [31:0] _GEN_2211 = _T_525 == 32'h2 ? _i_vn_1_T_23 : _GEN_2209; // @[ivncontrol4.scala 463:143 467:22]
  wire [31:0] _GEN_2212 = _T_525 == 32'h3 ? _i_vn_1_T_23 : _GEN_1646; // @[ivncontrol4.scala 456:145 458:23]
  wire [31:0] _GEN_2213 = _T_525 == 32'h3 ? _i_vn_1_T_23 : _GEN_2210; // @[ivncontrol4.scala 456:145 459:22]
  wire [31:0] _GEN_2214 = _T_525 == 32'h3 ? _i_vn_1_T_23 : _GEN_2211; // @[ivncontrol4.scala 456:145 460:22]
  wire [31:0] _GEN_2215 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_1645; // @[ivncontrol4.scala 450:143 452:22]
  wire [31:0] _GEN_2216 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_2212; // @[ivncontrol4.scala 450:143 453:22]
  wire [31:0] _GEN_2217 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_2213; // @[ivncontrol4.scala 450:143 454:22]
  wire [31:0] _GEN_2218 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_2214; // @[ivncontrol4.scala 450:143 455:22]
  wire [31:0] _GEN_2219 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_1644; // @[ivncontrol4.scala 443:143 445:23]
  wire [31:0] _GEN_2220 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2215; // @[ivncontrol4.scala 443:143 446:22]
  wire [31:0] _GEN_2221 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2216; // @[ivncontrol4.scala 443:143 447:22]
  wire [31:0] _GEN_2222 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2217; // @[ivncontrol4.scala 443:143 448:22]
  wire [31:0] _GEN_2223 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2218; // @[ivncontrol4.scala 443:143 449:22]
  wire [31:0] _GEN_2224 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_1643; // @[ivncontrol4.scala 435:143 437:22]
  wire [31:0] _GEN_2225 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2219; // @[ivncontrol4.scala 435:143 438:21]
  wire [31:0] _GEN_2226 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2220; // @[ivncontrol4.scala 435:143 439:22]
  wire [31:0] _GEN_2227 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2221; // @[ivncontrol4.scala 435:143 440:22]
  wire [31:0] _GEN_2228 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2222; // @[ivncontrol4.scala 435:143 441:22]
  wire [31:0] _GEN_2229 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2223; // @[ivncontrol4.scala 435:143 442:22]
  wire [31:0] _GEN_2230 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_1642; // @[ivncontrol4.scala 426:140 427:22]
  wire [31:0] _GEN_2231 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2224; // @[ivncontrol4.scala 426:140 428:21]
  wire [31:0] _GEN_2232 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2225; // @[ivncontrol4.scala 426:140 429:21]
  wire [31:0] _GEN_2233 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2226; // @[ivncontrol4.scala 426:140 430:22]
  wire [31:0] _GEN_2234 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2227; // @[ivncontrol4.scala 426:140 431:22]
  wire [31:0] _GEN_2235 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2228; // @[ivncontrol4.scala 426:140 432:22]
  wire [31:0] _GEN_2236 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2229; // @[ivncontrol4.scala 426:140 433:22]
  wire [31:0] _GEN_2318 = 4'h1 == _i_vn_1_T_23[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2319 = 4'h2 == _i_vn_1_T_23[3:0] ? rowcount_2 : _GEN_2318; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2320 = 4'h3 == _i_vn_1_T_23[3:0] ? rowcount_3 : _GEN_2319; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2321 = 4'h4 == _i_vn_1_T_23[3:0] ? rowcount_4 : _GEN_2320; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2322 = 4'h5 == _i_vn_1_T_23[3:0] ? rowcount_5 : _GEN_2321; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2323 = 4'h6 == _i_vn_1_T_23[3:0] ? rowcount_6 : _GEN_2322; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2324 = 4'h7 == _i_vn_1_T_23[3:0] ? rowcount_7 : _GEN_2323; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2325 = 4'h8 == _i_vn_1_T_23[3:0] ? rowcount_8 : _GEN_2324; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2326 = 4'h9 == _i_vn_1_T_23[3:0] ? rowcount_9 : _GEN_2325; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2327 = 4'ha == _i_vn_1_T_23[3:0] ? rowcount_10 : _GEN_2326; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2328 = 4'hb == _i_vn_1_T_23[3:0] ? rowcount_11 : _GEN_2327; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2329 = 4'hc == _i_vn_1_T_23[3:0] ? rowcount_12 : _GEN_2328; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2330 = 4'hd == _i_vn_1_T_23[3:0] ? rowcount_13 : _GEN_2329; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2331 = 4'he == _i_vn_1_T_23[3:0] ? rowcount_14 : _GEN_2330; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2332 = 4'hf == _i_vn_1_T_23[3:0] ? rowcount_15 : _GEN_2331; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _T_710 = _T_523 + _GEN_2332; // @[ivncontrol4.scala 477:130]
  wire [31:0] _T_712 = 32'h8 - _T_710; // @[ivncontrol4.scala 477:19]
  wire [31:0] _i_vn_1_T_25 = 32'h6 + pin; // @[ivncontrol4.scala 478:29]
  wire [31:0] _GEN_2909 = _T_712 == 32'h1 ? _i_vn_1_T_25 : _GEN_2236; // @[ivncontrol4.scala 520:166 523:22]
  wire [31:0] _GEN_2910 = _T_712 == 32'h2 ? _i_vn_1_T_25 : _GEN_2235; // @[ivncontrol4.scala 514:166 517:22]
  wire [31:0] _GEN_2911 = _T_712 == 32'h2 ? _i_vn_1_T_25 : _GEN_2909; // @[ivncontrol4.scala 514:166 518:22]
  wire [31:0] _GEN_2912 = _T_712 == 32'h3 ? _i_vn_1_T_25 : _GEN_2234; // @[ivncontrol4.scala 507:168 509:23]
  wire [31:0] _GEN_2913 = _T_712 == 32'h3 ? _i_vn_1_T_25 : _GEN_2910; // @[ivncontrol4.scala 507:168 510:22]
  wire [31:0] _GEN_2914 = _T_712 == 32'h3 ? _i_vn_1_T_25 : _GEN_2911; // @[ivncontrol4.scala 507:168 511:22]
  wire [31:0] _GEN_2915 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2233; // @[ivncontrol4.scala 501:166 503:22]
  wire [31:0] _GEN_2916 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2912; // @[ivncontrol4.scala 501:166 504:22]
  wire [31:0] _GEN_2917 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2913; // @[ivncontrol4.scala 501:166 505:22]
  wire [31:0] _GEN_2918 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2914; // @[ivncontrol4.scala 501:166 506:22]
  wire [31:0] _GEN_2919 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2232; // @[ivncontrol4.scala 494:166 496:23]
  wire [31:0] _GEN_2920 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2915; // @[ivncontrol4.scala 494:166 497:22]
  wire [31:0] _GEN_2921 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2916; // @[ivncontrol4.scala 494:166 498:22]
  wire [31:0] _GEN_2922 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2917; // @[ivncontrol4.scala 494:166 499:22]
  wire [31:0] _GEN_2923 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2918; // @[ivncontrol4.scala 494:166 500:22]
  wire [31:0] _GEN_2924 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2231; // @[ivncontrol4.scala 486:166 488:22]
  wire [31:0] _GEN_2925 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2919; // @[ivncontrol4.scala 486:166 489:21]
  wire [31:0] _GEN_2926 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2920; // @[ivncontrol4.scala 486:166 490:22]
  wire [31:0] _GEN_2927 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2921; // @[ivncontrol4.scala 486:166 491:22]
  wire [31:0] _GEN_2928 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2922; // @[ivncontrol4.scala 486:166 492:22]
  wire [31:0] _GEN_2929 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2923; // @[ivncontrol4.scala 486:166 493:22]
  wire [31:0] _GEN_2930 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2230; // @[ivncontrol4.scala 477:162 478:22]
  wire [31:0] _GEN_2931 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2924; // @[ivncontrol4.scala 477:162 479:21]
  wire [31:0] _GEN_2932 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2925; // @[ivncontrol4.scala 477:162 480:21]
  wire [31:0] _GEN_2933 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2926; // @[ivncontrol4.scala 477:162 481:22]
  wire [31:0] _GEN_2934 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2927; // @[ivncontrol4.scala 477:162 482:22]
  wire [31:0] _GEN_2935 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2928; // @[ivncontrol4.scala 477:162 483:22]
  wire [31:0] _GEN_2936 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2929; // @[ivncontrol4.scala 477:162 484:22]
  wire [31:0] _GEN_3034 = 4'h1 == _i_vn_1_T_25[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3035 = 4'h2 == _i_vn_1_T_25[3:0] ? rowcount_2 : _GEN_3034; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3036 = 4'h3 == _i_vn_1_T_25[3:0] ? rowcount_3 : _GEN_3035; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3037 = 4'h4 == _i_vn_1_T_25[3:0] ? rowcount_4 : _GEN_3036; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3038 = 4'h5 == _i_vn_1_T_25[3:0] ? rowcount_5 : _GEN_3037; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3039 = 4'h6 == _i_vn_1_T_25[3:0] ? rowcount_6 : _GEN_3038; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3040 = 4'h7 == _i_vn_1_T_25[3:0] ? rowcount_7 : _GEN_3039; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3041 = 4'h8 == _i_vn_1_T_25[3:0] ? rowcount_8 : _GEN_3040; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3042 = 4'h9 == _i_vn_1_T_25[3:0] ? rowcount_9 : _GEN_3041; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3043 = 4'ha == _i_vn_1_T_25[3:0] ? rowcount_10 : _GEN_3042; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3044 = 4'hb == _i_vn_1_T_25[3:0] ? rowcount_11 : _GEN_3043; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3045 = 4'hc == _i_vn_1_T_25[3:0] ? rowcount_12 : _GEN_3044; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3046 = 4'hd == _i_vn_1_T_25[3:0] ? rowcount_13 : _GEN_3045; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3047 = 4'he == _i_vn_1_T_25[3:0] ? rowcount_14 : _GEN_3046; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3048 = 4'hf == _i_vn_1_T_25[3:0] ? rowcount_15 : _GEN_3047; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _T_932 = _T_710 + _GEN_3048; // @[ivncontrol4.scala 528:152]
  wire [31:0] _T_934 = 32'h8 - _T_932; // @[ivncontrol4.scala 528:19]
  wire [31:0] _i_vn_1_T_27 = 32'h7 + pin; // @[ivncontrol4.scala 529:29]
  wire [31:0] _GEN_3721 = _T_934 == 32'h1 ? _i_vn_1_T_27 : _GEN_2936; // @[ivncontrol4.scala 571:188 574:22]
  wire [31:0] _GEN_3722 = _T_934 == 32'h2 ? _i_vn_1_T_27 : _GEN_2935; // @[ivncontrol4.scala 565:188 568:22]
  wire [31:0] _GEN_3723 = _T_934 == 32'h2 ? _i_vn_1_T_27 : _GEN_3721; // @[ivncontrol4.scala 565:188 569:22]
  wire [31:0] _GEN_3724 = _T_934 == 32'h3 ? _i_vn_1_T_27 : _GEN_2934; // @[ivncontrol4.scala 558:190 560:23]
  wire [31:0] _GEN_3725 = _T_934 == 32'h3 ? _i_vn_1_T_27 : _GEN_3722; // @[ivncontrol4.scala 558:190 561:22]
  wire [31:0] _GEN_3726 = _T_934 == 32'h3 ? _i_vn_1_T_27 : _GEN_3723; // @[ivncontrol4.scala 558:190 562:22]
  wire [31:0] _GEN_3727 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_2933; // @[ivncontrol4.scala 552:188 554:22]
  wire [31:0] _GEN_3728 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_3724; // @[ivncontrol4.scala 552:188 555:22]
  wire [31:0] _GEN_3729 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_3725; // @[ivncontrol4.scala 552:188 556:22]
  wire [31:0] _GEN_3730 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_3726; // @[ivncontrol4.scala 552:188 557:22]
  wire [31:0] _GEN_3731 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_2932; // @[ivncontrol4.scala 545:188 547:23]
  wire [31:0] _GEN_3732 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3727; // @[ivncontrol4.scala 545:188 548:22]
  wire [31:0] _GEN_3733 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3728; // @[ivncontrol4.scala 545:188 549:22]
  wire [31:0] _GEN_3734 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3729; // @[ivncontrol4.scala 545:188 550:22]
  wire [31:0] _GEN_3735 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3730; // @[ivncontrol4.scala 545:188 551:22]
  wire [31:0] _GEN_3736 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_2931; // @[ivncontrol4.scala 537:188 539:22]
  wire [31:0] _GEN_3737 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3731; // @[ivncontrol4.scala 537:188 540:21]
  wire [31:0] _GEN_3738 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3732; // @[ivncontrol4.scala 537:188 541:22]
  wire [31:0] _GEN_3739 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3733; // @[ivncontrol4.scala 537:188 542:22]
  wire [31:0] _GEN_3740 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3734; // @[ivncontrol4.scala 537:188 543:22]
  wire [31:0] _GEN_3741 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3735; // @[ivncontrol4.scala 537:188 544:22]
  wire [31:0] _GEN_3742 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_2930; // @[ivncontrol4.scala 528:184 529:22]
  wire [31:0] _GEN_3743 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3736; // @[ivncontrol4.scala 528:184 530:21]
  wire [31:0] _GEN_3744 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3737; // @[ivncontrol4.scala 528:184 531:21]
  wire [31:0] _GEN_3745 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3738; // @[ivncontrol4.scala 528:184 532:22]
  wire [31:0] _GEN_3746 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3739; // @[ivncontrol4.scala 528:184 533:22]
  wire [31:0] _GEN_3747 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3740; // @[ivncontrol4.scala 528:184 534:22]
  wire [31:0] _GEN_3748 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3741; // @[ivncontrol4.scala 528:184 535:22]
  wire [31:0] _GEN_3749 = _GEN_244 ? _GEN_409 : 32'h1f; // @[ivncontrol4.scala 125:17 172:28]
  wire [31:0] _GEN_3750 = _GEN_244 ? _GEN_3742 : 32'h16; // @[ivncontrol4.scala 125:17 172:28]
  wire [31:0] _GEN_3751 = _GEN_244 ? _GEN_3743 : 32'h7; // @[ivncontrol4.scala 125:17 172:28]
  wire [31:0] _GEN_3752 = _GEN_244 ? _GEN_3744 : 32'h7; // @[ivncontrol4.scala 125:17 172:28]
  wire [31:0] _GEN_3753 = _GEN_244 ? _GEN_3745 : 32'h3; // @[ivncontrol4.scala 126:18 172:28]
  wire [31:0] _GEN_3754 = _GEN_244 ? _GEN_3746 : 32'h19; // @[ivncontrol4.scala 126:18 172:28]
  wire [31:0] _GEN_3755 = _GEN_244 ? _GEN_3747 : 32'hb; // @[ivncontrol4.scala 126:18 172:28]
  wire [31:0] _GEN_3756 = _GEN_244 ? _GEN_3748 : 32'h1f; // @[ivncontrol4.scala 126:18 172:28]
  wire [31:0] _GEN_4137 = reset ? 32'h0 : _GEN_3749; // @[ivncontrol4.scala 16:{23,23}]
  wire [31:0] _GEN_4138 = reset ? 32'h0 : _GEN_3750; // @[ivncontrol4.scala 16:{23,23}]
  wire [31:0] _GEN_4139 = reset ? 32'h0 : _GEN_3751; // @[ivncontrol4.scala 16:{23,23}]
  wire [31:0] _GEN_4140 = reset ? 32'h0 : _GEN_3752; // @[ivncontrol4.scala 16:{23,23}]
  wire [31:0] _GEN_4141 = reset ? 32'h0 : _GEN_3753; // @[ivncontrol4.scala 17:{24,24}]
  wire [31:0] _GEN_4142 = reset ? 32'h0 : _GEN_3754; // @[ivncontrol4.scala 17:{24,24}]
  wire [31:0] _GEN_4143 = reset ? 32'h0 : _GEN_3755; // @[ivncontrol4.scala 17:{24,24}]
  wire [31:0] _GEN_4144 = reset ? 32'h0 : _GEN_3756; // @[ivncontrol4.scala 17:{24,24}]
  assign io_o_vn_0 = i_vn_0; // @[ivncontrol4.scala 121:13]
  assign io_o_vn_1 = i_vn_1; // @[ivncontrol4.scala 121:13]
  assign io_o_vn_2 = i_vn_2; // @[ivncontrol4.scala 121:13]
  assign io_o_vn_3 = i_vn_3; // @[ivncontrol4.scala 121:13]
  assign io_o_vn2_0 = i_vn2_0; // @[ivncontrol4.scala 122:14]
  assign io_o_vn2_1 = i_vn2_1; // @[ivncontrol4.scala 122:14]
  assign io_o_vn2_2 = i_vn2_2; // @[ivncontrol4.scala 122:14]
  assign io_o_vn2_3 = i_vn2_3; // @[ivncontrol4.scala 122:14]
  always @(posedge clock) begin
    i_vn_0 <= _GEN_4137[4:0]; // @[ivncontrol4.scala 16:{23,23}]
    i_vn_1 <= _GEN_4138[4:0]; // @[ivncontrol4.scala 16:{23,23}]
    i_vn_2 <= _GEN_4139[4:0]; // @[ivncontrol4.scala 16:{23,23}]
    i_vn_3 <= _GEN_4140[4:0]; // @[ivncontrol4.scala 16:{23,23}]
    i_vn2_0 <= _GEN_4141[4:0]; // @[ivncontrol4.scala 17:{24,24}]
    i_vn2_1 <= _GEN_4142[4:0]; // @[ivncontrol4.scala 17:{24,24}]
    i_vn2_2 <= _GEN_4143[4:0]; // @[ivncontrol4.scala 17:{24,24}]
    i_vn2_3 <= _GEN_4144[4:0]; // @[ivncontrol4.scala 17:{24,24}]
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_0 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_0 <= count_0; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_1 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_1 <= count_1; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_2 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_2 <= count_2; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_3 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_3 <= count_3; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_4 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_4 <= count_4; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_5 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_5 <= count_5; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_6 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_6 <= count_6; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_7 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_7 <= count_7; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_8 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_8 <= 32'h0; // @[ivncontrol4.scala 81:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_9 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_9 <= 32'h0; // @[ivncontrol4.scala 81:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_10 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_10 <= 32'h0; // @[ivncontrol4.scala 81:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_11 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_11 <= 32'h0; // @[ivncontrol4.scala 81:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_12 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_12 <= 32'h0; // @[ivncontrol4.scala 81:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_13 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_13 <= 32'h0; // @[ivncontrol4.scala 81:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_14 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_14 <= 32'h0; // @[ivncontrol4.scala 81:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_15 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end
    if (reset) begin // @[ivncontrol4.scala 31:22]
      pin <= 32'h0; // @[ivncontrol4.scala 31:22]
    end else if (_T_72 & rowcount_6 == 32'h0 & rowcount_7 != 32'h0) begin // @[ivncontrol4.scala 166:192]
      pin <= 32'h7; // @[ivncontrol4.scala 167:13]
    end else if (_T_59 & rowcount_5 == 32'h0 & rowcount_6 != 32'h0) begin // @[ivncontrol4.scala 163:169]
      pin <= 32'h6; // @[ivncontrol4.scala 164:13]
    end else if (_T_48 & rowcount_4 == 32'h0 & rowcount_5 != 32'h0) begin // @[ivncontrol4.scala 160:146]
      pin <= 32'h5; // @[ivncontrol4.scala 161:13]
    end else begin
      pin <= _GEN_249;
    end
    if (reset) begin // @[ivncontrol4.scala 35:20]
      i <= 32'h0; // @[ivncontrol4.scala 35:20]
    end else if (i < 32'h7 & _k_T_1) begin // @[ivncontrol4.scala 103:74]
      i <= _i_T_1; // @[ivncontrol4.scala 104:11]
    end
    if (reset) begin // @[ivncontrol4.scala 36:20]
      j <= 32'h0; // @[ivncontrol4.scala 36:20]
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 107:71]
      j <= _j_T_1; // @[ivncontrol4.scala 108:11]
    end else if (!(_k_T_2)) begin // @[ivncontrol4.scala 110:81]
      j <= 32'h0; // @[ivncontrol4.scala 114:11]
    end
    if (3'h0 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h0 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h0 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h0 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h0 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h0 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h0 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h0 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h0 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_0 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h1 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_1 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h2 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_2 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h3 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_3 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h4 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_4 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h5 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_5 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h6 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_6 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h7 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_7 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  i_vn_0 = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  i_vn_1 = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  i_vn_2 = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  i_vn_3 = _RAND_3[4:0];
  _RAND_4 = {1{`RANDOM}};
  i_vn2_0 = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  i_vn2_1 = _RAND_5[4:0];
  _RAND_6 = {1{`RANDOM}};
  i_vn2_2 = _RAND_6[4:0];
  _RAND_7 = {1{`RANDOM}};
  i_vn2_3 = _RAND_7[4:0];
  _RAND_8 = {1{`RANDOM}};
  rowcount_0 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  rowcount_1 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  rowcount_2 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  rowcount_3 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  rowcount_4 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  rowcount_5 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  rowcount_6 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  rowcount_7 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  rowcount_8 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  rowcount_9 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  rowcount_10 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  rowcount_11 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  rowcount_12 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  rowcount_13 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  rowcount_14 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  rowcount_15 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  pin = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  i = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  j = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  mat_0_0 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  mat_0_1 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  mat_0_2 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  mat_0_3 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  mat_0_4 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  mat_0_5 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  mat_0_6 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  mat_0_7 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  mat_1_0 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  mat_1_1 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  mat_1_2 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  mat_1_3 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  mat_1_4 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  mat_1_5 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  mat_1_6 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  mat_1_7 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  mat_2_0 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  mat_2_1 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  mat_2_2 = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  mat_2_3 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  mat_2_4 = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  mat_2_5 = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  mat_2_6 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  mat_2_7 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  mat_3_0 = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  mat_3_1 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  mat_3_2 = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  mat_3_3 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  mat_3_4 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  mat_3_5 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  mat_3_6 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  mat_3_7 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  mat_4_0 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  mat_4_1 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  mat_4_2 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  mat_4_3 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  mat_4_4 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  mat_4_5 = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  mat_4_6 = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  mat_4_7 = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  mat_5_0 = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  mat_5_1 = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  mat_5_2 = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  mat_5_3 = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  mat_5_4 = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  mat_5_5 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  mat_5_6 = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  mat_5_7 = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  mat_6_0 = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  mat_6_1 = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  mat_6_2 = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  mat_6_3 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  mat_6_4 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  mat_6_5 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  mat_6_6 = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  mat_6_7 = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  mat_7_0 = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  mat_7_1 = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  mat_7_2 = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  mat_7_3 = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  mat_7_4 = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  mat_7_5 = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  mat_7_6 = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  mat_7_7 = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  count_0 = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  count_1 = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  count_2 = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  count_3 = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  count_4 = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  count_5 = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  count_6 = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  count_7 = _RAND_98[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ivncontrol4_4(
  input         clock,
  input         reset,
  input  [15:0] io_Stationary_matrix_0_0,
  input  [15:0] io_Stationary_matrix_0_1,
  input  [15:0] io_Stationary_matrix_0_2,
  input  [15:0] io_Stationary_matrix_0_3,
  input  [15:0] io_Stationary_matrix_0_4,
  input  [15:0] io_Stationary_matrix_0_5,
  input  [15:0] io_Stationary_matrix_0_6,
  input  [15:0] io_Stationary_matrix_0_7,
  input  [15:0] io_Stationary_matrix_1_0,
  input  [15:0] io_Stationary_matrix_1_1,
  input  [15:0] io_Stationary_matrix_1_2,
  input  [15:0] io_Stationary_matrix_1_3,
  input  [15:0] io_Stationary_matrix_1_4,
  input  [15:0] io_Stationary_matrix_1_5,
  input  [15:0] io_Stationary_matrix_1_6,
  input  [15:0] io_Stationary_matrix_1_7,
  input  [15:0] io_Stationary_matrix_2_0,
  input  [15:0] io_Stationary_matrix_2_1,
  input  [15:0] io_Stationary_matrix_2_2,
  input  [15:0] io_Stationary_matrix_2_3,
  input  [15:0] io_Stationary_matrix_2_4,
  input  [15:0] io_Stationary_matrix_2_5,
  input  [15:0] io_Stationary_matrix_2_6,
  input  [15:0] io_Stationary_matrix_2_7,
  input  [15:0] io_Stationary_matrix_3_0,
  input  [15:0] io_Stationary_matrix_3_1,
  input  [15:0] io_Stationary_matrix_3_2,
  input  [15:0] io_Stationary_matrix_3_3,
  input  [15:0] io_Stationary_matrix_3_4,
  input  [15:0] io_Stationary_matrix_3_5,
  input  [15:0] io_Stationary_matrix_3_6,
  input  [15:0] io_Stationary_matrix_3_7,
  input  [15:0] io_Stationary_matrix_4_0,
  input  [15:0] io_Stationary_matrix_4_1,
  input  [15:0] io_Stationary_matrix_4_2,
  input  [15:0] io_Stationary_matrix_4_3,
  input  [15:0] io_Stationary_matrix_4_4,
  input  [15:0] io_Stationary_matrix_4_5,
  input  [15:0] io_Stationary_matrix_4_6,
  input  [15:0] io_Stationary_matrix_4_7,
  input  [15:0] io_Stationary_matrix_5_0,
  input  [15:0] io_Stationary_matrix_5_1,
  input  [15:0] io_Stationary_matrix_5_2,
  input  [15:0] io_Stationary_matrix_5_3,
  input  [15:0] io_Stationary_matrix_5_4,
  input  [15:0] io_Stationary_matrix_5_5,
  input  [15:0] io_Stationary_matrix_5_6,
  input  [15:0] io_Stationary_matrix_5_7,
  input  [15:0] io_Stationary_matrix_6_0,
  input  [15:0] io_Stationary_matrix_6_1,
  input  [15:0] io_Stationary_matrix_6_2,
  input  [15:0] io_Stationary_matrix_6_3,
  input  [15:0] io_Stationary_matrix_6_4,
  input  [15:0] io_Stationary_matrix_6_5,
  input  [15:0] io_Stationary_matrix_6_6,
  input  [15:0] io_Stationary_matrix_6_7,
  input  [15:0] io_Stationary_matrix_7_0,
  input  [15:0] io_Stationary_matrix_7_1,
  input  [15:0] io_Stationary_matrix_7_2,
  input  [15:0] io_Stationary_matrix_7_3,
  input  [15:0] io_Stationary_matrix_7_4,
  input  [15:0] io_Stationary_matrix_7_5,
  input  [15:0] io_Stationary_matrix_7_6,
  input  [15:0] io_Stationary_matrix_7_7,
  output [4:0]  io_o_vn_0,
  output [4:0]  io_o_vn_1,
  output [4:0]  io_o_vn_2,
  output [4:0]  io_o_vn_3,
  output [4:0]  io_o_vn2_0,
  output [4:0]  io_o_vn2_1,
  output [4:0]  io_o_vn2_2,
  output [4:0]  io_o_vn2_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
`endif // RANDOMIZE_REG_INIT
  reg [4:0] i_vn_0; // @[ivncontrol4.scala 16:23]
  reg [4:0] i_vn_1; // @[ivncontrol4.scala 16:23]
  reg [4:0] i_vn_2; // @[ivncontrol4.scala 16:23]
  reg [4:0] i_vn_3; // @[ivncontrol4.scala 16:23]
  reg [4:0] i_vn2_0; // @[ivncontrol4.scala 17:24]
  reg [4:0] i_vn2_1; // @[ivncontrol4.scala 17:24]
  reg [4:0] i_vn2_2; // @[ivncontrol4.scala 17:24]
  reg [4:0] i_vn2_3; // @[ivncontrol4.scala 17:24]
  reg [31:0] rowcount_0; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_1; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_2; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_3; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_4; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_5; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_6; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_7; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_8; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_9; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_10; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_11; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_12; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_13; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_14; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_15; // @[ivncontrol4.scala 21:27]
  reg [31:0] pin; // @[ivncontrol4.scala 31:22]
  reg [31:0] i; // @[ivncontrol4.scala 35:20]
  reg [31:0] j; // @[ivncontrol4.scala 36:20]
  wire  _k_T_1 = j == 32'h7; // @[ivncontrol4.scala 38:37]
  wire  _k_T_2 = i == 32'h7 & j == 32'h7; // @[ivncontrol4.scala 38:31]
  reg [31:0] mat_0_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_0_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_0_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_0_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_0_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_0_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_0_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_0_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] count_0; // @[ivncontrol4.scala 52:20]
  reg [31:0] count_1; // @[ivncontrol4.scala 52:20]
  reg [31:0] count_2; // @[ivncontrol4.scala 52:20]
  reg [31:0] count_3; // @[ivncontrol4.scala 52:20]
  reg [31:0] count_4; // @[ivncontrol4.scala 52:20]
  reg [31:0] count_5; // @[ivncontrol4.scala 52:20]
  reg [31:0] count_6; // @[ivncontrol4.scala 52:20]
  reg [31:0] count_7; // @[ivncontrol4.scala 52:20]
  wire [15:0] _GEN_66 = 3'h0 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_0_1 : io_Stationary_matrix_0_0; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_67 = 3'h0 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_0_2 : _GEN_66; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_68 = 3'h0 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_0_3 : _GEN_67; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_69 = 3'h0 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_0_4 : _GEN_68; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_70 = 3'h0 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_0_5 : _GEN_69; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_71 = 3'h0 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_0_6 : _GEN_70; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_72 = 3'h0 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_0_7 : _GEN_71; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_73 = 3'h1 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_1_0 : _GEN_72; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_74 = 3'h1 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_1_1 : _GEN_73; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_75 = 3'h1 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_1_2 : _GEN_74; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_76 = 3'h1 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_1_3 : _GEN_75; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_77 = 3'h1 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_1_4 : _GEN_76; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_78 = 3'h1 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_1_5 : _GEN_77; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_79 = 3'h1 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_1_6 : _GEN_78; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_80 = 3'h1 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_1_7 : _GEN_79; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_81 = 3'h2 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_2_0 : _GEN_80; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_82 = 3'h2 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_2_1 : _GEN_81; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_83 = 3'h2 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_2_2 : _GEN_82; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_84 = 3'h2 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_2_3 : _GEN_83; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_85 = 3'h2 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_2_4 : _GEN_84; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_86 = 3'h2 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_2_5 : _GEN_85; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_87 = 3'h2 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_2_6 : _GEN_86; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_88 = 3'h2 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_2_7 : _GEN_87; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_89 = 3'h3 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_3_0 : _GEN_88; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_90 = 3'h3 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_3_1 : _GEN_89; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_91 = 3'h3 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_3_2 : _GEN_90; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_92 = 3'h3 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_3_3 : _GEN_91; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_93 = 3'h3 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_3_4 : _GEN_92; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_94 = 3'h3 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_3_5 : _GEN_93; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_95 = 3'h3 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_3_6 : _GEN_94; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_96 = 3'h3 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_3_7 : _GEN_95; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_97 = 3'h4 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_4_0 : _GEN_96; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_98 = 3'h4 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_4_1 : _GEN_97; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_99 = 3'h4 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_4_2 : _GEN_98; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_100 = 3'h4 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_4_3 : _GEN_99; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_101 = 3'h4 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_4_4 : _GEN_100; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_102 = 3'h4 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_4_5 : _GEN_101; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_103 = 3'h4 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_4_6 : _GEN_102; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_104 = 3'h4 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_4_7 : _GEN_103; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_105 = 3'h5 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_5_0 : _GEN_104; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_106 = 3'h5 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_5_1 : _GEN_105; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_107 = 3'h5 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_5_2 : _GEN_106; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_108 = 3'h5 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_5_3 : _GEN_107; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_109 = 3'h5 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_5_4 : _GEN_108; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_110 = 3'h5 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_5_5 : _GEN_109; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_111 = 3'h5 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_5_6 : _GEN_110; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_112 = 3'h5 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_5_7 : _GEN_111; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_113 = 3'h6 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_6_0 : _GEN_112; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_114 = 3'h6 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_6_1 : _GEN_113; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_115 = 3'h6 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_6_2 : _GEN_114; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_116 = 3'h6 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_6_3 : _GEN_115; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_117 = 3'h6 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_6_4 : _GEN_116; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_118 = 3'h6 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_6_5 : _GEN_117; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_119 = 3'h6 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_6_6 : _GEN_118; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_120 = 3'h6 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_6_7 : _GEN_119; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_121 = 3'h7 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_7_0 : _GEN_120; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_122 = 3'h7 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_7_1 : _GEN_121; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_123 = 3'h7 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_7_2 : _GEN_122; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_124 = 3'h7 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_7_3 : _GEN_123; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_125 = 3'h7 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_7_4 : _GEN_124; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_126 = 3'h7 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_7_5 : _GEN_125; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_127 = 3'h7 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_7_6 : _GEN_126; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_128 = 3'h7 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_7_7 : _GEN_127; // @[ivncontrol4.scala 57:{15,15}]
  wire [31:0] _mat_T_3_T_4 = {{16'd0}, _GEN_128}; // @[ivncontrol4.scala 57:{15,15}]
  wire  _GEN_225 = count_7 >= 32'h8; // @[ivncontrol4.scala 66:28 67:16]
  wire  valid1 = count_7 >= 32'h8; // @[ivncontrol4.scala 66:28 67:16]
  wire [31:0] _GEN_194 = 3'h1 == i[2:0] ? count_1 : count_0; // @[ivncontrol4.scala 60:{33,33}]
  wire [31:0] _GEN_195 = 3'h2 == i[2:0] ? count_2 : _GEN_194; // @[ivncontrol4.scala 60:{33,33}]
  wire [31:0] _GEN_196 = 3'h3 == i[2:0] ? count_3 : _GEN_195; // @[ivncontrol4.scala 60:{33,33}]
  wire [31:0] _GEN_197 = 3'h4 == i[2:0] ? count_4 : _GEN_196; // @[ivncontrol4.scala 60:{33,33}]
  wire [31:0] _GEN_198 = 3'h5 == i[2:0] ? count_5 : _GEN_197; // @[ivncontrol4.scala 60:{33,33}]
  wire [31:0] _GEN_199 = 3'h6 == i[2:0] ? count_6 : _GEN_198; // @[ivncontrol4.scala 60:{33,33}]
  wire [31:0] _GEN_200 = 3'h7 == i[2:0] ? count_7 : _GEN_199; // @[ivncontrol4.scala 60:{33,33}]
  wire [31:0] _count_T_2 = _GEN_200 + 32'h1; // @[ivncontrol4.scala 60:33]
  wire [31:0] _i_T_1 = i + 32'h1; // @[ivncontrol4.scala 104:16]
  wire [31:0] _j_T_1 = j + 32'h1; // @[ivncontrol4.scala 108:16]
  wire  _GEN_244 = _k_T_2; // @[ivncontrol4.scala 136:75 137:14 139:14]
  wire [31:0] _GEN_245 = rowcount_0 != 32'h0 ? 32'h0 : pin; // @[ivncontrol4.scala 145:30 146:13 31:22]
  wire  _T_27 = rowcount_0 == 32'h0; // @[ivncontrol4.scala 148:23]
  wire [31:0] _GEN_246 = rowcount_0 == 32'h0 & rowcount_1 != 32'h0 ? 32'h1 : _GEN_245; // @[ivncontrol4.scala 148:54 149:13]
  wire  _T_32 = _T_27 & rowcount_1 == 32'h0; // @[ivncontrol4.scala 151:31]
  wire [31:0] _GEN_247 = _T_27 & rowcount_1 == 32'h0 & rowcount_2 != 32'h0 ? 32'h2 : _GEN_246; // @[ivncontrol4.scala 151:77 152:13]
  wire  _T_39 = _T_32 & rowcount_2 == 32'h0; // @[ivncontrol4.scala 154:54]
  wire [31:0] _GEN_248 = _T_32 & rowcount_2 == 32'h0 & rowcount_3 != 32'h0 ? 32'h3 : _GEN_247; // @[ivncontrol4.scala 154:100 155:13]
  wire  _T_48 = _T_39 & rowcount_3 == 32'h0; // @[ivncontrol4.scala 157:77]
  wire [31:0] _GEN_249 = _T_39 & rowcount_3 == 32'h0 & rowcount_4 != 32'h0 ? 32'h4 : _GEN_248; // @[ivncontrol4.scala 157:123 158:13]
  wire  _T_59 = _T_48 & rowcount_4 == 32'h0; // @[ivncontrol4.scala 160:100]
  wire  _T_72 = _T_59 & rowcount_5 == 32'h0; // @[ivncontrol4.scala 163:123]
  wire  valid = _k_T_2; // @[ivncontrol4.scala 136:75 137:14 139:14]
  wire [32:0] _T_91 = {{1'd0}, pin}; // @[ivncontrol4.scala 174:27]
  wire [31:0] _GEN_254 = 4'h1 == _T_91[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_255 = 4'h2 == _T_91[3:0] ? rowcount_2 : _GEN_254; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_256 = 4'h3 == _T_91[3:0] ? rowcount_3 : _GEN_255; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_257 = 4'h4 == _T_91[3:0] ? rowcount_4 : _GEN_256; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_258 = 4'h5 == _T_91[3:0] ? rowcount_5 : _GEN_257; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_259 = 4'h6 == _T_91[3:0] ? rowcount_6 : _GEN_258; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_260 = 4'h7 == _T_91[3:0] ? rowcount_7 : _GEN_259; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_261 = 4'h8 == _T_91[3:0] ? rowcount_8 : _GEN_260; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_262 = 4'h9 == _T_91[3:0] ? rowcount_9 : _GEN_261; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_263 = 4'ha == _T_91[3:0] ? rowcount_10 : _GEN_262; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_264 = 4'hb == _T_91[3:0] ? rowcount_11 : _GEN_263; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_265 = 4'hc == _T_91[3:0] ? rowcount_12 : _GEN_264; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_266 = 4'hd == _T_91[3:0] ? rowcount_13 : _GEN_265; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_267 = 4'he == _T_91[3:0] ? rowcount_14 : _GEN_266; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_268 = 4'hf == _T_91[3:0] ? rowcount_15 : _GEN_267; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_381 = _GEN_268 == 32'h1 ? _T_91[31:0] : 32'h19; // @[ivncontrol4.scala 125:17 224:50 225:21]
  wire [31:0] _GEN_382 = _GEN_268 == 32'h2 ? _T_91[31:0] : _GEN_381; // @[ivncontrol4.scala 220:51 221:21]
  wire [31:0] _GEN_383 = _GEN_268 == 32'h2 ? _T_91[31:0] : 32'ha; // @[ivncontrol4.scala 125:17 220:51 222:21]
  wire [31:0] _GEN_384 = _GEN_268 == 32'h3 ? _T_91[31:0] : _GEN_382; // @[ivncontrol4.scala 215:50 216:21]
  wire [31:0] _GEN_385 = _GEN_268 == 32'h3 ? _T_91[31:0] : _GEN_383; // @[ivncontrol4.scala 215:50 217:21]
  wire [31:0] _GEN_386 = _GEN_268 == 32'h3 ? _T_91[31:0] : 32'he; // @[ivncontrol4.scala 125:17 215:50 218:21]
  wire [31:0] _GEN_387 = _GEN_268 == 32'h4 ? _T_91[31:0] : _GEN_384; // @[ivncontrol4.scala 207:50 208:21]
  wire [31:0] _GEN_388 = _GEN_268 == 32'h4 ? _T_91[31:0] : _GEN_385; // @[ivncontrol4.scala 207:50 209:21]
  wire [31:0] _GEN_389 = _GEN_268 == 32'h4 ? _T_91[31:0] : _GEN_386; // @[ivncontrol4.scala 207:50 210:21]
  wire [31:0] _GEN_390 = _GEN_268 == 32'h4 ? _T_91[31:0] : 32'h4; // @[ivncontrol4.scala 125:17 207:50 211:21]
  wire [31:0] _GEN_391 = _GEN_268 == 32'h5 ? _T_91[31:0] : _GEN_387; // @[ivncontrol4.scala 200:50 201:21]
  wire [31:0] _GEN_392 = _GEN_268 == 32'h5 ? _T_91[31:0] : _GEN_388; // @[ivncontrol4.scala 200:50 202:21]
  wire [31:0] _GEN_393 = _GEN_268 == 32'h5 ? _T_91[31:0] : _GEN_389; // @[ivncontrol4.scala 200:50 203:21]
  wire [31:0] _GEN_394 = _GEN_268 == 32'h5 ? _T_91[31:0] : _GEN_390; // @[ivncontrol4.scala 200:50 204:21]
  wire [31:0] _GEN_395 = _GEN_268 == 32'h5 ? _T_91[31:0] : 32'h10; // @[ivncontrol4.scala 126:18 200:50 205:22]
  wire [31:0] _GEN_396 = _GEN_268 == 32'h6 ? _T_91[31:0] : _GEN_391; // @[ivncontrol4.scala 192:52 193:21]
  wire [31:0] _GEN_397 = _GEN_268 == 32'h6 ? _T_91[31:0] : _GEN_392; // @[ivncontrol4.scala 192:52 194:21]
  wire [31:0] _GEN_398 = _GEN_268 == 32'h6 ? _T_91[31:0] : _GEN_393; // @[ivncontrol4.scala 192:52 195:21]
  wire [31:0] _GEN_399 = _GEN_268 == 32'h6 ? _T_91[31:0] : _GEN_394; // @[ivncontrol4.scala 192:52 196:21]
  wire [31:0] _GEN_400 = _GEN_268 == 32'h6 ? _T_91[31:0] : _GEN_395; // @[ivncontrol4.scala 192:52 197:22]
  wire [31:0] _GEN_401 = _GEN_268 == 32'h6 ? _T_91[31:0] : 32'he; // @[ivncontrol4.scala 126:18 192:52 198:22]
  wire [31:0] _GEN_402 = _GEN_268 == 32'h7 ? _T_91[31:0] : _GEN_396; // @[ivncontrol4.scala 184:52 185:21]
  wire [31:0] _GEN_403 = _GEN_268 == 32'h7 ? _T_91[31:0] : _GEN_397; // @[ivncontrol4.scala 184:52 186:21]
  wire [31:0] _GEN_404 = _GEN_268 == 32'h7 ? _T_91[31:0] : _GEN_398; // @[ivncontrol4.scala 184:52 187:21]
  wire [31:0] _GEN_405 = _GEN_268 == 32'h7 ? _T_91[31:0] : _GEN_399; // @[ivncontrol4.scala 184:52 188:21]
  wire [31:0] _GEN_406 = _GEN_268 == 32'h7 ? _T_91[31:0] : _GEN_400; // @[ivncontrol4.scala 184:52 189:22]
  wire [31:0] _GEN_407 = _GEN_268 == 32'h7 ? _T_91[31:0] : _GEN_401; // @[ivncontrol4.scala 184:52 190:22]
  wire [31:0] _GEN_408 = _GEN_268 == 32'h7 ? _T_91[31:0] : 32'ha; // @[ivncontrol4.scala 126:18 184:52 191:22]
  wire [31:0] _GEN_409 = _GEN_268 >= 32'h8 ? _T_91[31:0] : _GEN_402; // @[ivncontrol4.scala 174:42 175:21]
  wire [31:0] _GEN_410 = _GEN_268 >= 32'h8 ? _T_91[31:0] : _GEN_403; // @[ivncontrol4.scala 174:42 176:21]
  wire [31:0] _GEN_411 = _GEN_268 >= 32'h8 ? _T_91[31:0] : _GEN_404; // @[ivncontrol4.scala 174:42 177:21]
  wire [31:0] _GEN_412 = _GEN_268 >= 32'h8 ? _T_91[31:0] : _GEN_405; // @[ivncontrol4.scala 174:42 178:21]
  wire [31:0] _GEN_413 = _GEN_268 >= 32'h8 ? _T_91[31:0] : _GEN_406; // @[ivncontrol4.scala 174:42 179:22]
  wire [31:0] _GEN_414 = _GEN_268 >= 32'h8 ? _T_91[31:0] : _GEN_407; // @[ivncontrol4.scala 174:42 180:22]
  wire [31:0] _GEN_415 = _GEN_268 >= 32'h8 ? _T_91[31:0] : _GEN_408; // @[ivncontrol4.scala 174:42 181:22]
  wire [31:0] _GEN_416 = _GEN_268 >= 32'h8 ? _T_91[31:0] : 32'h1; // @[ivncontrol4.scala 126:18 174:42 182:22]
  wire [31:0] _T_127 = 32'h8 - _GEN_268; // @[ivncontrol4.scala 228:18]
  wire [31:0] _i_vn_1_T_15 = 32'h1 + pin; // @[ivncontrol4.scala 229:29]
  wire [31:0] _GEN_529 = _T_127 == 32'h1 ? _i_vn_1_T_15 : _GEN_416; // @[ivncontrol4.scala 269:54 272:22]
  wire [31:0] _GEN_530 = _T_127 == 32'h2 ? _i_vn_1_T_15 : _GEN_415; // @[ivncontrol4.scala 264:54 267:22]
  wire [31:0] _GEN_531 = _T_127 == 32'h2 ? _i_vn_1_T_15 : _GEN_529; // @[ivncontrol4.scala 264:54 268:22]
  wire [31:0] _GEN_532 = _T_127 == 32'h3 ? _i_vn_1_T_15 : _GEN_414; // @[ivncontrol4.scala 257:54 259:22]
  wire [31:0] _GEN_533 = _T_127 == 32'h3 ? _i_vn_1_T_15 : _GEN_530; // @[ivncontrol4.scala 257:54 260:22]
  wire [31:0] _GEN_534 = _T_127 == 32'h3 ? _i_vn_1_T_15 : _GEN_531; // @[ivncontrol4.scala 257:54 261:22]
  wire [31:0] _GEN_535 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_413; // @[ivncontrol4.scala 251:54 253:22]
  wire [31:0] _GEN_536 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_532; // @[ivncontrol4.scala 251:54 254:22]
  wire [31:0] _GEN_537 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_533; // @[ivncontrol4.scala 251:54 255:22]
  wire [31:0] _GEN_538 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_534; // @[ivncontrol4.scala 251:54 256:22]
  wire [31:0] _GEN_539 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_412; // @[ivncontrol4.scala 244:54 246:21]
  wire [31:0] _GEN_540 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_535; // @[ivncontrol4.scala 244:54 247:22]
  wire [31:0] _GEN_541 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_536; // @[ivncontrol4.scala 244:54 248:22]
  wire [31:0] _GEN_542 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_537; // @[ivncontrol4.scala 244:54 249:22]
  wire [31:0] _GEN_543 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_538; // @[ivncontrol4.scala 244:54 250:22]
  wire [31:0] _GEN_544 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_411; // @[ivncontrol4.scala 237:54 238:22]
  wire [31:0] _GEN_545 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_539; // @[ivncontrol4.scala 237:54 239:21]
  wire [31:0] _GEN_546 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_540; // @[ivncontrol4.scala 237:54 240:22]
  wire [31:0] _GEN_547 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_541; // @[ivncontrol4.scala 237:54 241:22]
  wire [31:0] _GEN_548 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_542; // @[ivncontrol4.scala 237:54 242:22]
  wire [31:0] _GEN_549 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_543; // @[ivncontrol4.scala 237:54 243:22]
  wire [31:0] _GEN_550 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_410; // @[ivncontrol4.scala 228:49 229:22]
  wire [31:0] _GEN_551 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_544; // @[ivncontrol4.scala 228:49 230:21]
  wire [31:0] _GEN_552 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_545; // @[ivncontrol4.scala 228:49 231:21]
  wire [31:0] _GEN_553 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_546; // @[ivncontrol4.scala 228:49 232:22]
  wire [31:0] _GEN_554 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_547; // @[ivncontrol4.scala 228:49 233:22]
  wire [31:0] _GEN_555 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_548; // @[ivncontrol4.scala 228:49 234:22]
  wire [31:0] _GEN_556 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_549; // @[ivncontrol4.scala 228:49 235:22]
  wire [31:0] _GEN_574 = 4'h1 == _i_vn_1_T_15[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_575 = 4'h2 == _i_vn_1_T_15[3:0] ? rowcount_2 : _GEN_574; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_576 = 4'h3 == _i_vn_1_T_15[3:0] ? rowcount_3 : _GEN_575; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_577 = 4'h4 == _i_vn_1_T_15[3:0] ? rowcount_4 : _GEN_576; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_578 = 4'h5 == _i_vn_1_T_15[3:0] ? rowcount_5 : _GEN_577; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_579 = 4'h6 == _i_vn_1_T_15[3:0] ? rowcount_6 : _GEN_578; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_580 = 4'h7 == _i_vn_1_T_15[3:0] ? rowcount_7 : _GEN_579; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_581 = 4'h8 == _i_vn_1_T_15[3:0] ? rowcount_8 : _GEN_580; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_582 = 4'h9 == _i_vn_1_T_15[3:0] ? rowcount_9 : _GEN_581; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_583 = 4'ha == _i_vn_1_T_15[3:0] ? rowcount_10 : _GEN_582; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_584 = 4'hb == _i_vn_1_T_15[3:0] ? rowcount_11 : _GEN_583; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_585 = 4'hc == _i_vn_1_T_15[3:0] ? rowcount_12 : _GEN_584; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_586 = 4'hd == _i_vn_1_T_15[3:0] ? rowcount_13 : _GEN_585; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_587 = 4'he == _i_vn_1_T_15[3:0] ? rowcount_14 : _GEN_586; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_588 = 4'hf == _i_vn_1_T_15[3:0] ? rowcount_15 : _GEN_587; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _T_172 = _GEN_268 + _GEN_588; // @[ivncontrol4.scala 275:41]
  wire [31:0] _T_174 = 32'h8 - _T_172; // @[ivncontrol4.scala 275:18]
  wire [31:0] _i_vn_1_T_17 = 32'h2 + pin; // @[ivncontrol4.scala 276:29]
  wire [31:0] _GEN_781 = _T_174 == 32'h1 ? _i_vn_1_T_17 : _GEN_556; // @[ivncontrol4.scala 318:78 321:22]
  wire [31:0] _GEN_782 = _T_174 == 32'h2 ? _i_vn_1_T_17 : _GEN_555; // @[ivncontrol4.scala 312:76 315:22]
  wire [31:0] _GEN_783 = _T_174 == 32'h2 ? _i_vn_1_T_17 : _GEN_781; // @[ivncontrol4.scala 312:76 316:22]
  wire [31:0] _GEN_784 = _T_174 == 32'h3 ? _i_vn_1_T_17 : _GEN_554; // @[ivncontrol4.scala 305:78 307:23]
  wire [31:0] _GEN_785 = _T_174 == 32'h3 ? _i_vn_1_T_17 : _GEN_782; // @[ivncontrol4.scala 305:78 308:22]
  wire [31:0] _GEN_786 = _T_174 == 32'h3 ? _i_vn_1_T_17 : _GEN_783; // @[ivncontrol4.scala 305:78 309:22]
  wire [31:0] _GEN_787 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_553; // @[ivncontrol4.scala 299:78 301:22]
  wire [31:0] _GEN_788 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_784; // @[ivncontrol4.scala 299:78 302:22]
  wire [31:0] _GEN_789 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_785; // @[ivncontrol4.scala 299:78 303:22]
  wire [31:0] _GEN_790 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_786; // @[ivncontrol4.scala 299:78 304:22]
  wire [31:0] _GEN_791 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_552; // @[ivncontrol4.scala 292:76 294:23]
  wire [31:0] _GEN_792 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_787; // @[ivncontrol4.scala 292:76 295:22]
  wire [31:0] _GEN_793 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_788; // @[ivncontrol4.scala 292:76 296:22]
  wire [31:0] _GEN_794 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_789; // @[ivncontrol4.scala 292:76 297:22]
  wire [31:0] _GEN_795 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_790; // @[ivncontrol4.scala 292:76 298:22]
  wire [31:0] _GEN_796 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_551; // @[ivncontrol4.scala 284:77 286:22]
  wire [31:0] _GEN_797 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_791; // @[ivncontrol4.scala 284:77 287:21]
  wire [31:0] _GEN_798 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_792; // @[ivncontrol4.scala 284:77 288:22]
  wire [31:0] _GEN_799 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_793; // @[ivncontrol4.scala 284:77 289:22]
  wire [31:0] _GEN_800 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_794; // @[ivncontrol4.scala 284:77 290:22]
  wire [31:0] _GEN_801 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_795; // @[ivncontrol4.scala 284:77 291:22]
  wire [31:0] _GEN_802 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_550; // @[ivncontrol4.scala 275:73 276:22]
  wire [31:0] _GEN_803 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_796; // @[ivncontrol4.scala 275:73 277:21]
  wire [31:0] _GEN_804 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_797; // @[ivncontrol4.scala 275:73 278:21]
  wire [31:0] _GEN_805 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_798; // @[ivncontrol4.scala 275:73 279:22]
  wire [31:0] _GEN_806 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_799; // @[ivncontrol4.scala 275:73 280:22]
  wire [31:0] _GEN_807 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_800; // @[ivncontrol4.scala 275:73 281:22]
  wire [31:0] _GEN_808 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_801; // @[ivncontrol4.scala 275:73 282:22]
  wire [31:0] _GEN_842 = 4'h1 == _i_vn_1_T_17[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_843 = 4'h2 == _i_vn_1_T_17[3:0] ? rowcount_2 : _GEN_842; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_844 = 4'h3 == _i_vn_1_T_17[3:0] ? rowcount_3 : _GEN_843; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_845 = 4'h4 == _i_vn_1_T_17[3:0] ? rowcount_4 : _GEN_844; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_846 = 4'h5 == _i_vn_1_T_17[3:0] ? rowcount_5 : _GEN_845; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_847 = 4'h6 == _i_vn_1_T_17[3:0] ? rowcount_6 : _GEN_846; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_848 = 4'h7 == _i_vn_1_T_17[3:0] ? rowcount_7 : _GEN_847; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_849 = 4'h8 == _i_vn_1_T_17[3:0] ? rowcount_8 : _GEN_848; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_850 = 4'h9 == _i_vn_1_T_17[3:0] ? rowcount_9 : _GEN_849; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_851 = 4'ha == _i_vn_1_T_17[3:0] ? rowcount_10 : _GEN_850; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_852 = 4'hb == _i_vn_1_T_17[3:0] ? rowcount_11 : _GEN_851; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_853 = 4'hc == _i_vn_1_T_17[3:0] ? rowcount_12 : _GEN_852; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_854 = 4'hd == _i_vn_1_T_17[3:0] ? rowcount_13 : _GEN_853; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_855 = 4'he == _i_vn_1_T_17[3:0] ? rowcount_14 : _GEN_854; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_856 = 4'hf == _i_vn_1_T_17[3:0] ? rowcount_15 : _GEN_855; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _T_254 = _T_172 + _GEN_856; // @[ivncontrol4.scala 326:62]
  wire [31:0] _T_256 = 32'h8 - _T_254; // @[ivncontrol4.scala 326:17]
  wire [31:0] _i_vn_1_T_19 = 32'h3 + pin; // @[ivncontrol4.scala 327:29]
  wire [31:0] _GEN_1145 = _T_256 == 32'h1 ? _i_vn_1_T_19 : _GEN_808; // @[ivncontrol4.scala 369:100 372:22]
  wire [31:0] _GEN_1146 = _T_256 == 32'h2 ? _i_vn_1_T_19 : _GEN_807; // @[ivncontrol4.scala 363:98 366:22]
  wire [31:0] _GEN_1147 = _T_256 == 32'h2 ? _i_vn_1_T_19 : _GEN_1145; // @[ivncontrol4.scala 363:98 367:22]
  wire [31:0] _GEN_1148 = _T_256 == 32'h3 ? _i_vn_1_T_19 : _GEN_806; // @[ivncontrol4.scala 356:100 358:23]
  wire [31:0] _GEN_1149 = _T_256 == 32'h3 ? _i_vn_1_T_19 : _GEN_1146; // @[ivncontrol4.scala 356:100 359:22]
  wire [31:0] _GEN_1150 = _T_256 == 32'h3 ? _i_vn_1_T_19 : _GEN_1147; // @[ivncontrol4.scala 356:100 360:22]
  wire [31:0] _GEN_1151 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_805; // @[ivncontrol4.scala 350:100 352:22]
  wire [31:0] _GEN_1152 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_1148; // @[ivncontrol4.scala 350:100 353:22]
  wire [31:0] _GEN_1153 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_1149; // @[ivncontrol4.scala 350:100 354:22]
  wire [31:0] _GEN_1154 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_1150; // @[ivncontrol4.scala 350:100 355:22]
  wire [31:0] _GEN_1155 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_804; // @[ivncontrol4.scala 343:98 345:23]
  wire [31:0] _GEN_1156 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1151; // @[ivncontrol4.scala 343:98 346:22]
  wire [31:0] _GEN_1157 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1152; // @[ivncontrol4.scala 343:98 347:22]
  wire [31:0] _GEN_1158 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1153; // @[ivncontrol4.scala 343:98 348:22]
  wire [31:0] _GEN_1159 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1154; // @[ivncontrol4.scala 343:98 349:22]
  wire [31:0] _GEN_1160 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_803; // @[ivncontrol4.scala 335:99 337:22]
  wire [31:0] _GEN_1161 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1155; // @[ivncontrol4.scala 335:99 338:21]
  wire [31:0] _GEN_1162 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1156; // @[ivncontrol4.scala 335:99 339:22]
  wire [31:0] _GEN_1163 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1157; // @[ivncontrol4.scala 335:99 340:22]
  wire [31:0] _GEN_1164 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1158; // @[ivncontrol4.scala 335:99 341:22]
  wire [31:0] _GEN_1165 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1159; // @[ivncontrol4.scala 335:99 342:22]
  wire [31:0] _GEN_1166 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_802; // @[ivncontrol4.scala 326:94 327:22]
  wire [31:0] _GEN_1167 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1160; // @[ivncontrol4.scala 326:94 328:21]
  wire [31:0] _GEN_1168 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1161; // @[ivncontrol4.scala 326:94 329:21]
  wire [31:0] _GEN_1169 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1162; // @[ivncontrol4.scala 326:94 330:22]
  wire [31:0] _GEN_1170 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1163; // @[ivncontrol4.scala 326:94 331:22]
  wire [31:0] _GEN_1171 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1164; // @[ivncontrol4.scala 326:94 332:22]
  wire [31:0] _GEN_1172 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1165; // @[ivncontrol4.scala 326:94 333:22]
  wire [31:0] _GEN_1222 = 4'h1 == _i_vn_1_T_19[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1223 = 4'h2 == _i_vn_1_T_19[3:0] ? rowcount_2 : _GEN_1222; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1224 = 4'h3 == _i_vn_1_T_19[3:0] ? rowcount_3 : _GEN_1223; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1225 = 4'h4 == _i_vn_1_T_19[3:0] ? rowcount_4 : _GEN_1224; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1226 = 4'h5 == _i_vn_1_T_19[3:0] ? rowcount_5 : _GEN_1225; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1227 = 4'h6 == _i_vn_1_T_19[3:0] ? rowcount_6 : _GEN_1226; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1228 = 4'h7 == _i_vn_1_T_19[3:0] ? rowcount_7 : _GEN_1227; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1229 = 4'h8 == _i_vn_1_T_19[3:0] ? rowcount_8 : _GEN_1228; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1230 = 4'h9 == _i_vn_1_T_19[3:0] ? rowcount_9 : _GEN_1229; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1231 = 4'ha == _i_vn_1_T_19[3:0] ? rowcount_10 : _GEN_1230; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1232 = 4'hb == _i_vn_1_T_19[3:0] ? rowcount_11 : _GEN_1231; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1233 = 4'hc == _i_vn_1_T_19[3:0] ? rowcount_12 : _GEN_1232; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1234 = 4'hd == _i_vn_1_T_19[3:0] ? rowcount_13 : _GEN_1233; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1235 = 4'he == _i_vn_1_T_19[3:0] ? rowcount_14 : _GEN_1234; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1236 = 4'hf == _i_vn_1_T_19[3:0] ? rowcount_15 : _GEN_1235; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _T_371 = _T_254 + _GEN_1236; // @[ivncontrol4.scala 376:86]
  wire [31:0] _T_373 = 32'h8 - _T_371; // @[ivncontrol4.scala 376:19]
  wire [31:0] _i_vn_1_T_21 = 32'h4 + pin; // @[ivncontrol4.scala 377:29]
  wire [31:0] _GEN_1621 = _T_373 == 32'h1 ? _i_vn_1_T_21 : _GEN_1172; // @[ivncontrol4.scala 419:122 422:22]
  wire [31:0] _GEN_1622 = _T_373 == 32'h2 ? _i_vn_1_T_21 : _GEN_1171; // @[ivncontrol4.scala 413:121 416:22]
  wire [31:0] _GEN_1623 = _T_373 == 32'h2 ? _i_vn_1_T_21 : _GEN_1621; // @[ivncontrol4.scala 413:121 417:22]
  wire [31:0] _GEN_1624 = _T_373 == 32'h3 ? _i_vn_1_T_21 : _GEN_1170; // @[ivncontrol4.scala 406:123 408:23]
  wire [31:0] _GEN_1625 = _T_373 == 32'h3 ? _i_vn_1_T_21 : _GEN_1622; // @[ivncontrol4.scala 406:123 409:22]
  wire [31:0] _GEN_1626 = _T_373 == 32'h3 ? _i_vn_1_T_21 : _GEN_1623; // @[ivncontrol4.scala 406:123 410:22]
  wire [31:0] _GEN_1627 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1169; // @[ivncontrol4.scala 400:122 402:22]
  wire [31:0] _GEN_1628 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1624; // @[ivncontrol4.scala 400:122 403:22]
  wire [31:0] _GEN_1629 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1625; // @[ivncontrol4.scala 400:122 404:22]
  wire [31:0] _GEN_1630 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1626; // @[ivncontrol4.scala 400:122 405:22]
  wire [31:0] _GEN_1631 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1168; // @[ivncontrol4.scala 393:121 395:23]
  wire [31:0] _GEN_1632 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1627; // @[ivncontrol4.scala 393:121 396:22]
  wire [31:0] _GEN_1633 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1628; // @[ivncontrol4.scala 393:121 397:22]
  wire [31:0] _GEN_1634 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1629; // @[ivncontrol4.scala 393:121 398:22]
  wire [31:0] _GEN_1635 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1630; // @[ivncontrol4.scala 393:121 399:22]
  wire [31:0] _GEN_1636 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1167; // @[ivncontrol4.scala 385:121 387:22]
  wire [31:0] _GEN_1637 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1631; // @[ivncontrol4.scala 385:121 388:21]
  wire [31:0] _GEN_1638 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1632; // @[ivncontrol4.scala 385:121 389:22]
  wire [31:0] _GEN_1639 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1633; // @[ivncontrol4.scala 385:121 390:22]
  wire [31:0] _GEN_1640 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1634; // @[ivncontrol4.scala 385:121 391:22]
  wire [31:0] _GEN_1641 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1635; // @[ivncontrol4.scala 385:121 392:22]
  wire [31:0] _GEN_1642 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1166; // @[ivncontrol4.scala 376:118 377:22]
  wire [31:0] _GEN_1643 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1636; // @[ivncontrol4.scala 376:118 378:21]
  wire [31:0] _GEN_1644 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1637; // @[ivncontrol4.scala 376:118 379:21]
  wire [31:0] _GEN_1645 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1638; // @[ivncontrol4.scala 376:118 380:22]
  wire [31:0] _GEN_1646 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1639; // @[ivncontrol4.scala 376:118 381:22]
  wire [31:0] _GEN_1647 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1640; // @[ivncontrol4.scala 376:118 382:22]
  wire [31:0] _GEN_1648 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1641; // @[ivncontrol4.scala 376:118 383:22]
  wire [31:0] _GEN_1714 = 4'h1 == _i_vn_1_T_21[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1715 = 4'h2 == _i_vn_1_T_21[3:0] ? rowcount_2 : _GEN_1714; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1716 = 4'h3 == _i_vn_1_T_21[3:0] ? rowcount_3 : _GEN_1715; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1717 = 4'h4 == _i_vn_1_T_21[3:0] ? rowcount_4 : _GEN_1716; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1718 = 4'h5 == _i_vn_1_T_21[3:0] ? rowcount_5 : _GEN_1717; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1719 = 4'h6 == _i_vn_1_T_21[3:0] ? rowcount_6 : _GEN_1718; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1720 = 4'h7 == _i_vn_1_T_21[3:0] ? rowcount_7 : _GEN_1719; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1721 = 4'h8 == _i_vn_1_T_21[3:0] ? rowcount_8 : _GEN_1720; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1722 = 4'h9 == _i_vn_1_T_21[3:0] ? rowcount_9 : _GEN_1721; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1723 = 4'ha == _i_vn_1_T_21[3:0] ? rowcount_10 : _GEN_1722; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1724 = 4'hb == _i_vn_1_T_21[3:0] ? rowcount_11 : _GEN_1723; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1725 = 4'hc == _i_vn_1_T_21[3:0] ? rowcount_12 : _GEN_1724; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1726 = 4'hd == _i_vn_1_T_21[3:0] ? rowcount_13 : _GEN_1725; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1727 = 4'he == _i_vn_1_T_21[3:0] ? rowcount_14 : _GEN_1726; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1728 = 4'hf == _i_vn_1_T_21[3:0] ? rowcount_15 : _GEN_1727; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _T_523 = _T_371 + _GEN_1728; // @[ivncontrol4.scala 426:108]
  wire [31:0] _T_525 = 32'h8 - _T_523; // @[ivncontrol4.scala 426:19]
  wire [31:0] _i_vn_1_T_23 = 32'h5 + pin; // @[ivncontrol4.scala 427:29]
  wire [31:0] _GEN_2209 = _T_525 == 32'h1 ? _i_vn_1_T_23 : _GEN_1648; // @[ivncontrol4.scala 469:144 472:22]
  wire [31:0] _GEN_2210 = _T_525 == 32'h2 ? _i_vn_1_T_23 : _GEN_1647; // @[ivncontrol4.scala 463:143 466:22]
  wire [31:0] _GEN_2211 = _T_525 == 32'h2 ? _i_vn_1_T_23 : _GEN_2209; // @[ivncontrol4.scala 463:143 467:22]
  wire [31:0] _GEN_2212 = _T_525 == 32'h3 ? _i_vn_1_T_23 : _GEN_1646; // @[ivncontrol4.scala 456:145 458:23]
  wire [31:0] _GEN_2213 = _T_525 == 32'h3 ? _i_vn_1_T_23 : _GEN_2210; // @[ivncontrol4.scala 456:145 459:22]
  wire [31:0] _GEN_2214 = _T_525 == 32'h3 ? _i_vn_1_T_23 : _GEN_2211; // @[ivncontrol4.scala 456:145 460:22]
  wire [31:0] _GEN_2215 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_1645; // @[ivncontrol4.scala 450:143 452:22]
  wire [31:0] _GEN_2216 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_2212; // @[ivncontrol4.scala 450:143 453:22]
  wire [31:0] _GEN_2217 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_2213; // @[ivncontrol4.scala 450:143 454:22]
  wire [31:0] _GEN_2218 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_2214; // @[ivncontrol4.scala 450:143 455:22]
  wire [31:0] _GEN_2219 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_1644; // @[ivncontrol4.scala 443:143 445:23]
  wire [31:0] _GEN_2220 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2215; // @[ivncontrol4.scala 443:143 446:22]
  wire [31:0] _GEN_2221 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2216; // @[ivncontrol4.scala 443:143 447:22]
  wire [31:0] _GEN_2222 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2217; // @[ivncontrol4.scala 443:143 448:22]
  wire [31:0] _GEN_2223 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2218; // @[ivncontrol4.scala 443:143 449:22]
  wire [31:0] _GEN_2224 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_1643; // @[ivncontrol4.scala 435:143 437:22]
  wire [31:0] _GEN_2225 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2219; // @[ivncontrol4.scala 435:143 438:21]
  wire [31:0] _GEN_2226 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2220; // @[ivncontrol4.scala 435:143 439:22]
  wire [31:0] _GEN_2227 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2221; // @[ivncontrol4.scala 435:143 440:22]
  wire [31:0] _GEN_2228 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2222; // @[ivncontrol4.scala 435:143 441:22]
  wire [31:0] _GEN_2229 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2223; // @[ivncontrol4.scala 435:143 442:22]
  wire [31:0] _GEN_2230 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_1642; // @[ivncontrol4.scala 426:140 427:22]
  wire [31:0] _GEN_2231 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2224; // @[ivncontrol4.scala 426:140 428:21]
  wire [31:0] _GEN_2232 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2225; // @[ivncontrol4.scala 426:140 429:21]
  wire [31:0] _GEN_2233 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2226; // @[ivncontrol4.scala 426:140 430:22]
  wire [31:0] _GEN_2234 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2227; // @[ivncontrol4.scala 426:140 431:22]
  wire [31:0] _GEN_2235 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2228; // @[ivncontrol4.scala 426:140 432:22]
  wire [31:0] _GEN_2236 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2229; // @[ivncontrol4.scala 426:140 433:22]
  wire [31:0] _GEN_2318 = 4'h1 == _i_vn_1_T_23[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2319 = 4'h2 == _i_vn_1_T_23[3:0] ? rowcount_2 : _GEN_2318; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2320 = 4'h3 == _i_vn_1_T_23[3:0] ? rowcount_3 : _GEN_2319; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2321 = 4'h4 == _i_vn_1_T_23[3:0] ? rowcount_4 : _GEN_2320; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2322 = 4'h5 == _i_vn_1_T_23[3:0] ? rowcount_5 : _GEN_2321; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2323 = 4'h6 == _i_vn_1_T_23[3:0] ? rowcount_6 : _GEN_2322; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2324 = 4'h7 == _i_vn_1_T_23[3:0] ? rowcount_7 : _GEN_2323; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2325 = 4'h8 == _i_vn_1_T_23[3:0] ? rowcount_8 : _GEN_2324; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2326 = 4'h9 == _i_vn_1_T_23[3:0] ? rowcount_9 : _GEN_2325; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2327 = 4'ha == _i_vn_1_T_23[3:0] ? rowcount_10 : _GEN_2326; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2328 = 4'hb == _i_vn_1_T_23[3:0] ? rowcount_11 : _GEN_2327; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2329 = 4'hc == _i_vn_1_T_23[3:0] ? rowcount_12 : _GEN_2328; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2330 = 4'hd == _i_vn_1_T_23[3:0] ? rowcount_13 : _GEN_2329; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2331 = 4'he == _i_vn_1_T_23[3:0] ? rowcount_14 : _GEN_2330; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2332 = 4'hf == _i_vn_1_T_23[3:0] ? rowcount_15 : _GEN_2331; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _T_710 = _T_523 + _GEN_2332; // @[ivncontrol4.scala 477:130]
  wire [31:0] _T_712 = 32'h8 - _T_710; // @[ivncontrol4.scala 477:19]
  wire [31:0] _i_vn_1_T_25 = 32'h6 + pin; // @[ivncontrol4.scala 478:29]
  wire [31:0] _GEN_2909 = _T_712 == 32'h1 ? _i_vn_1_T_25 : _GEN_2236; // @[ivncontrol4.scala 520:166 523:22]
  wire [31:0] _GEN_2910 = _T_712 == 32'h2 ? _i_vn_1_T_25 : _GEN_2235; // @[ivncontrol4.scala 514:166 517:22]
  wire [31:0] _GEN_2911 = _T_712 == 32'h2 ? _i_vn_1_T_25 : _GEN_2909; // @[ivncontrol4.scala 514:166 518:22]
  wire [31:0] _GEN_2912 = _T_712 == 32'h3 ? _i_vn_1_T_25 : _GEN_2234; // @[ivncontrol4.scala 507:168 509:23]
  wire [31:0] _GEN_2913 = _T_712 == 32'h3 ? _i_vn_1_T_25 : _GEN_2910; // @[ivncontrol4.scala 507:168 510:22]
  wire [31:0] _GEN_2914 = _T_712 == 32'h3 ? _i_vn_1_T_25 : _GEN_2911; // @[ivncontrol4.scala 507:168 511:22]
  wire [31:0] _GEN_2915 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2233; // @[ivncontrol4.scala 501:166 503:22]
  wire [31:0] _GEN_2916 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2912; // @[ivncontrol4.scala 501:166 504:22]
  wire [31:0] _GEN_2917 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2913; // @[ivncontrol4.scala 501:166 505:22]
  wire [31:0] _GEN_2918 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2914; // @[ivncontrol4.scala 501:166 506:22]
  wire [31:0] _GEN_2919 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2232; // @[ivncontrol4.scala 494:166 496:23]
  wire [31:0] _GEN_2920 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2915; // @[ivncontrol4.scala 494:166 497:22]
  wire [31:0] _GEN_2921 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2916; // @[ivncontrol4.scala 494:166 498:22]
  wire [31:0] _GEN_2922 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2917; // @[ivncontrol4.scala 494:166 499:22]
  wire [31:0] _GEN_2923 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2918; // @[ivncontrol4.scala 494:166 500:22]
  wire [31:0] _GEN_2924 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2231; // @[ivncontrol4.scala 486:166 488:22]
  wire [31:0] _GEN_2925 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2919; // @[ivncontrol4.scala 486:166 489:21]
  wire [31:0] _GEN_2926 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2920; // @[ivncontrol4.scala 486:166 490:22]
  wire [31:0] _GEN_2927 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2921; // @[ivncontrol4.scala 486:166 491:22]
  wire [31:0] _GEN_2928 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2922; // @[ivncontrol4.scala 486:166 492:22]
  wire [31:0] _GEN_2929 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2923; // @[ivncontrol4.scala 486:166 493:22]
  wire [31:0] _GEN_2930 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2230; // @[ivncontrol4.scala 477:162 478:22]
  wire [31:0] _GEN_2931 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2924; // @[ivncontrol4.scala 477:162 479:21]
  wire [31:0] _GEN_2932 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2925; // @[ivncontrol4.scala 477:162 480:21]
  wire [31:0] _GEN_2933 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2926; // @[ivncontrol4.scala 477:162 481:22]
  wire [31:0] _GEN_2934 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2927; // @[ivncontrol4.scala 477:162 482:22]
  wire [31:0] _GEN_2935 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2928; // @[ivncontrol4.scala 477:162 483:22]
  wire [31:0] _GEN_2936 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2929; // @[ivncontrol4.scala 477:162 484:22]
  wire [31:0] _GEN_3034 = 4'h1 == _i_vn_1_T_25[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3035 = 4'h2 == _i_vn_1_T_25[3:0] ? rowcount_2 : _GEN_3034; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3036 = 4'h3 == _i_vn_1_T_25[3:0] ? rowcount_3 : _GEN_3035; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3037 = 4'h4 == _i_vn_1_T_25[3:0] ? rowcount_4 : _GEN_3036; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3038 = 4'h5 == _i_vn_1_T_25[3:0] ? rowcount_5 : _GEN_3037; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3039 = 4'h6 == _i_vn_1_T_25[3:0] ? rowcount_6 : _GEN_3038; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3040 = 4'h7 == _i_vn_1_T_25[3:0] ? rowcount_7 : _GEN_3039; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3041 = 4'h8 == _i_vn_1_T_25[3:0] ? rowcount_8 : _GEN_3040; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3042 = 4'h9 == _i_vn_1_T_25[3:0] ? rowcount_9 : _GEN_3041; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3043 = 4'ha == _i_vn_1_T_25[3:0] ? rowcount_10 : _GEN_3042; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3044 = 4'hb == _i_vn_1_T_25[3:0] ? rowcount_11 : _GEN_3043; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3045 = 4'hc == _i_vn_1_T_25[3:0] ? rowcount_12 : _GEN_3044; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3046 = 4'hd == _i_vn_1_T_25[3:0] ? rowcount_13 : _GEN_3045; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3047 = 4'he == _i_vn_1_T_25[3:0] ? rowcount_14 : _GEN_3046; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3048 = 4'hf == _i_vn_1_T_25[3:0] ? rowcount_15 : _GEN_3047; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _T_932 = _T_710 + _GEN_3048; // @[ivncontrol4.scala 528:152]
  wire [31:0] _T_934 = 32'h8 - _T_932; // @[ivncontrol4.scala 528:19]
  wire [31:0] _i_vn_1_T_27 = 32'h7 + pin; // @[ivncontrol4.scala 529:29]
  wire [31:0] _GEN_3721 = _T_934 == 32'h1 ? _i_vn_1_T_27 : _GEN_2936; // @[ivncontrol4.scala 571:188 574:22]
  wire [31:0] _GEN_3722 = _T_934 == 32'h2 ? _i_vn_1_T_27 : _GEN_2935; // @[ivncontrol4.scala 565:188 568:22]
  wire [31:0] _GEN_3723 = _T_934 == 32'h2 ? _i_vn_1_T_27 : _GEN_3721; // @[ivncontrol4.scala 565:188 569:22]
  wire [31:0] _GEN_3724 = _T_934 == 32'h3 ? _i_vn_1_T_27 : _GEN_2934; // @[ivncontrol4.scala 558:190 560:23]
  wire [31:0] _GEN_3725 = _T_934 == 32'h3 ? _i_vn_1_T_27 : _GEN_3722; // @[ivncontrol4.scala 558:190 561:22]
  wire [31:0] _GEN_3726 = _T_934 == 32'h3 ? _i_vn_1_T_27 : _GEN_3723; // @[ivncontrol4.scala 558:190 562:22]
  wire [31:0] _GEN_3727 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_2933; // @[ivncontrol4.scala 552:188 554:22]
  wire [31:0] _GEN_3728 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_3724; // @[ivncontrol4.scala 552:188 555:22]
  wire [31:0] _GEN_3729 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_3725; // @[ivncontrol4.scala 552:188 556:22]
  wire [31:0] _GEN_3730 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_3726; // @[ivncontrol4.scala 552:188 557:22]
  wire [31:0] _GEN_3731 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_2932; // @[ivncontrol4.scala 545:188 547:23]
  wire [31:0] _GEN_3732 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3727; // @[ivncontrol4.scala 545:188 548:22]
  wire [31:0] _GEN_3733 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3728; // @[ivncontrol4.scala 545:188 549:22]
  wire [31:0] _GEN_3734 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3729; // @[ivncontrol4.scala 545:188 550:22]
  wire [31:0] _GEN_3735 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3730; // @[ivncontrol4.scala 545:188 551:22]
  wire [31:0] _GEN_3736 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_2931; // @[ivncontrol4.scala 537:188 539:22]
  wire [31:0] _GEN_3737 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3731; // @[ivncontrol4.scala 537:188 540:21]
  wire [31:0] _GEN_3738 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3732; // @[ivncontrol4.scala 537:188 541:22]
  wire [31:0] _GEN_3739 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3733; // @[ivncontrol4.scala 537:188 542:22]
  wire [31:0] _GEN_3740 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3734; // @[ivncontrol4.scala 537:188 543:22]
  wire [31:0] _GEN_3741 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3735; // @[ivncontrol4.scala 537:188 544:22]
  wire [31:0] _GEN_3742 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_2930; // @[ivncontrol4.scala 528:184 529:22]
  wire [31:0] _GEN_3743 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3736; // @[ivncontrol4.scala 528:184 530:21]
  wire [31:0] _GEN_3744 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3737; // @[ivncontrol4.scala 528:184 531:21]
  wire [31:0] _GEN_3745 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3738; // @[ivncontrol4.scala 528:184 532:22]
  wire [31:0] _GEN_3746 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3739; // @[ivncontrol4.scala 528:184 533:22]
  wire [31:0] _GEN_3747 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3740; // @[ivncontrol4.scala 528:184 534:22]
  wire [31:0] _GEN_3748 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3741; // @[ivncontrol4.scala 528:184 535:22]
  wire [31:0] _GEN_3749 = _GEN_244 ? _GEN_409 : 32'h19; // @[ivncontrol4.scala 125:17 172:28]
  wire [31:0] _GEN_3750 = _GEN_244 ? _GEN_3742 : 32'ha; // @[ivncontrol4.scala 125:17 172:28]
  wire [31:0] _GEN_3751 = _GEN_244 ? _GEN_3743 : 32'he; // @[ivncontrol4.scala 125:17 172:28]
  wire [31:0] _GEN_3752 = _GEN_244 ? _GEN_3744 : 32'h4; // @[ivncontrol4.scala 125:17 172:28]
  wire [31:0] _GEN_3753 = _GEN_244 ? _GEN_3745 : 32'h10; // @[ivncontrol4.scala 126:18 172:28]
  wire [31:0] _GEN_3754 = _GEN_244 ? _GEN_3746 : 32'he; // @[ivncontrol4.scala 126:18 172:28]
  wire [31:0] _GEN_3755 = _GEN_244 ? _GEN_3747 : 32'ha; // @[ivncontrol4.scala 126:18 172:28]
  wire [31:0] _GEN_3756 = _GEN_244 ? _GEN_3748 : 32'h1; // @[ivncontrol4.scala 126:18 172:28]
  wire [31:0] _GEN_4137 = reset ? 32'h0 : _GEN_3749; // @[ivncontrol4.scala 16:{23,23}]
  wire [31:0] _GEN_4138 = reset ? 32'h0 : _GEN_3750; // @[ivncontrol4.scala 16:{23,23}]
  wire [31:0] _GEN_4139 = reset ? 32'h0 : _GEN_3751; // @[ivncontrol4.scala 16:{23,23}]
  wire [31:0] _GEN_4140 = reset ? 32'h0 : _GEN_3752; // @[ivncontrol4.scala 16:{23,23}]
  wire [31:0] _GEN_4141 = reset ? 32'h0 : _GEN_3753; // @[ivncontrol4.scala 17:{24,24}]
  wire [31:0] _GEN_4142 = reset ? 32'h0 : _GEN_3754; // @[ivncontrol4.scala 17:{24,24}]
  wire [31:0] _GEN_4143 = reset ? 32'h0 : _GEN_3755; // @[ivncontrol4.scala 17:{24,24}]
  wire [31:0] _GEN_4144 = reset ? 32'h0 : _GEN_3756; // @[ivncontrol4.scala 17:{24,24}]
  assign io_o_vn_0 = i_vn_0; // @[ivncontrol4.scala 121:13]
  assign io_o_vn_1 = i_vn_1; // @[ivncontrol4.scala 121:13]
  assign io_o_vn_2 = i_vn_2; // @[ivncontrol4.scala 121:13]
  assign io_o_vn_3 = i_vn_3; // @[ivncontrol4.scala 121:13]
  assign io_o_vn2_0 = i_vn2_0; // @[ivncontrol4.scala 122:14]
  assign io_o_vn2_1 = i_vn2_1; // @[ivncontrol4.scala 122:14]
  assign io_o_vn2_2 = i_vn2_2; // @[ivncontrol4.scala 122:14]
  assign io_o_vn2_3 = i_vn2_3; // @[ivncontrol4.scala 122:14]
  always @(posedge clock) begin
    i_vn_0 <= _GEN_4137[4:0]; // @[ivncontrol4.scala 16:{23,23}]
    i_vn_1 <= _GEN_4138[4:0]; // @[ivncontrol4.scala 16:{23,23}]
    i_vn_2 <= _GEN_4139[4:0]; // @[ivncontrol4.scala 16:{23,23}]
    i_vn_3 <= _GEN_4140[4:0]; // @[ivncontrol4.scala 16:{23,23}]
    i_vn2_0 <= _GEN_4141[4:0]; // @[ivncontrol4.scala 17:{24,24}]
    i_vn2_1 <= _GEN_4142[4:0]; // @[ivncontrol4.scala 17:{24,24}]
    i_vn2_2 <= _GEN_4143[4:0]; // @[ivncontrol4.scala 17:{24,24}]
    i_vn2_3 <= _GEN_4144[4:0]; // @[ivncontrol4.scala 17:{24,24}]
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_0 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_0 <= count_0; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_1 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_1 <= count_1; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_2 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_2 <= count_2; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_3 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_3 <= count_3; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_4 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_4 <= count_4; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_5 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_5 <= count_5; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_6 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_6 <= count_6; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_7 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_7 <= count_7; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_8 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_8 <= 32'h0; // @[ivncontrol4.scala 81:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_9 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_9 <= 32'h0; // @[ivncontrol4.scala 81:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_10 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_10 <= 32'h0; // @[ivncontrol4.scala 81:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_11 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_11 <= 32'h0; // @[ivncontrol4.scala 81:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_12 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_12 <= 32'h0; // @[ivncontrol4.scala 81:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_13 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_13 <= 32'h0; // @[ivncontrol4.scala 81:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_14 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_14 <= 32'h0; // @[ivncontrol4.scala 81:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_15 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end
    if (reset) begin // @[ivncontrol4.scala 31:22]
      pin <= 32'h0; // @[ivncontrol4.scala 31:22]
    end else if (_T_72 & rowcount_6 == 32'h0 & rowcount_7 != 32'h0) begin // @[ivncontrol4.scala 166:192]
      pin <= 32'h7; // @[ivncontrol4.scala 167:13]
    end else if (_T_59 & rowcount_5 == 32'h0 & rowcount_6 != 32'h0) begin // @[ivncontrol4.scala 163:169]
      pin <= 32'h6; // @[ivncontrol4.scala 164:13]
    end else if (_T_48 & rowcount_4 == 32'h0 & rowcount_5 != 32'h0) begin // @[ivncontrol4.scala 160:146]
      pin <= 32'h5; // @[ivncontrol4.scala 161:13]
    end else begin
      pin <= _GEN_249;
    end
    if (reset) begin // @[ivncontrol4.scala 35:20]
      i <= 32'h0; // @[ivncontrol4.scala 35:20]
    end else if (i < 32'h7 & _k_T_1) begin // @[ivncontrol4.scala 103:74]
      i <= _i_T_1; // @[ivncontrol4.scala 104:11]
    end
    if (reset) begin // @[ivncontrol4.scala 36:20]
      j <= 32'h0; // @[ivncontrol4.scala 36:20]
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 107:71]
      j <= _j_T_1; // @[ivncontrol4.scala 108:11]
    end else if (!(_k_T_2)) begin // @[ivncontrol4.scala 110:81]
      j <= 32'h0; // @[ivncontrol4.scala 114:11]
    end
    if (3'h0 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h0 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h0 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h0 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h0 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h0 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h0 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h0 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h0 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_0 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h1 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_1 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h2 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_2 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h3 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_3 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h4 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_4 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h5 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_5 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h6 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_6 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h7 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_7 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  i_vn_0 = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  i_vn_1 = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  i_vn_2 = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  i_vn_3 = _RAND_3[4:0];
  _RAND_4 = {1{`RANDOM}};
  i_vn2_0 = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  i_vn2_1 = _RAND_5[4:0];
  _RAND_6 = {1{`RANDOM}};
  i_vn2_2 = _RAND_6[4:0];
  _RAND_7 = {1{`RANDOM}};
  i_vn2_3 = _RAND_7[4:0];
  _RAND_8 = {1{`RANDOM}};
  rowcount_0 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  rowcount_1 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  rowcount_2 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  rowcount_3 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  rowcount_4 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  rowcount_5 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  rowcount_6 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  rowcount_7 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  rowcount_8 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  rowcount_9 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  rowcount_10 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  rowcount_11 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  rowcount_12 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  rowcount_13 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  rowcount_14 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  rowcount_15 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  pin = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  i = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  j = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  mat_0_0 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  mat_0_1 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  mat_0_2 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  mat_0_3 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  mat_0_4 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  mat_0_5 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  mat_0_6 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  mat_0_7 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  mat_1_0 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  mat_1_1 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  mat_1_2 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  mat_1_3 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  mat_1_4 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  mat_1_5 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  mat_1_6 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  mat_1_7 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  mat_2_0 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  mat_2_1 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  mat_2_2 = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  mat_2_3 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  mat_2_4 = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  mat_2_5 = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  mat_2_6 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  mat_2_7 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  mat_3_0 = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  mat_3_1 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  mat_3_2 = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  mat_3_3 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  mat_3_4 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  mat_3_5 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  mat_3_6 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  mat_3_7 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  mat_4_0 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  mat_4_1 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  mat_4_2 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  mat_4_3 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  mat_4_4 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  mat_4_5 = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  mat_4_6 = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  mat_4_7 = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  mat_5_0 = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  mat_5_1 = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  mat_5_2 = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  mat_5_3 = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  mat_5_4 = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  mat_5_5 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  mat_5_6 = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  mat_5_7 = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  mat_6_0 = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  mat_6_1 = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  mat_6_2 = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  mat_6_3 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  mat_6_4 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  mat_6_5 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  mat_6_6 = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  mat_6_7 = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  mat_7_0 = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  mat_7_1 = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  mat_7_2 = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  mat_7_3 = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  mat_7_4 = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  mat_7_5 = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  mat_7_6 = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  mat_7_7 = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  count_0 = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  count_1 = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  count_2 = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  count_3 = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  count_4 = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  count_5 = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  count_6 = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  count_7 = _RAND_98[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ivncontrol4_5(
  input         clock,
  input         reset,
  input  [15:0] io_Stationary_matrix_0_0,
  input  [15:0] io_Stationary_matrix_0_1,
  input  [15:0] io_Stationary_matrix_0_2,
  input  [15:0] io_Stationary_matrix_0_3,
  input  [15:0] io_Stationary_matrix_0_4,
  input  [15:0] io_Stationary_matrix_0_5,
  input  [15:0] io_Stationary_matrix_0_6,
  input  [15:0] io_Stationary_matrix_0_7,
  input  [15:0] io_Stationary_matrix_1_0,
  input  [15:0] io_Stationary_matrix_1_1,
  input  [15:0] io_Stationary_matrix_1_2,
  input  [15:0] io_Stationary_matrix_1_3,
  input  [15:0] io_Stationary_matrix_1_4,
  input  [15:0] io_Stationary_matrix_1_5,
  input  [15:0] io_Stationary_matrix_1_6,
  input  [15:0] io_Stationary_matrix_1_7,
  input  [15:0] io_Stationary_matrix_2_0,
  input  [15:0] io_Stationary_matrix_2_1,
  input  [15:0] io_Stationary_matrix_2_2,
  input  [15:0] io_Stationary_matrix_2_3,
  input  [15:0] io_Stationary_matrix_2_4,
  input  [15:0] io_Stationary_matrix_2_5,
  input  [15:0] io_Stationary_matrix_2_6,
  input  [15:0] io_Stationary_matrix_2_7,
  input  [15:0] io_Stationary_matrix_3_0,
  input  [15:0] io_Stationary_matrix_3_1,
  input  [15:0] io_Stationary_matrix_3_2,
  input  [15:0] io_Stationary_matrix_3_3,
  input  [15:0] io_Stationary_matrix_3_4,
  input  [15:0] io_Stationary_matrix_3_5,
  input  [15:0] io_Stationary_matrix_3_6,
  input  [15:0] io_Stationary_matrix_3_7,
  input  [15:0] io_Stationary_matrix_4_0,
  input  [15:0] io_Stationary_matrix_4_1,
  input  [15:0] io_Stationary_matrix_4_2,
  input  [15:0] io_Stationary_matrix_4_3,
  input  [15:0] io_Stationary_matrix_4_4,
  input  [15:0] io_Stationary_matrix_4_5,
  input  [15:0] io_Stationary_matrix_4_6,
  input  [15:0] io_Stationary_matrix_4_7,
  input  [15:0] io_Stationary_matrix_5_0,
  input  [15:0] io_Stationary_matrix_5_1,
  input  [15:0] io_Stationary_matrix_5_2,
  input  [15:0] io_Stationary_matrix_5_3,
  input  [15:0] io_Stationary_matrix_5_4,
  input  [15:0] io_Stationary_matrix_5_5,
  input  [15:0] io_Stationary_matrix_5_6,
  input  [15:0] io_Stationary_matrix_5_7,
  input  [15:0] io_Stationary_matrix_6_0,
  input  [15:0] io_Stationary_matrix_6_1,
  input  [15:0] io_Stationary_matrix_6_2,
  input  [15:0] io_Stationary_matrix_6_3,
  input  [15:0] io_Stationary_matrix_6_4,
  input  [15:0] io_Stationary_matrix_6_5,
  input  [15:0] io_Stationary_matrix_6_6,
  input  [15:0] io_Stationary_matrix_6_7,
  input  [15:0] io_Stationary_matrix_7_0,
  input  [15:0] io_Stationary_matrix_7_1,
  input  [15:0] io_Stationary_matrix_7_2,
  input  [15:0] io_Stationary_matrix_7_3,
  input  [15:0] io_Stationary_matrix_7_4,
  input  [15:0] io_Stationary_matrix_7_5,
  input  [15:0] io_Stationary_matrix_7_6,
  input  [15:0] io_Stationary_matrix_7_7,
  output [4:0]  io_o_vn_0,
  output [4:0]  io_o_vn_1,
  output [4:0]  io_o_vn_2,
  output [4:0]  io_o_vn_3,
  output [4:0]  io_o_vn2_0,
  output [4:0]  io_o_vn2_1,
  output [4:0]  io_o_vn2_2,
  output [4:0]  io_o_vn2_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
`endif // RANDOMIZE_REG_INIT
  reg [4:0] i_vn_0; // @[ivncontrol4.scala 16:23]
  reg [4:0] i_vn_1; // @[ivncontrol4.scala 16:23]
  reg [4:0] i_vn_2; // @[ivncontrol4.scala 16:23]
  reg [4:0] i_vn_3; // @[ivncontrol4.scala 16:23]
  reg [4:0] i_vn2_0; // @[ivncontrol4.scala 17:24]
  reg [4:0] i_vn2_1; // @[ivncontrol4.scala 17:24]
  reg [4:0] i_vn2_2; // @[ivncontrol4.scala 17:24]
  reg [4:0] i_vn2_3; // @[ivncontrol4.scala 17:24]
  reg [31:0] rowcount_0; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_1; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_2; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_3; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_4; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_5; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_6; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_7; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_8; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_9; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_10; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_11; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_12; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_13; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_14; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_15; // @[ivncontrol4.scala 21:27]
  reg [31:0] pin; // @[ivncontrol4.scala 31:22]
  reg [31:0] i; // @[ivncontrol4.scala 35:20]
  reg [31:0] j; // @[ivncontrol4.scala 36:20]
  wire  _k_T_1 = j == 32'h7; // @[ivncontrol4.scala 38:37]
  wire  _k_T_2 = i == 32'h7 & j == 32'h7; // @[ivncontrol4.scala 38:31]
  reg [31:0] mat_0_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_0_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_0_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_0_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_0_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_0_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_0_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_0_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] count_0; // @[ivncontrol4.scala 52:20]
  reg [31:0] count_1; // @[ivncontrol4.scala 52:20]
  reg [31:0] count_2; // @[ivncontrol4.scala 52:20]
  reg [31:0] count_3; // @[ivncontrol4.scala 52:20]
  reg [31:0] count_4; // @[ivncontrol4.scala 52:20]
  reg [31:0] count_5; // @[ivncontrol4.scala 52:20]
  reg [31:0] count_6; // @[ivncontrol4.scala 52:20]
  reg [31:0] count_7; // @[ivncontrol4.scala 52:20]
  wire [15:0] _GEN_66 = 3'h0 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_0_1 : io_Stationary_matrix_0_0; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_67 = 3'h0 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_0_2 : _GEN_66; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_68 = 3'h0 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_0_3 : _GEN_67; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_69 = 3'h0 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_0_4 : _GEN_68; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_70 = 3'h0 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_0_5 : _GEN_69; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_71 = 3'h0 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_0_6 : _GEN_70; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_72 = 3'h0 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_0_7 : _GEN_71; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_73 = 3'h1 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_1_0 : _GEN_72; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_74 = 3'h1 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_1_1 : _GEN_73; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_75 = 3'h1 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_1_2 : _GEN_74; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_76 = 3'h1 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_1_3 : _GEN_75; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_77 = 3'h1 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_1_4 : _GEN_76; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_78 = 3'h1 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_1_5 : _GEN_77; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_79 = 3'h1 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_1_6 : _GEN_78; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_80 = 3'h1 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_1_7 : _GEN_79; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_81 = 3'h2 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_2_0 : _GEN_80; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_82 = 3'h2 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_2_1 : _GEN_81; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_83 = 3'h2 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_2_2 : _GEN_82; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_84 = 3'h2 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_2_3 : _GEN_83; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_85 = 3'h2 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_2_4 : _GEN_84; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_86 = 3'h2 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_2_5 : _GEN_85; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_87 = 3'h2 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_2_6 : _GEN_86; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_88 = 3'h2 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_2_7 : _GEN_87; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_89 = 3'h3 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_3_0 : _GEN_88; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_90 = 3'h3 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_3_1 : _GEN_89; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_91 = 3'h3 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_3_2 : _GEN_90; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_92 = 3'h3 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_3_3 : _GEN_91; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_93 = 3'h3 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_3_4 : _GEN_92; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_94 = 3'h3 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_3_5 : _GEN_93; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_95 = 3'h3 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_3_6 : _GEN_94; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_96 = 3'h3 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_3_7 : _GEN_95; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_97 = 3'h4 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_4_0 : _GEN_96; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_98 = 3'h4 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_4_1 : _GEN_97; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_99 = 3'h4 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_4_2 : _GEN_98; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_100 = 3'h4 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_4_3 : _GEN_99; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_101 = 3'h4 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_4_4 : _GEN_100; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_102 = 3'h4 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_4_5 : _GEN_101; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_103 = 3'h4 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_4_6 : _GEN_102; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_104 = 3'h4 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_4_7 : _GEN_103; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_105 = 3'h5 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_5_0 : _GEN_104; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_106 = 3'h5 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_5_1 : _GEN_105; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_107 = 3'h5 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_5_2 : _GEN_106; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_108 = 3'h5 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_5_3 : _GEN_107; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_109 = 3'h5 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_5_4 : _GEN_108; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_110 = 3'h5 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_5_5 : _GEN_109; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_111 = 3'h5 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_5_6 : _GEN_110; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_112 = 3'h5 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_5_7 : _GEN_111; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_113 = 3'h6 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_6_0 : _GEN_112; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_114 = 3'h6 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_6_1 : _GEN_113; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_115 = 3'h6 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_6_2 : _GEN_114; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_116 = 3'h6 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_6_3 : _GEN_115; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_117 = 3'h6 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_6_4 : _GEN_116; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_118 = 3'h6 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_6_5 : _GEN_117; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_119 = 3'h6 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_6_6 : _GEN_118; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_120 = 3'h6 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_6_7 : _GEN_119; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_121 = 3'h7 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_7_0 : _GEN_120; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_122 = 3'h7 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_7_1 : _GEN_121; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_123 = 3'h7 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_7_2 : _GEN_122; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_124 = 3'h7 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_7_3 : _GEN_123; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_125 = 3'h7 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_7_4 : _GEN_124; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_126 = 3'h7 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_7_5 : _GEN_125; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_127 = 3'h7 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_7_6 : _GEN_126; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_128 = 3'h7 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_7_7 : _GEN_127; // @[ivncontrol4.scala 57:{15,15}]
  wire [31:0] _mat_T_3_T_4 = {{16'd0}, _GEN_128}; // @[ivncontrol4.scala 57:{15,15}]
  wire  _GEN_225 = count_7 >= 32'h8; // @[ivncontrol4.scala 66:28 67:16]
  wire  valid1 = count_7 >= 32'h8; // @[ivncontrol4.scala 66:28 67:16]
  wire [31:0] _GEN_194 = 3'h1 == i[2:0] ? count_1 : count_0; // @[ivncontrol4.scala 60:{33,33}]
  wire [31:0] _GEN_195 = 3'h2 == i[2:0] ? count_2 : _GEN_194; // @[ivncontrol4.scala 60:{33,33}]
  wire [31:0] _GEN_196 = 3'h3 == i[2:0] ? count_3 : _GEN_195; // @[ivncontrol4.scala 60:{33,33}]
  wire [31:0] _GEN_197 = 3'h4 == i[2:0] ? count_4 : _GEN_196; // @[ivncontrol4.scala 60:{33,33}]
  wire [31:0] _GEN_198 = 3'h5 == i[2:0] ? count_5 : _GEN_197; // @[ivncontrol4.scala 60:{33,33}]
  wire [31:0] _GEN_199 = 3'h6 == i[2:0] ? count_6 : _GEN_198; // @[ivncontrol4.scala 60:{33,33}]
  wire [31:0] _GEN_200 = 3'h7 == i[2:0] ? count_7 : _GEN_199; // @[ivncontrol4.scala 60:{33,33}]
  wire [31:0] _count_T_2 = _GEN_200 + 32'h1; // @[ivncontrol4.scala 60:33]
  wire [31:0] _i_T_1 = i + 32'h1; // @[ivncontrol4.scala 104:16]
  wire [31:0] _j_T_1 = j + 32'h1; // @[ivncontrol4.scala 108:16]
  wire  _GEN_244 = _k_T_2; // @[ivncontrol4.scala 136:75 137:14 139:14]
  wire [31:0] _GEN_245 = rowcount_0 != 32'h0 ? 32'h0 : pin; // @[ivncontrol4.scala 145:30 146:13 31:22]
  wire  _T_27 = rowcount_0 == 32'h0; // @[ivncontrol4.scala 148:23]
  wire [31:0] _GEN_246 = rowcount_0 == 32'h0 & rowcount_1 != 32'h0 ? 32'h1 : _GEN_245; // @[ivncontrol4.scala 148:54 149:13]
  wire  _T_32 = _T_27 & rowcount_1 == 32'h0; // @[ivncontrol4.scala 151:31]
  wire [31:0] _GEN_247 = _T_27 & rowcount_1 == 32'h0 & rowcount_2 != 32'h0 ? 32'h2 : _GEN_246; // @[ivncontrol4.scala 151:77 152:13]
  wire  _T_39 = _T_32 & rowcount_2 == 32'h0; // @[ivncontrol4.scala 154:54]
  wire [31:0] _GEN_248 = _T_32 & rowcount_2 == 32'h0 & rowcount_3 != 32'h0 ? 32'h3 : _GEN_247; // @[ivncontrol4.scala 154:100 155:13]
  wire  _T_48 = _T_39 & rowcount_3 == 32'h0; // @[ivncontrol4.scala 157:77]
  wire [31:0] _GEN_249 = _T_39 & rowcount_3 == 32'h0 & rowcount_4 != 32'h0 ? 32'h4 : _GEN_248; // @[ivncontrol4.scala 157:123 158:13]
  wire  _T_59 = _T_48 & rowcount_4 == 32'h0; // @[ivncontrol4.scala 160:100]
  wire  _T_72 = _T_59 & rowcount_5 == 32'h0; // @[ivncontrol4.scala 163:123]
  wire  valid = _k_T_2; // @[ivncontrol4.scala 136:75 137:14 139:14]
  wire [32:0] _T_91 = {{1'd0}, pin}; // @[ivncontrol4.scala 174:27]
  wire [31:0] _GEN_254 = 4'h1 == _T_91[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_255 = 4'h2 == _T_91[3:0] ? rowcount_2 : _GEN_254; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_256 = 4'h3 == _T_91[3:0] ? rowcount_3 : _GEN_255; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_257 = 4'h4 == _T_91[3:0] ? rowcount_4 : _GEN_256; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_258 = 4'h5 == _T_91[3:0] ? rowcount_5 : _GEN_257; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_259 = 4'h6 == _T_91[3:0] ? rowcount_6 : _GEN_258; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_260 = 4'h7 == _T_91[3:0] ? rowcount_7 : _GEN_259; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_261 = 4'h8 == _T_91[3:0] ? rowcount_8 : _GEN_260; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_262 = 4'h9 == _T_91[3:0] ? rowcount_9 : _GEN_261; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_263 = 4'ha == _T_91[3:0] ? rowcount_10 : _GEN_262; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_264 = 4'hb == _T_91[3:0] ? rowcount_11 : _GEN_263; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_265 = 4'hc == _T_91[3:0] ? rowcount_12 : _GEN_264; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_266 = 4'hd == _T_91[3:0] ? rowcount_13 : _GEN_265; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_267 = 4'he == _T_91[3:0] ? rowcount_14 : _GEN_266; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_268 = 4'hf == _T_91[3:0] ? rowcount_15 : _GEN_267; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_381 = _GEN_268 == 32'h1 ? _T_91[31:0] : 32'h13; // @[ivncontrol4.scala 125:17 224:50 225:21]
  wire [31:0] _GEN_382 = _GEN_268 == 32'h2 ? _T_91[31:0] : _GEN_381; // @[ivncontrol4.scala 220:51 221:21]
  wire [31:0] _GEN_383 = _GEN_268 == 32'h2 ? _T_91[31:0] : 32'h1e; // @[ivncontrol4.scala 125:17 220:51 222:21]
  wire [31:0] _GEN_384 = _GEN_268 == 32'h3 ? _T_91[31:0] : _GEN_382; // @[ivncontrol4.scala 215:50 216:21]
  wire [31:0] _GEN_385 = _GEN_268 == 32'h3 ? _T_91[31:0] : _GEN_383; // @[ivncontrol4.scala 215:50 217:21]
  wire [31:0] _GEN_386 = _GEN_268 == 32'h3 ? _T_91[31:0] : 32'hc; // @[ivncontrol4.scala 125:17 215:50 218:21]
  wire [31:0] _GEN_387 = _GEN_268 == 32'h4 ? _T_91[31:0] : _GEN_384; // @[ivncontrol4.scala 207:50 208:21]
  wire [31:0] _GEN_388 = _GEN_268 == 32'h4 ? _T_91[31:0] : _GEN_385; // @[ivncontrol4.scala 207:50 209:21]
  wire [31:0] _GEN_389 = _GEN_268 == 32'h4 ? _T_91[31:0] : _GEN_386; // @[ivncontrol4.scala 207:50 210:21]
  wire [31:0] _GEN_390 = _GEN_268 == 32'h4 ? _T_91[31:0] : 32'h1d; // @[ivncontrol4.scala 125:17 207:50 211:21]
  wire [31:0] _GEN_391 = _GEN_268 == 32'h5 ? _T_91[31:0] : _GEN_387; // @[ivncontrol4.scala 200:50 201:21]
  wire [31:0] _GEN_392 = _GEN_268 == 32'h5 ? _T_91[31:0] : _GEN_388; // @[ivncontrol4.scala 200:50 202:21]
  wire [31:0] _GEN_393 = _GEN_268 == 32'h5 ? _T_91[31:0] : _GEN_389; // @[ivncontrol4.scala 200:50 203:21]
  wire [31:0] _GEN_394 = _GEN_268 == 32'h5 ? _T_91[31:0] : _GEN_390; // @[ivncontrol4.scala 200:50 204:21]
  wire [31:0] _GEN_395 = _GEN_268 == 32'h5 ? _T_91[31:0] : 32'h12; // @[ivncontrol4.scala 126:18 200:50 205:22]
  wire [31:0] _GEN_396 = _GEN_268 == 32'h6 ? _T_91[31:0] : _GEN_391; // @[ivncontrol4.scala 192:52 193:21]
  wire [31:0] _GEN_397 = _GEN_268 == 32'h6 ? _T_91[31:0] : _GEN_392; // @[ivncontrol4.scala 192:52 194:21]
  wire [31:0] _GEN_398 = _GEN_268 == 32'h6 ? _T_91[31:0] : _GEN_393; // @[ivncontrol4.scala 192:52 195:21]
  wire [31:0] _GEN_399 = _GEN_268 == 32'h6 ? _T_91[31:0] : _GEN_394; // @[ivncontrol4.scala 192:52 196:21]
  wire [31:0] _GEN_400 = _GEN_268 == 32'h6 ? _T_91[31:0] : _GEN_395; // @[ivncontrol4.scala 192:52 197:22]
  wire [31:0] _GEN_401 = _GEN_268 == 32'h6 ? _T_91[31:0] : 32'he; // @[ivncontrol4.scala 126:18 192:52 198:22]
  wire [31:0] _GEN_402 = _GEN_268 == 32'h7 ? _T_91[31:0] : _GEN_396; // @[ivncontrol4.scala 184:52 185:21]
  wire [31:0] _GEN_403 = _GEN_268 == 32'h7 ? _T_91[31:0] : _GEN_397; // @[ivncontrol4.scala 184:52 186:21]
  wire [31:0] _GEN_404 = _GEN_268 == 32'h7 ? _T_91[31:0] : _GEN_398; // @[ivncontrol4.scala 184:52 187:21]
  wire [31:0] _GEN_405 = _GEN_268 == 32'h7 ? _T_91[31:0] : _GEN_399; // @[ivncontrol4.scala 184:52 188:21]
  wire [31:0] _GEN_406 = _GEN_268 == 32'h7 ? _T_91[31:0] : _GEN_400; // @[ivncontrol4.scala 184:52 189:22]
  wire [31:0] _GEN_407 = _GEN_268 == 32'h7 ? _T_91[31:0] : _GEN_401; // @[ivncontrol4.scala 184:52 190:22]
  wire [31:0] _GEN_408 = _GEN_268 == 32'h7 ? _T_91[31:0] : 32'h1f; // @[ivncontrol4.scala 126:18 184:52 191:22]
  wire [31:0] _GEN_409 = _GEN_268 >= 32'h8 ? _T_91[31:0] : _GEN_402; // @[ivncontrol4.scala 174:42 175:21]
  wire [31:0] _GEN_410 = _GEN_268 >= 32'h8 ? _T_91[31:0] : _GEN_403; // @[ivncontrol4.scala 174:42 176:21]
  wire [31:0] _GEN_411 = _GEN_268 >= 32'h8 ? _T_91[31:0] : _GEN_404; // @[ivncontrol4.scala 174:42 177:21]
  wire [31:0] _GEN_412 = _GEN_268 >= 32'h8 ? _T_91[31:0] : _GEN_405; // @[ivncontrol4.scala 174:42 178:21]
  wire [31:0] _GEN_413 = _GEN_268 >= 32'h8 ? _T_91[31:0] : _GEN_406; // @[ivncontrol4.scala 174:42 179:22]
  wire [31:0] _GEN_414 = _GEN_268 >= 32'h8 ? _T_91[31:0] : _GEN_407; // @[ivncontrol4.scala 174:42 180:22]
  wire [31:0] _GEN_415 = _GEN_268 >= 32'h8 ? _T_91[31:0] : _GEN_408; // @[ivncontrol4.scala 174:42 181:22]
  wire [31:0] _GEN_416 = _GEN_268 >= 32'h8 ? _T_91[31:0] : 32'hb; // @[ivncontrol4.scala 126:18 174:42 182:22]
  wire [31:0] _T_127 = 32'h8 - _GEN_268; // @[ivncontrol4.scala 228:18]
  wire [31:0] _i_vn_1_T_15 = 32'h1 + pin; // @[ivncontrol4.scala 229:29]
  wire [31:0] _GEN_529 = _T_127 == 32'h1 ? _i_vn_1_T_15 : _GEN_416; // @[ivncontrol4.scala 269:54 272:22]
  wire [31:0] _GEN_530 = _T_127 == 32'h2 ? _i_vn_1_T_15 : _GEN_415; // @[ivncontrol4.scala 264:54 267:22]
  wire [31:0] _GEN_531 = _T_127 == 32'h2 ? _i_vn_1_T_15 : _GEN_529; // @[ivncontrol4.scala 264:54 268:22]
  wire [31:0] _GEN_532 = _T_127 == 32'h3 ? _i_vn_1_T_15 : _GEN_414; // @[ivncontrol4.scala 257:54 259:22]
  wire [31:0] _GEN_533 = _T_127 == 32'h3 ? _i_vn_1_T_15 : _GEN_530; // @[ivncontrol4.scala 257:54 260:22]
  wire [31:0] _GEN_534 = _T_127 == 32'h3 ? _i_vn_1_T_15 : _GEN_531; // @[ivncontrol4.scala 257:54 261:22]
  wire [31:0] _GEN_535 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_413; // @[ivncontrol4.scala 251:54 253:22]
  wire [31:0] _GEN_536 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_532; // @[ivncontrol4.scala 251:54 254:22]
  wire [31:0] _GEN_537 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_533; // @[ivncontrol4.scala 251:54 255:22]
  wire [31:0] _GEN_538 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_534; // @[ivncontrol4.scala 251:54 256:22]
  wire [31:0] _GEN_539 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_412; // @[ivncontrol4.scala 244:54 246:21]
  wire [31:0] _GEN_540 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_535; // @[ivncontrol4.scala 244:54 247:22]
  wire [31:0] _GEN_541 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_536; // @[ivncontrol4.scala 244:54 248:22]
  wire [31:0] _GEN_542 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_537; // @[ivncontrol4.scala 244:54 249:22]
  wire [31:0] _GEN_543 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_538; // @[ivncontrol4.scala 244:54 250:22]
  wire [31:0] _GEN_544 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_411; // @[ivncontrol4.scala 237:54 238:22]
  wire [31:0] _GEN_545 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_539; // @[ivncontrol4.scala 237:54 239:21]
  wire [31:0] _GEN_546 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_540; // @[ivncontrol4.scala 237:54 240:22]
  wire [31:0] _GEN_547 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_541; // @[ivncontrol4.scala 237:54 241:22]
  wire [31:0] _GEN_548 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_542; // @[ivncontrol4.scala 237:54 242:22]
  wire [31:0] _GEN_549 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_543; // @[ivncontrol4.scala 237:54 243:22]
  wire [31:0] _GEN_550 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_410; // @[ivncontrol4.scala 228:49 229:22]
  wire [31:0] _GEN_551 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_544; // @[ivncontrol4.scala 228:49 230:21]
  wire [31:0] _GEN_552 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_545; // @[ivncontrol4.scala 228:49 231:21]
  wire [31:0] _GEN_553 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_546; // @[ivncontrol4.scala 228:49 232:22]
  wire [31:0] _GEN_554 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_547; // @[ivncontrol4.scala 228:49 233:22]
  wire [31:0] _GEN_555 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_548; // @[ivncontrol4.scala 228:49 234:22]
  wire [31:0] _GEN_556 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_549; // @[ivncontrol4.scala 228:49 235:22]
  wire [31:0] _GEN_574 = 4'h1 == _i_vn_1_T_15[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_575 = 4'h2 == _i_vn_1_T_15[3:0] ? rowcount_2 : _GEN_574; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_576 = 4'h3 == _i_vn_1_T_15[3:0] ? rowcount_3 : _GEN_575; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_577 = 4'h4 == _i_vn_1_T_15[3:0] ? rowcount_4 : _GEN_576; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_578 = 4'h5 == _i_vn_1_T_15[3:0] ? rowcount_5 : _GEN_577; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_579 = 4'h6 == _i_vn_1_T_15[3:0] ? rowcount_6 : _GEN_578; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_580 = 4'h7 == _i_vn_1_T_15[3:0] ? rowcount_7 : _GEN_579; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_581 = 4'h8 == _i_vn_1_T_15[3:0] ? rowcount_8 : _GEN_580; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_582 = 4'h9 == _i_vn_1_T_15[3:0] ? rowcount_9 : _GEN_581; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_583 = 4'ha == _i_vn_1_T_15[3:0] ? rowcount_10 : _GEN_582; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_584 = 4'hb == _i_vn_1_T_15[3:0] ? rowcount_11 : _GEN_583; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_585 = 4'hc == _i_vn_1_T_15[3:0] ? rowcount_12 : _GEN_584; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_586 = 4'hd == _i_vn_1_T_15[3:0] ? rowcount_13 : _GEN_585; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_587 = 4'he == _i_vn_1_T_15[3:0] ? rowcount_14 : _GEN_586; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_588 = 4'hf == _i_vn_1_T_15[3:0] ? rowcount_15 : _GEN_587; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _T_172 = _GEN_268 + _GEN_588; // @[ivncontrol4.scala 275:41]
  wire [31:0] _T_174 = 32'h8 - _T_172; // @[ivncontrol4.scala 275:18]
  wire [31:0] _i_vn_1_T_17 = 32'h2 + pin; // @[ivncontrol4.scala 276:29]
  wire [31:0] _GEN_781 = _T_174 == 32'h1 ? _i_vn_1_T_17 : _GEN_556; // @[ivncontrol4.scala 318:78 321:22]
  wire [31:0] _GEN_782 = _T_174 == 32'h2 ? _i_vn_1_T_17 : _GEN_555; // @[ivncontrol4.scala 312:76 315:22]
  wire [31:0] _GEN_783 = _T_174 == 32'h2 ? _i_vn_1_T_17 : _GEN_781; // @[ivncontrol4.scala 312:76 316:22]
  wire [31:0] _GEN_784 = _T_174 == 32'h3 ? _i_vn_1_T_17 : _GEN_554; // @[ivncontrol4.scala 305:78 307:23]
  wire [31:0] _GEN_785 = _T_174 == 32'h3 ? _i_vn_1_T_17 : _GEN_782; // @[ivncontrol4.scala 305:78 308:22]
  wire [31:0] _GEN_786 = _T_174 == 32'h3 ? _i_vn_1_T_17 : _GEN_783; // @[ivncontrol4.scala 305:78 309:22]
  wire [31:0] _GEN_787 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_553; // @[ivncontrol4.scala 299:78 301:22]
  wire [31:0] _GEN_788 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_784; // @[ivncontrol4.scala 299:78 302:22]
  wire [31:0] _GEN_789 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_785; // @[ivncontrol4.scala 299:78 303:22]
  wire [31:0] _GEN_790 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_786; // @[ivncontrol4.scala 299:78 304:22]
  wire [31:0] _GEN_791 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_552; // @[ivncontrol4.scala 292:76 294:23]
  wire [31:0] _GEN_792 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_787; // @[ivncontrol4.scala 292:76 295:22]
  wire [31:0] _GEN_793 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_788; // @[ivncontrol4.scala 292:76 296:22]
  wire [31:0] _GEN_794 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_789; // @[ivncontrol4.scala 292:76 297:22]
  wire [31:0] _GEN_795 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_790; // @[ivncontrol4.scala 292:76 298:22]
  wire [31:0] _GEN_796 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_551; // @[ivncontrol4.scala 284:77 286:22]
  wire [31:0] _GEN_797 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_791; // @[ivncontrol4.scala 284:77 287:21]
  wire [31:0] _GEN_798 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_792; // @[ivncontrol4.scala 284:77 288:22]
  wire [31:0] _GEN_799 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_793; // @[ivncontrol4.scala 284:77 289:22]
  wire [31:0] _GEN_800 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_794; // @[ivncontrol4.scala 284:77 290:22]
  wire [31:0] _GEN_801 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_795; // @[ivncontrol4.scala 284:77 291:22]
  wire [31:0] _GEN_802 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_550; // @[ivncontrol4.scala 275:73 276:22]
  wire [31:0] _GEN_803 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_796; // @[ivncontrol4.scala 275:73 277:21]
  wire [31:0] _GEN_804 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_797; // @[ivncontrol4.scala 275:73 278:21]
  wire [31:0] _GEN_805 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_798; // @[ivncontrol4.scala 275:73 279:22]
  wire [31:0] _GEN_806 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_799; // @[ivncontrol4.scala 275:73 280:22]
  wire [31:0] _GEN_807 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_800; // @[ivncontrol4.scala 275:73 281:22]
  wire [31:0] _GEN_808 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_801; // @[ivncontrol4.scala 275:73 282:22]
  wire [31:0] _GEN_842 = 4'h1 == _i_vn_1_T_17[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_843 = 4'h2 == _i_vn_1_T_17[3:0] ? rowcount_2 : _GEN_842; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_844 = 4'h3 == _i_vn_1_T_17[3:0] ? rowcount_3 : _GEN_843; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_845 = 4'h4 == _i_vn_1_T_17[3:0] ? rowcount_4 : _GEN_844; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_846 = 4'h5 == _i_vn_1_T_17[3:0] ? rowcount_5 : _GEN_845; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_847 = 4'h6 == _i_vn_1_T_17[3:0] ? rowcount_6 : _GEN_846; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_848 = 4'h7 == _i_vn_1_T_17[3:0] ? rowcount_7 : _GEN_847; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_849 = 4'h8 == _i_vn_1_T_17[3:0] ? rowcount_8 : _GEN_848; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_850 = 4'h9 == _i_vn_1_T_17[3:0] ? rowcount_9 : _GEN_849; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_851 = 4'ha == _i_vn_1_T_17[3:0] ? rowcount_10 : _GEN_850; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_852 = 4'hb == _i_vn_1_T_17[3:0] ? rowcount_11 : _GEN_851; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_853 = 4'hc == _i_vn_1_T_17[3:0] ? rowcount_12 : _GEN_852; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_854 = 4'hd == _i_vn_1_T_17[3:0] ? rowcount_13 : _GEN_853; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_855 = 4'he == _i_vn_1_T_17[3:0] ? rowcount_14 : _GEN_854; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_856 = 4'hf == _i_vn_1_T_17[3:0] ? rowcount_15 : _GEN_855; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _T_254 = _T_172 + _GEN_856; // @[ivncontrol4.scala 326:62]
  wire [31:0] _T_256 = 32'h8 - _T_254; // @[ivncontrol4.scala 326:17]
  wire [31:0] _i_vn_1_T_19 = 32'h3 + pin; // @[ivncontrol4.scala 327:29]
  wire [31:0] _GEN_1145 = _T_256 == 32'h1 ? _i_vn_1_T_19 : _GEN_808; // @[ivncontrol4.scala 369:100 372:22]
  wire [31:0] _GEN_1146 = _T_256 == 32'h2 ? _i_vn_1_T_19 : _GEN_807; // @[ivncontrol4.scala 363:98 366:22]
  wire [31:0] _GEN_1147 = _T_256 == 32'h2 ? _i_vn_1_T_19 : _GEN_1145; // @[ivncontrol4.scala 363:98 367:22]
  wire [31:0] _GEN_1148 = _T_256 == 32'h3 ? _i_vn_1_T_19 : _GEN_806; // @[ivncontrol4.scala 356:100 358:23]
  wire [31:0] _GEN_1149 = _T_256 == 32'h3 ? _i_vn_1_T_19 : _GEN_1146; // @[ivncontrol4.scala 356:100 359:22]
  wire [31:0] _GEN_1150 = _T_256 == 32'h3 ? _i_vn_1_T_19 : _GEN_1147; // @[ivncontrol4.scala 356:100 360:22]
  wire [31:0] _GEN_1151 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_805; // @[ivncontrol4.scala 350:100 352:22]
  wire [31:0] _GEN_1152 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_1148; // @[ivncontrol4.scala 350:100 353:22]
  wire [31:0] _GEN_1153 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_1149; // @[ivncontrol4.scala 350:100 354:22]
  wire [31:0] _GEN_1154 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_1150; // @[ivncontrol4.scala 350:100 355:22]
  wire [31:0] _GEN_1155 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_804; // @[ivncontrol4.scala 343:98 345:23]
  wire [31:0] _GEN_1156 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1151; // @[ivncontrol4.scala 343:98 346:22]
  wire [31:0] _GEN_1157 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1152; // @[ivncontrol4.scala 343:98 347:22]
  wire [31:0] _GEN_1158 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1153; // @[ivncontrol4.scala 343:98 348:22]
  wire [31:0] _GEN_1159 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1154; // @[ivncontrol4.scala 343:98 349:22]
  wire [31:0] _GEN_1160 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_803; // @[ivncontrol4.scala 335:99 337:22]
  wire [31:0] _GEN_1161 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1155; // @[ivncontrol4.scala 335:99 338:21]
  wire [31:0] _GEN_1162 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1156; // @[ivncontrol4.scala 335:99 339:22]
  wire [31:0] _GEN_1163 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1157; // @[ivncontrol4.scala 335:99 340:22]
  wire [31:0] _GEN_1164 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1158; // @[ivncontrol4.scala 335:99 341:22]
  wire [31:0] _GEN_1165 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1159; // @[ivncontrol4.scala 335:99 342:22]
  wire [31:0] _GEN_1166 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_802; // @[ivncontrol4.scala 326:94 327:22]
  wire [31:0] _GEN_1167 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1160; // @[ivncontrol4.scala 326:94 328:21]
  wire [31:0] _GEN_1168 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1161; // @[ivncontrol4.scala 326:94 329:21]
  wire [31:0] _GEN_1169 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1162; // @[ivncontrol4.scala 326:94 330:22]
  wire [31:0] _GEN_1170 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1163; // @[ivncontrol4.scala 326:94 331:22]
  wire [31:0] _GEN_1171 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1164; // @[ivncontrol4.scala 326:94 332:22]
  wire [31:0] _GEN_1172 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1165; // @[ivncontrol4.scala 326:94 333:22]
  wire [31:0] _GEN_1222 = 4'h1 == _i_vn_1_T_19[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1223 = 4'h2 == _i_vn_1_T_19[3:0] ? rowcount_2 : _GEN_1222; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1224 = 4'h3 == _i_vn_1_T_19[3:0] ? rowcount_3 : _GEN_1223; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1225 = 4'h4 == _i_vn_1_T_19[3:0] ? rowcount_4 : _GEN_1224; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1226 = 4'h5 == _i_vn_1_T_19[3:0] ? rowcount_5 : _GEN_1225; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1227 = 4'h6 == _i_vn_1_T_19[3:0] ? rowcount_6 : _GEN_1226; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1228 = 4'h7 == _i_vn_1_T_19[3:0] ? rowcount_7 : _GEN_1227; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1229 = 4'h8 == _i_vn_1_T_19[3:0] ? rowcount_8 : _GEN_1228; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1230 = 4'h9 == _i_vn_1_T_19[3:0] ? rowcount_9 : _GEN_1229; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1231 = 4'ha == _i_vn_1_T_19[3:0] ? rowcount_10 : _GEN_1230; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1232 = 4'hb == _i_vn_1_T_19[3:0] ? rowcount_11 : _GEN_1231; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1233 = 4'hc == _i_vn_1_T_19[3:0] ? rowcount_12 : _GEN_1232; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1234 = 4'hd == _i_vn_1_T_19[3:0] ? rowcount_13 : _GEN_1233; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1235 = 4'he == _i_vn_1_T_19[3:0] ? rowcount_14 : _GEN_1234; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1236 = 4'hf == _i_vn_1_T_19[3:0] ? rowcount_15 : _GEN_1235; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _T_371 = _T_254 + _GEN_1236; // @[ivncontrol4.scala 376:86]
  wire [31:0] _T_373 = 32'h8 - _T_371; // @[ivncontrol4.scala 376:19]
  wire [31:0] _i_vn_1_T_21 = 32'h4 + pin; // @[ivncontrol4.scala 377:29]
  wire [31:0] _GEN_1621 = _T_373 == 32'h1 ? _i_vn_1_T_21 : _GEN_1172; // @[ivncontrol4.scala 419:122 422:22]
  wire [31:0] _GEN_1622 = _T_373 == 32'h2 ? _i_vn_1_T_21 : _GEN_1171; // @[ivncontrol4.scala 413:121 416:22]
  wire [31:0] _GEN_1623 = _T_373 == 32'h2 ? _i_vn_1_T_21 : _GEN_1621; // @[ivncontrol4.scala 413:121 417:22]
  wire [31:0] _GEN_1624 = _T_373 == 32'h3 ? _i_vn_1_T_21 : _GEN_1170; // @[ivncontrol4.scala 406:123 408:23]
  wire [31:0] _GEN_1625 = _T_373 == 32'h3 ? _i_vn_1_T_21 : _GEN_1622; // @[ivncontrol4.scala 406:123 409:22]
  wire [31:0] _GEN_1626 = _T_373 == 32'h3 ? _i_vn_1_T_21 : _GEN_1623; // @[ivncontrol4.scala 406:123 410:22]
  wire [31:0] _GEN_1627 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1169; // @[ivncontrol4.scala 400:122 402:22]
  wire [31:0] _GEN_1628 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1624; // @[ivncontrol4.scala 400:122 403:22]
  wire [31:0] _GEN_1629 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1625; // @[ivncontrol4.scala 400:122 404:22]
  wire [31:0] _GEN_1630 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1626; // @[ivncontrol4.scala 400:122 405:22]
  wire [31:0] _GEN_1631 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1168; // @[ivncontrol4.scala 393:121 395:23]
  wire [31:0] _GEN_1632 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1627; // @[ivncontrol4.scala 393:121 396:22]
  wire [31:0] _GEN_1633 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1628; // @[ivncontrol4.scala 393:121 397:22]
  wire [31:0] _GEN_1634 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1629; // @[ivncontrol4.scala 393:121 398:22]
  wire [31:0] _GEN_1635 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1630; // @[ivncontrol4.scala 393:121 399:22]
  wire [31:0] _GEN_1636 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1167; // @[ivncontrol4.scala 385:121 387:22]
  wire [31:0] _GEN_1637 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1631; // @[ivncontrol4.scala 385:121 388:21]
  wire [31:0] _GEN_1638 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1632; // @[ivncontrol4.scala 385:121 389:22]
  wire [31:0] _GEN_1639 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1633; // @[ivncontrol4.scala 385:121 390:22]
  wire [31:0] _GEN_1640 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1634; // @[ivncontrol4.scala 385:121 391:22]
  wire [31:0] _GEN_1641 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1635; // @[ivncontrol4.scala 385:121 392:22]
  wire [31:0] _GEN_1642 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1166; // @[ivncontrol4.scala 376:118 377:22]
  wire [31:0] _GEN_1643 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1636; // @[ivncontrol4.scala 376:118 378:21]
  wire [31:0] _GEN_1644 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1637; // @[ivncontrol4.scala 376:118 379:21]
  wire [31:0] _GEN_1645 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1638; // @[ivncontrol4.scala 376:118 380:22]
  wire [31:0] _GEN_1646 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1639; // @[ivncontrol4.scala 376:118 381:22]
  wire [31:0] _GEN_1647 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1640; // @[ivncontrol4.scala 376:118 382:22]
  wire [31:0] _GEN_1648 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1641; // @[ivncontrol4.scala 376:118 383:22]
  wire [31:0] _GEN_1714 = 4'h1 == _i_vn_1_T_21[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1715 = 4'h2 == _i_vn_1_T_21[3:0] ? rowcount_2 : _GEN_1714; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1716 = 4'h3 == _i_vn_1_T_21[3:0] ? rowcount_3 : _GEN_1715; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1717 = 4'h4 == _i_vn_1_T_21[3:0] ? rowcount_4 : _GEN_1716; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1718 = 4'h5 == _i_vn_1_T_21[3:0] ? rowcount_5 : _GEN_1717; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1719 = 4'h6 == _i_vn_1_T_21[3:0] ? rowcount_6 : _GEN_1718; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1720 = 4'h7 == _i_vn_1_T_21[3:0] ? rowcount_7 : _GEN_1719; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1721 = 4'h8 == _i_vn_1_T_21[3:0] ? rowcount_8 : _GEN_1720; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1722 = 4'h9 == _i_vn_1_T_21[3:0] ? rowcount_9 : _GEN_1721; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1723 = 4'ha == _i_vn_1_T_21[3:0] ? rowcount_10 : _GEN_1722; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1724 = 4'hb == _i_vn_1_T_21[3:0] ? rowcount_11 : _GEN_1723; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1725 = 4'hc == _i_vn_1_T_21[3:0] ? rowcount_12 : _GEN_1724; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1726 = 4'hd == _i_vn_1_T_21[3:0] ? rowcount_13 : _GEN_1725; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1727 = 4'he == _i_vn_1_T_21[3:0] ? rowcount_14 : _GEN_1726; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1728 = 4'hf == _i_vn_1_T_21[3:0] ? rowcount_15 : _GEN_1727; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _T_523 = _T_371 + _GEN_1728; // @[ivncontrol4.scala 426:108]
  wire [31:0] _T_525 = 32'h8 - _T_523; // @[ivncontrol4.scala 426:19]
  wire [31:0] _i_vn_1_T_23 = 32'h5 + pin; // @[ivncontrol4.scala 427:29]
  wire [31:0] _GEN_2209 = _T_525 == 32'h1 ? _i_vn_1_T_23 : _GEN_1648; // @[ivncontrol4.scala 469:144 472:22]
  wire [31:0] _GEN_2210 = _T_525 == 32'h2 ? _i_vn_1_T_23 : _GEN_1647; // @[ivncontrol4.scala 463:143 466:22]
  wire [31:0] _GEN_2211 = _T_525 == 32'h2 ? _i_vn_1_T_23 : _GEN_2209; // @[ivncontrol4.scala 463:143 467:22]
  wire [31:0] _GEN_2212 = _T_525 == 32'h3 ? _i_vn_1_T_23 : _GEN_1646; // @[ivncontrol4.scala 456:145 458:23]
  wire [31:0] _GEN_2213 = _T_525 == 32'h3 ? _i_vn_1_T_23 : _GEN_2210; // @[ivncontrol4.scala 456:145 459:22]
  wire [31:0] _GEN_2214 = _T_525 == 32'h3 ? _i_vn_1_T_23 : _GEN_2211; // @[ivncontrol4.scala 456:145 460:22]
  wire [31:0] _GEN_2215 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_1645; // @[ivncontrol4.scala 450:143 452:22]
  wire [31:0] _GEN_2216 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_2212; // @[ivncontrol4.scala 450:143 453:22]
  wire [31:0] _GEN_2217 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_2213; // @[ivncontrol4.scala 450:143 454:22]
  wire [31:0] _GEN_2218 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_2214; // @[ivncontrol4.scala 450:143 455:22]
  wire [31:0] _GEN_2219 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_1644; // @[ivncontrol4.scala 443:143 445:23]
  wire [31:0] _GEN_2220 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2215; // @[ivncontrol4.scala 443:143 446:22]
  wire [31:0] _GEN_2221 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2216; // @[ivncontrol4.scala 443:143 447:22]
  wire [31:0] _GEN_2222 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2217; // @[ivncontrol4.scala 443:143 448:22]
  wire [31:0] _GEN_2223 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2218; // @[ivncontrol4.scala 443:143 449:22]
  wire [31:0] _GEN_2224 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_1643; // @[ivncontrol4.scala 435:143 437:22]
  wire [31:0] _GEN_2225 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2219; // @[ivncontrol4.scala 435:143 438:21]
  wire [31:0] _GEN_2226 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2220; // @[ivncontrol4.scala 435:143 439:22]
  wire [31:0] _GEN_2227 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2221; // @[ivncontrol4.scala 435:143 440:22]
  wire [31:0] _GEN_2228 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2222; // @[ivncontrol4.scala 435:143 441:22]
  wire [31:0] _GEN_2229 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2223; // @[ivncontrol4.scala 435:143 442:22]
  wire [31:0] _GEN_2230 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_1642; // @[ivncontrol4.scala 426:140 427:22]
  wire [31:0] _GEN_2231 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2224; // @[ivncontrol4.scala 426:140 428:21]
  wire [31:0] _GEN_2232 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2225; // @[ivncontrol4.scala 426:140 429:21]
  wire [31:0] _GEN_2233 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2226; // @[ivncontrol4.scala 426:140 430:22]
  wire [31:0] _GEN_2234 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2227; // @[ivncontrol4.scala 426:140 431:22]
  wire [31:0] _GEN_2235 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2228; // @[ivncontrol4.scala 426:140 432:22]
  wire [31:0] _GEN_2236 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2229; // @[ivncontrol4.scala 426:140 433:22]
  wire [31:0] _GEN_2318 = 4'h1 == _i_vn_1_T_23[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2319 = 4'h2 == _i_vn_1_T_23[3:0] ? rowcount_2 : _GEN_2318; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2320 = 4'h3 == _i_vn_1_T_23[3:0] ? rowcount_3 : _GEN_2319; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2321 = 4'h4 == _i_vn_1_T_23[3:0] ? rowcount_4 : _GEN_2320; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2322 = 4'h5 == _i_vn_1_T_23[3:0] ? rowcount_5 : _GEN_2321; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2323 = 4'h6 == _i_vn_1_T_23[3:0] ? rowcount_6 : _GEN_2322; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2324 = 4'h7 == _i_vn_1_T_23[3:0] ? rowcount_7 : _GEN_2323; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2325 = 4'h8 == _i_vn_1_T_23[3:0] ? rowcount_8 : _GEN_2324; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2326 = 4'h9 == _i_vn_1_T_23[3:0] ? rowcount_9 : _GEN_2325; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2327 = 4'ha == _i_vn_1_T_23[3:0] ? rowcount_10 : _GEN_2326; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2328 = 4'hb == _i_vn_1_T_23[3:0] ? rowcount_11 : _GEN_2327; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2329 = 4'hc == _i_vn_1_T_23[3:0] ? rowcount_12 : _GEN_2328; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2330 = 4'hd == _i_vn_1_T_23[3:0] ? rowcount_13 : _GEN_2329; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2331 = 4'he == _i_vn_1_T_23[3:0] ? rowcount_14 : _GEN_2330; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2332 = 4'hf == _i_vn_1_T_23[3:0] ? rowcount_15 : _GEN_2331; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _T_710 = _T_523 + _GEN_2332; // @[ivncontrol4.scala 477:130]
  wire [31:0] _T_712 = 32'h8 - _T_710; // @[ivncontrol4.scala 477:19]
  wire [31:0] _i_vn_1_T_25 = 32'h6 + pin; // @[ivncontrol4.scala 478:29]
  wire [31:0] _GEN_2909 = _T_712 == 32'h1 ? _i_vn_1_T_25 : _GEN_2236; // @[ivncontrol4.scala 520:166 523:22]
  wire [31:0] _GEN_2910 = _T_712 == 32'h2 ? _i_vn_1_T_25 : _GEN_2235; // @[ivncontrol4.scala 514:166 517:22]
  wire [31:0] _GEN_2911 = _T_712 == 32'h2 ? _i_vn_1_T_25 : _GEN_2909; // @[ivncontrol4.scala 514:166 518:22]
  wire [31:0] _GEN_2912 = _T_712 == 32'h3 ? _i_vn_1_T_25 : _GEN_2234; // @[ivncontrol4.scala 507:168 509:23]
  wire [31:0] _GEN_2913 = _T_712 == 32'h3 ? _i_vn_1_T_25 : _GEN_2910; // @[ivncontrol4.scala 507:168 510:22]
  wire [31:0] _GEN_2914 = _T_712 == 32'h3 ? _i_vn_1_T_25 : _GEN_2911; // @[ivncontrol4.scala 507:168 511:22]
  wire [31:0] _GEN_2915 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2233; // @[ivncontrol4.scala 501:166 503:22]
  wire [31:0] _GEN_2916 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2912; // @[ivncontrol4.scala 501:166 504:22]
  wire [31:0] _GEN_2917 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2913; // @[ivncontrol4.scala 501:166 505:22]
  wire [31:0] _GEN_2918 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2914; // @[ivncontrol4.scala 501:166 506:22]
  wire [31:0] _GEN_2919 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2232; // @[ivncontrol4.scala 494:166 496:23]
  wire [31:0] _GEN_2920 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2915; // @[ivncontrol4.scala 494:166 497:22]
  wire [31:0] _GEN_2921 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2916; // @[ivncontrol4.scala 494:166 498:22]
  wire [31:0] _GEN_2922 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2917; // @[ivncontrol4.scala 494:166 499:22]
  wire [31:0] _GEN_2923 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2918; // @[ivncontrol4.scala 494:166 500:22]
  wire [31:0] _GEN_2924 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2231; // @[ivncontrol4.scala 486:166 488:22]
  wire [31:0] _GEN_2925 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2919; // @[ivncontrol4.scala 486:166 489:21]
  wire [31:0] _GEN_2926 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2920; // @[ivncontrol4.scala 486:166 490:22]
  wire [31:0] _GEN_2927 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2921; // @[ivncontrol4.scala 486:166 491:22]
  wire [31:0] _GEN_2928 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2922; // @[ivncontrol4.scala 486:166 492:22]
  wire [31:0] _GEN_2929 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2923; // @[ivncontrol4.scala 486:166 493:22]
  wire [31:0] _GEN_2930 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2230; // @[ivncontrol4.scala 477:162 478:22]
  wire [31:0] _GEN_2931 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2924; // @[ivncontrol4.scala 477:162 479:21]
  wire [31:0] _GEN_2932 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2925; // @[ivncontrol4.scala 477:162 480:21]
  wire [31:0] _GEN_2933 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2926; // @[ivncontrol4.scala 477:162 481:22]
  wire [31:0] _GEN_2934 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2927; // @[ivncontrol4.scala 477:162 482:22]
  wire [31:0] _GEN_2935 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2928; // @[ivncontrol4.scala 477:162 483:22]
  wire [31:0] _GEN_2936 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2929; // @[ivncontrol4.scala 477:162 484:22]
  wire [31:0] _GEN_3034 = 4'h1 == _i_vn_1_T_25[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3035 = 4'h2 == _i_vn_1_T_25[3:0] ? rowcount_2 : _GEN_3034; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3036 = 4'h3 == _i_vn_1_T_25[3:0] ? rowcount_3 : _GEN_3035; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3037 = 4'h4 == _i_vn_1_T_25[3:0] ? rowcount_4 : _GEN_3036; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3038 = 4'h5 == _i_vn_1_T_25[3:0] ? rowcount_5 : _GEN_3037; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3039 = 4'h6 == _i_vn_1_T_25[3:0] ? rowcount_6 : _GEN_3038; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3040 = 4'h7 == _i_vn_1_T_25[3:0] ? rowcount_7 : _GEN_3039; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3041 = 4'h8 == _i_vn_1_T_25[3:0] ? rowcount_8 : _GEN_3040; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3042 = 4'h9 == _i_vn_1_T_25[3:0] ? rowcount_9 : _GEN_3041; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3043 = 4'ha == _i_vn_1_T_25[3:0] ? rowcount_10 : _GEN_3042; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3044 = 4'hb == _i_vn_1_T_25[3:0] ? rowcount_11 : _GEN_3043; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3045 = 4'hc == _i_vn_1_T_25[3:0] ? rowcount_12 : _GEN_3044; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3046 = 4'hd == _i_vn_1_T_25[3:0] ? rowcount_13 : _GEN_3045; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3047 = 4'he == _i_vn_1_T_25[3:0] ? rowcount_14 : _GEN_3046; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3048 = 4'hf == _i_vn_1_T_25[3:0] ? rowcount_15 : _GEN_3047; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _T_932 = _T_710 + _GEN_3048; // @[ivncontrol4.scala 528:152]
  wire [31:0] _T_934 = 32'h8 - _T_932; // @[ivncontrol4.scala 528:19]
  wire [31:0] _i_vn_1_T_27 = 32'h7 + pin; // @[ivncontrol4.scala 529:29]
  wire [31:0] _GEN_3721 = _T_934 == 32'h1 ? _i_vn_1_T_27 : _GEN_2936; // @[ivncontrol4.scala 571:188 574:22]
  wire [31:0] _GEN_3722 = _T_934 == 32'h2 ? _i_vn_1_T_27 : _GEN_2935; // @[ivncontrol4.scala 565:188 568:22]
  wire [31:0] _GEN_3723 = _T_934 == 32'h2 ? _i_vn_1_T_27 : _GEN_3721; // @[ivncontrol4.scala 565:188 569:22]
  wire [31:0] _GEN_3724 = _T_934 == 32'h3 ? _i_vn_1_T_27 : _GEN_2934; // @[ivncontrol4.scala 558:190 560:23]
  wire [31:0] _GEN_3725 = _T_934 == 32'h3 ? _i_vn_1_T_27 : _GEN_3722; // @[ivncontrol4.scala 558:190 561:22]
  wire [31:0] _GEN_3726 = _T_934 == 32'h3 ? _i_vn_1_T_27 : _GEN_3723; // @[ivncontrol4.scala 558:190 562:22]
  wire [31:0] _GEN_3727 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_2933; // @[ivncontrol4.scala 552:188 554:22]
  wire [31:0] _GEN_3728 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_3724; // @[ivncontrol4.scala 552:188 555:22]
  wire [31:0] _GEN_3729 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_3725; // @[ivncontrol4.scala 552:188 556:22]
  wire [31:0] _GEN_3730 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_3726; // @[ivncontrol4.scala 552:188 557:22]
  wire [31:0] _GEN_3731 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_2932; // @[ivncontrol4.scala 545:188 547:23]
  wire [31:0] _GEN_3732 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3727; // @[ivncontrol4.scala 545:188 548:22]
  wire [31:0] _GEN_3733 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3728; // @[ivncontrol4.scala 545:188 549:22]
  wire [31:0] _GEN_3734 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3729; // @[ivncontrol4.scala 545:188 550:22]
  wire [31:0] _GEN_3735 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3730; // @[ivncontrol4.scala 545:188 551:22]
  wire [31:0] _GEN_3736 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_2931; // @[ivncontrol4.scala 537:188 539:22]
  wire [31:0] _GEN_3737 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3731; // @[ivncontrol4.scala 537:188 540:21]
  wire [31:0] _GEN_3738 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3732; // @[ivncontrol4.scala 537:188 541:22]
  wire [31:0] _GEN_3739 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3733; // @[ivncontrol4.scala 537:188 542:22]
  wire [31:0] _GEN_3740 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3734; // @[ivncontrol4.scala 537:188 543:22]
  wire [31:0] _GEN_3741 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3735; // @[ivncontrol4.scala 537:188 544:22]
  wire [31:0] _GEN_3742 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_2930; // @[ivncontrol4.scala 528:184 529:22]
  wire [31:0] _GEN_3743 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3736; // @[ivncontrol4.scala 528:184 530:21]
  wire [31:0] _GEN_3744 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3737; // @[ivncontrol4.scala 528:184 531:21]
  wire [31:0] _GEN_3745 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3738; // @[ivncontrol4.scala 528:184 532:22]
  wire [31:0] _GEN_3746 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3739; // @[ivncontrol4.scala 528:184 533:22]
  wire [31:0] _GEN_3747 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3740; // @[ivncontrol4.scala 528:184 534:22]
  wire [31:0] _GEN_3748 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3741; // @[ivncontrol4.scala 528:184 535:22]
  wire [31:0] _GEN_3749 = _GEN_244 ? _GEN_409 : 32'h13; // @[ivncontrol4.scala 125:17 172:28]
  wire [31:0] _GEN_3750 = _GEN_244 ? _GEN_3742 : 32'h1e; // @[ivncontrol4.scala 125:17 172:28]
  wire [31:0] _GEN_3751 = _GEN_244 ? _GEN_3743 : 32'hc; // @[ivncontrol4.scala 125:17 172:28]
  wire [31:0] _GEN_3752 = _GEN_244 ? _GEN_3744 : 32'h1d; // @[ivncontrol4.scala 125:17 172:28]
  wire [31:0] _GEN_3753 = _GEN_244 ? _GEN_3745 : 32'h12; // @[ivncontrol4.scala 126:18 172:28]
  wire [31:0] _GEN_3754 = _GEN_244 ? _GEN_3746 : 32'he; // @[ivncontrol4.scala 126:18 172:28]
  wire [31:0] _GEN_3755 = _GEN_244 ? _GEN_3747 : 32'h1f; // @[ivncontrol4.scala 126:18 172:28]
  wire [31:0] _GEN_3756 = _GEN_244 ? _GEN_3748 : 32'hb; // @[ivncontrol4.scala 126:18 172:28]
  wire [31:0] _GEN_4137 = reset ? 32'h0 : _GEN_3749; // @[ivncontrol4.scala 16:{23,23}]
  wire [31:0] _GEN_4138 = reset ? 32'h0 : _GEN_3750; // @[ivncontrol4.scala 16:{23,23}]
  wire [31:0] _GEN_4139 = reset ? 32'h0 : _GEN_3751; // @[ivncontrol4.scala 16:{23,23}]
  wire [31:0] _GEN_4140 = reset ? 32'h0 : _GEN_3752; // @[ivncontrol4.scala 16:{23,23}]
  wire [31:0] _GEN_4141 = reset ? 32'h0 : _GEN_3753; // @[ivncontrol4.scala 17:{24,24}]
  wire [31:0] _GEN_4142 = reset ? 32'h0 : _GEN_3754; // @[ivncontrol4.scala 17:{24,24}]
  wire [31:0] _GEN_4143 = reset ? 32'h0 : _GEN_3755; // @[ivncontrol4.scala 17:{24,24}]
  wire [31:0] _GEN_4144 = reset ? 32'h0 : _GEN_3756; // @[ivncontrol4.scala 17:{24,24}]
  assign io_o_vn_0 = i_vn_0; // @[ivncontrol4.scala 121:13]
  assign io_o_vn_1 = i_vn_1; // @[ivncontrol4.scala 121:13]
  assign io_o_vn_2 = i_vn_2; // @[ivncontrol4.scala 121:13]
  assign io_o_vn_3 = i_vn_3; // @[ivncontrol4.scala 121:13]
  assign io_o_vn2_0 = i_vn2_0; // @[ivncontrol4.scala 122:14]
  assign io_o_vn2_1 = i_vn2_1; // @[ivncontrol4.scala 122:14]
  assign io_o_vn2_2 = i_vn2_2; // @[ivncontrol4.scala 122:14]
  assign io_o_vn2_3 = i_vn2_3; // @[ivncontrol4.scala 122:14]
  always @(posedge clock) begin
    i_vn_0 <= _GEN_4137[4:0]; // @[ivncontrol4.scala 16:{23,23}]
    i_vn_1 <= _GEN_4138[4:0]; // @[ivncontrol4.scala 16:{23,23}]
    i_vn_2 <= _GEN_4139[4:0]; // @[ivncontrol4.scala 16:{23,23}]
    i_vn_3 <= _GEN_4140[4:0]; // @[ivncontrol4.scala 16:{23,23}]
    i_vn2_0 <= _GEN_4141[4:0]; // @[ivncontrol4.scala 17:{24,24}]
    i_vn2_1 <= _GEN_4142[4:0]; // @[ivncontrol4.scala 17:{24,24}]
    i_vn2_2 <= _GEN_4143[4:0]; // @[ivncontrol4.scala 17:{24,24}]
    i_vn2_3 <= _GEN_4144[4:0]; // @[ivncontrol4.scala 17:{24,24}]
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_0 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_0 <= count_0; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_1 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_1 <= count_1; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_2 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_2 <= count_2; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_3 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_3 <= count_3; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_4 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_4 <= count_4; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_5 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_5 <= count_5; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_6 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_6 <= count_6; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_7 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_7 <= count_7; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_8 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_8 <= 32'h0; // @[ivncontrol4.scala 81:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_9 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_9 <= 32'h0; // @[ivncontrol4.scala 81:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_10 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_10 <= 32'h0; // @[ivncontrol4.scala 81:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_11 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_11 <= 32'h0; // @[ivncontrol4.scala 81:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_12 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_12 <= 32'h0; // @[ivncontrol4.scala 81:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_13 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_13 <= 32'h0; // @[ivncontrol4.scala 81:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_14 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_14 <= 32'h0; // @[ivncontrol4.scala 81:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_15 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end
    if (reset) begin // @[ivncontrol4.scala 31:22]
      pin <= 32'h0; // @[ivncontrol4.scala 31:22]
    end else if (_T_72 & rowcount_6 == 32'h0 & rowcount_7 != 32'h0) begin // @[ivncontrol4.scala 166:192]
      pin <= 32'h7; // @[ivncontrol4.scala 167:13]
    end else if (_T_59 & rowcount_5 == 32'h0 & rowcount_6 != 32'h0) begin // @[ivncontrol4.scala 163:169]
      pin <= 32'h6; // @[ivncontrol4.scala 164:13]
    end else if (_T_48 & rowcount_4 == 32'h0 & rowcount_5 != 32'h0) begin // @[ivncontrol4.scala 160:146]
      pin <= 32'h5; // @[ivncontrol4.scala 161:13]
    end else begin
      pin <= _GEN_249;
    end
    if (reset) begin // @[ivncontrol4.scala 35:20]
      i <= 32'h0; // @[ivncontrol4.scala 35:20]
    end else if (i < 32'h7 & _k_T_1) begin // @[ivncontrol4.scala 103:74]
      i <= _i_T_1; // @[ivncontrol4.scala 104:11]
    end
    if (reset) begin // @[ivncontrol4.scala 36:20]
      j <= 32'h0; // @[ivncontrol4.scala 36:20]
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 107:71]
      j <= _j_T_1; // @[ivncontrol4.scala 108:11]
    end else if (!(_k_T_2)) begin // @[ivncontrol4.scala 110:81]
      j <= 32'h0; // @[ivncontrol4.scala 114:11]
    end
    if (3'h0 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h0 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h0 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h0 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h0 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h0 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h0 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h0 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h0 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_0 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h1 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_1 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h2 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_2 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h3 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_3 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h4 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_4 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h5 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_5 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h6 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_6 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h7 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_7 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  i_vn_0 = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  i_vn_1 = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  i_vn_2 = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  i_vn_3 = _RAND_3[4:0];
  _RAND_4 = {1{`RANDOM}};
  i_vn2_0 = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  i_vn2_1 = _RAND_5[4:0];
  _RAND_6 = {1{`RANDOM}};
  i_vn2_2 = _RAND_6[4:0];
  _RAND_7 = {1{`RANDOM}};
  i_vn2_3 = _RAND_7[4:0];
  _RAND_8 = {1{`RANDOM}};
  rowcount_0 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  rowcount_1 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  rowcount_2 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  rowcount_3 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  rowcount_4 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  rowcount_5 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  rowcount_6 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  rowcount_7 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  rowcount_8 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  rowcount_9 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  rowcount_10 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  rowcount_11 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  rowcount_12 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  rowcount_13 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  rowcount_14 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  rowcount_15 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  pin = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  i = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  j = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  mat_0_0 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  mat_0_1 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  mat_0_2 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  mat_0_3 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  mat_0_4 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  mat_0_5 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  mat_0_6 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  mat_0_7 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  mat_1_0 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  mat_1_1 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  mat_1_2 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  mat_1_3 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  mat_1_4 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  mat_1_5 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  mat_1_6 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  mat_1_7 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  mat_2_0 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  mat_2_1 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  mat_2_2 = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  mat_2_3 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  mat_2_4 = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  mat_2_5 = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  mat_2_6 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  mat_2_7 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  mat_3_0 = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  mat_3_1 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  mat_3_2 = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  mat_3_3 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  mat_3_4 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  mat_3_5 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  mat_3_6 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  mat_3_7 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  mat_4_0 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  mat_4_1 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  mat_4_2 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  mat_4_3 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  mat_4_4 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  mat_4_5 = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  mat_4_6 = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  mat_4_7 = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  mat_5_0 = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  mat_5_1 = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  mat_5_2 = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  mat_5_3 = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  mat_5_4 = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  mat_5_5 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  mat_5_6 = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  mat_5_7 = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  mat_6_0 = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  mat_6_1 = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  mat_6_2 = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  mat_6_3 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  mat_6_4 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  mat_6_5 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  mat_6_6 = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  mat_6_7 = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  mat_7_0 = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  mat_7_1 = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  mat_7_2 = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  mat_7_3 = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  mat_7_4 = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  mat_7_5 = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  mat_7_6 = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  mat_7_7 = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  count_0 = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  count_1 = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  count_2 = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  count_3 = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  count_4 = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  count_5 = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  count_6 = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  count_7 = _RAND_98[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ivncontrol4_6(
  input         clock,
  input         reset,
  input  [15:0] io_Stationary_matrix_0_0,
  input  [15:0] io_Stationary_matrix_0_1,
  input  [15:0] io_Stationary_matrix_0_2,
  input  [15:0] io_Stationary_matrix_0_3,
  input  [15:0] io_Stationary_matrix_0_4,
  input  [15:0] io_Stationary_matrix_0_5,
  input  [15:0] io_Stationary_matrix_0_6,
  input  [15:0] io_Stationary_matrix_0_7,
  input  [15:0] io_Stationary_matrix_1_0,
  input  [15:0] io_Stationary_matrix_1_1,
  input  [15:0] io_Stationary_matrix_1_2,
  input  [15:0] io_Stationary_matrix_1_3,
  input  [15:0] io_Stationary_matrix_1_4,
  input  [15:0] io_Stationary_matrix_1_5,
  input  [15:0] io_Stationary_matrix_1_6,
  input  [15:0] io_Stationary_matrix_1_7,
  input  [15:0] io_Stationary_matrix_2_0,
  input  [15:0] io_Stationary_matrix_2_1,
  input  [15:0] io_Stationary_matrix_2_2,
  input  [15:0] io_Stationary_matrix_2_3,
  input  [15:0] io_Stationary_matrix_2_4,
  input  [15:0] io_Stationary_matrix_2_5,
  input  [15:0] io_Stationary_matrix_2_6,
  input  [15:0] io_Stationary_matrix_2_7,
  input  [15:0] io_Stationary_matrix_3_0,
  input  [15:0] io_Stationary_matrix_3_1,
  input  [15:0] io_Stationary_matrix_3_2,
  input  [15:0] io_Stationary_matrix_3_3,
  input  [15:0] io_Stationary_matrix_3_4,
  input  [15:0] io_Stationary_matrix_3_5,
  input  [15:0] io_Stationary_matrix_3_6,
  input  [15:0] io_Stationary_matrix_3_7,
  input  [15:0] io_Stationary_matrix_4_0,
  input  [15:0] io_Stationary_matrix_4_1,
  input  [15:0] io_Stationary_matrix_4_2,
  input  [15:0] io_Stationary_matrix_4_3,
  input  [15:0] io_Stationary_matrix_4_4,
  input  [15:0] io_Stationary_matrix_4_5,
  input  [15:0] io_Stationary_matrix_4_6,
  input  [15:0] io_Stationary_matrix_4_7,
  input  [15:0] io_Stationary_matrix_5_0,
  input  [15:0] io_Stationary_matrix_5_1,
  input  [15:0] io_Stationary_matrix_5_2,
  input  [15:0] io_Stationary_matrix_5_3,
  input  [15:0] io_Stationary_matrix_5_4,
  input  [15:0] io_Stationary_matrix_5_5,
  input  [15:0] io_Stationary_matrix_5_6,
  input  [15:0] io_Stationary_matrix_5_7,
  input  [15:0] io_Stationary_matrix_6_0,
  input  [15:0] io_Stationary_matrix_6_1,
  input  [15:0] io_Stationary_matrix_6_2,
  input  [15:0] io_Stationary_matrix_6_3,
  input  [15:0] io_Stationary_matrix_6_4,
  input  [15:0] io_Stationary_matrix_6_5,
  input  [15:0] io_Stationary_matrix_6_6,
  input  [15:0] io_Stationary_matrix_6_7,
  input  [15:0] io_Stationary_matrix_7_0,
  input  [15:0] io_Stationary_matrix_7_1,
  input  [15:0] io_Stationary_matrix_7_2,
  input  [15:0] io_Stationary_matrix_7_3,
  input  [15:0] io_Stationary_matrix_7_4,
  input  [15:0] io_Stationary_matrix_7_5,
  input  [15:0] io_Stationary_matrix_7_6,
  input  [15:0] io_Stationary_matrix_7_7,
  output [4:0]  io_o_vn_0,
  output [4:0]  io_o_vn_1,
  output [4:0]  io_o_vn_2,
  output [4:0]  io_o_vn_3,
  output [4:0]  io_o_vn2_0,
  output [4:0]  io_o_vn2_1,
  output [4:0]  io_o_vn2_2,
  output [4:0]  io_o_vn2_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
`endif // RANDOMIZE_REG_INIT
  reg [4:0] i_vn_0; // @[ivncontrol4.scala 16:23]
  reg [4:0] i_vn_1; // @[ivncontrol4.scala 16:23]
  reg [4:0] i_vn_2; // @[ivncontrol4.scala 16:23]
  reg [4:0] i_vn_3; // @[ivncontrol4.scala 16:23]
  reg [4:0] i_vn2_0; // @[ivncontrol4.scala 17:24]
  reg [4:0] i_vn2_1; // @[ivncontrol4.scala 17:24]
  reg [4:0] i_vn2_2; // @[ivncontrol4.scala 17:24]
  reg [4:0] i_vn2_3; // @[ivncontrol4.scala 17:24]
  reg [31:0] rowcount_0; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_1; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_2; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_3; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_4; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_5; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_6; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_7; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_8; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_9; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_10; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_11; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_12; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_13; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_14; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_15; // @[ivncontrol4.scala 21:27]
  reg [31:0] pin; // @[ivncontrol4.scala 31:22]
  reg [31:0] i; // @[ivncontrol4.scala 35:20]
  reg [31:0] j; // @[ivncontrol4.scala 36:20]
  wire  _k_T_1 = j == 32'h7; // @[ivncontrol4.scala 38:37]
  wire  _k_T_2 = i == 32'h7 & j == 32'h7; // @[ivncontrol4.scala 38:31]
  reg [31:0] mat_0_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_0_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_0_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_0_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_0_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_0_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_0_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_0_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] count_0; // @[ivncontrol4.scala 52:20]
  reg [31:0] count_1; // @[ivncontrol4.scala 52:20]
  reg [31:0] count_2; // @[ivncontrol4.scala 52:20]
  reg [31:0] count_3; // @[ivncontrol4.scala 52:20]
  reg [31:0] count_4; // @[ivncontrol4.scala 52:20]
  reg [31:0] count_5; // @[ivncontrol4.scala 52:20]
  reg [31:0] count_6; // @[ivncontrol4.scala 52:20]
  reg [31:0] count_7; // @[ivncontrol4.scala 52:20]
  wire [15:0] _GEN_66 = 3'h0 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_0_1 : io_Stationary_matrix_0_0; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_67 = 3'h0 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_0_2 : _GEN_66; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_68 = 3'h0 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_0_3 : _GEN_67; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_69 = 3'h0 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_0_4 : _GEN_68; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_70 = 3'h0 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_0_5 : _GEN_69; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_71 = 3'h0 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_0_6 : _GEN_70; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_72 = 3'h0 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_0_7 : _GEN_71; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_73 = 3'h1 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_1_0 : _GEN_72; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_74 = 3'h1 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_1_1 : _GEN_73; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_75 = 3'h1 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_1_2 : _GEN_74; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_76 = 3'h1 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_1_3 : _GEN_75; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_77 = 3'h1 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_1_4 : _GEN_76; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_78 = 3'h1 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_1_5 : _GEN_77; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_79 = 3'h1 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_1_6 : _GEN_78; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_80 = 3'h1 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_1_7 : _GEN_79; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_81 = 3'h2 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_2_0 : _GEN_80; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_82 = 3'h2 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_2_1 : _GEN_81; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_83 = 3'h2 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_2_2 : _GEN_82; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_84 = 3'h2 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_2_3 : _GEN_83; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_85 = 3'h2 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_2_4 : _GEN_84; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_86 = 3'h2 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_2_5 : _GEN_85; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_87 = 3'h2 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_2_6 : _GEN_86; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_88 = 3'h2 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_2_7 : _GEN_87; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_89 = 3'h3 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_3_0 : _GEN_88; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_90 = 3'h3 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_3_1 : _GEN_89; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_91 = 3'h3 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_3_2 : _GEN_90; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_92 = 3'h3 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_3_3 : _GEN_91; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_93 = 3'h3 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_3_4 : _GEN_92; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_94 = 3'h3 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_3_5 : _GEN_93; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_95 = 3'h3 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_3_6 : _GEN_94; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_96 = 3'h3 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_3_7 : _GEN_95; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_97 = 3'h4 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_4_0 : _GEN_96; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_98 = 3'h4 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_4_1 : _GEN_97; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_99 = 3'h4 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_4_2 : _GEN_98; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_100 = 3'h4 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_4_3 : _GEN_99; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_101 = 3'h4 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_4_4 : _GEN_100; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_102 = 3'h4 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_4_5 : _GEN_101; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_103 = 3'h4 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_4_6 : _GEN_102; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_104 = 3'h4 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_4_7 : _GEN_103; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_105 = 3'h5 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_5_0 : _GEN_104; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_106 = 3'h5 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_5_1 : _GEN_105; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_107 = 3'h5 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_5_2 : _GEN_106; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_108 = 3'h5 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_5_3 : _GEN_107; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_109 = 3'h5 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_5_4 : _GEN_108; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_110 = 3'h5 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_5_5 : _GEN_109; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_111 = 3'h5 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_5_6 : _GEN_110; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_112 = 3'h5 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_5_7 : _GEN_111; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_113 = 3'h6 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_6_0 : _GEN_112; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_114 = 3'h6 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_6_1 : _GEN_113; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_115 = 3'h6 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_6_2 : _GEN_114; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_116 = 3'h6 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_6_3 : _GEN_115; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_117 = 3'h6 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_6_4 : _GEN_116; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_118 = 3'h6 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_6_5 : _GEN_117; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_119 = 3'h6 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_6_6 : _GEN_118; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_120 = 3'h6 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_6_7 : _GEN_119; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_121 = 3'h7 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_7_0 : _GEN_120; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_122 = 3'h7 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_7_1 : _GEN_121; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_123 = 3'h7 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_7_2 : _GEN_122; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_124 = 3'h7 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_7_3 : _GEN_123; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_125 = 3'h7 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_7_4 : _GEN_124; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_126 = 3'h7 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_7_5 : _GEN_125; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_127 = 3'h7 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_7_6 : _GEN_126; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_128 = 3'h7 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_7_7 : _GEN_127; // @[ivncontrol4.scala 57:{15,15}]
  wire [31:0] _mat_T_3_T_4 = {{16'd0}, _GEN_128}; // @[ivncontrol4.scala 57:{15,15}]
  wire  _GEN_225 = count_7 >= 32'h8; // @[ivncontrol4.scala 66:28 67:16]
  wire  valid1 = count_7 >= 32'h8; // @[ivncontrol4.scala 66:28 67:16]
  wire [31:0] _GEN_194 = 3'h1 == i[2:0] ? count_1 : count_0; // @[ivncontrol4.scala 60:{33,33}]
  wire [31:0] _GEN_195 = 3'h2 == i[2:0] ? count_2 : _GEN_194; // @[ivncontrol4.scala 60:{33,33}]
  wire [31:0] _GEN_196 = 3'h3 == i[2:0] ? count_3 : _GEN_195; // @[ivncontrol4.scala 60:{33,33}]
  wire [31:0] _GEN_197 = 3'h4 == i[2:0] ? count_4 : _GEN_196; // @[ivncontrol4.scala 60:{33,33}]
  wire [31:0] _GEN_198 = 3'h5 == i[2:0] ? count_5 : _GEN_197; // @[ivncontrol4.scala 60:{33,33}]
  wire [31:0] _GEN_199 = 3'h6 == i[2:0] ? count_6 : _GEN_198; // @[ivncontrol4.scala 60:{33,33}]
  wire [31:0] _GEN_200 = 3'h7 == i[2:0] ? count_7 : _GEN_199; // @[ivncontrol4.scala 60:{33,33}]
  wire [31:0] _count_T_2 = _GEN_200 + 32'h1; // @[ivncontrol4.scala 60:33]
  wire [31:0] _i_T_1 = i + 32'h1; // @[ivncontrol4.scala 104:16]
  wire [31:0] _j_T_1 = j + 32'h1; // @[ivncontrol4.scala 108:16]
  wire  _GEN_244 = _k_T_2; // @[ivncontrol4.scala 136:75 137:14 139:14]
  wire [31:0] _GEN_245 = rowcount_0 != 32'h0 ? 32'h0 : pin; // @[ivncontrol4.scala 145:30 146:13 31:22]
  wire  _T_27 = rowcount_0 == 32'h0; // @[ivncontrol4.scala 148:23]
  wire [31:0] _GEN_246 = rowcount_0 == 32'h0 & rowcount_1 != 32'h0 ? 32'h1 : _GEN_245; // @[ivncontrol4.scala 148:54 149:13]
  wire  _T_32 = _T_27 & rowcount_1 == 32'h0; // @[ivncontrol4.scala 151:31]
  wire [31:0] _GEN_247 = _T_27 & rowcount_1 == 32'h0 & rowcount_2 != 32'h0 ? 32'h2 : _GEN_246; // @[ivncontrol4.scala 151:77 152:13]
  wire  _T_39 = _T_32 & rowcount_2 == 32'h0; // @[ivncontrol4.scala 154:54]
  wire [31:0] _GEN_248 = _T_32 & rowcount_2 == 32'h0 & rowcount_3 != 32'h0 ? 32'h3 : _GEN_247; // @[ivncontrol4.scala 154:100 155:13]
  wire  _T_48 = _T_39 & rowcount_3 == 32'h0; // @[ivncontrol4.scala 157:77]
  wire [31:0] _GEN_249 = _T_39 & rowcount_3 == 32'h0 & rowcount_4 != 32'h0 ? 32'h4 : _GEN_248; // @[ivncontrol4.scala 157:123 158:13]
  wire  _T_59 = _T_48 & rowcount_4 == 32'h0; // @[ivncontrol4.scala 160:100]
  wire  _T_72 = _T_59 & rowcount_5 == 32'h0; // @[ivncontrol4.scala 163:123]
  wire  valid = _k_T_2; // @[ivncontrol4.scala 136:75 137:14 139:14]
  wire [32:0] _T_91 = {{1'd0}, pin}; // @[ivncontrol4.scala 174:27]
  wire [31:0] _GEN_254 = 4'h1 == _T_91[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_255 = 4'h2 == _T_91[3:0] ? rowcount_2 : _GEN_254; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_256 = 4'h3 == _T_91[3:0] ? rowcount_3 : _GEN_255; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_257 = 4'h4 == _T_91[3:0] ? rowcount_4 : _GEN_256; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_258 = 4'h5 == _T_91[3:0] ? rowcount_5 : _GEN_257; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_259 = 4'h6 == _T_91[3:0] ? rowcount_6 : _GEN_258; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_260 = 4'h7 == _T_91[3:0] ? rowcount_7 : _GEN_259; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_261 = 4'h8 == _T_91[3:0] ? rowcount_8 : _GEN_260; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_262 = 4'h9 == _T_91[3:0] ? rowcount_9 : _GEN_261; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_263 = 4'ha == _T_91[3:0] ? rowcount_10 : _GEN_262; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_264 = 4'hb == _T_91[3:0] ? rowcount_11 : _GEN_263; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_265 = 4'hc == _T_91[3:0] ? rowcount_12 : _GEN_264; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_266 = 4'hd == _T_91[3:0] ? rowcount_13 : _GEN_265; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_267 = 4'he == _T_91[3:0] ? rowcount_14 : _GEN_266; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_268 = 4'hf == _T_91[3:0] ? rowcount_15 : _GEN_267; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_381 = _GEN_268 == 32'h1 ? _T_91[31:0] : 32'h10; // @[ivncontrol4.scala 125:17 224:50 225:21]
  wire [31:0] _GEN_382 = _GEN_268 == 32'h2 ? _T_91[31:0] : _GEN_381; // @[ivncontrol4.scala 220:51 221:21]
  wire [31:0] _GEN_383 = _GEN_268 == 32'h2 ? _T_91[31:0] : 32'h16; // @[ivncontrol4.scala 125:17 220:51 222:21]
  wire [31:0] _GEN_384 = _GEN_268 == 32'h3 ? _T_91[31:0] : _GEN_382; // @[ivncontrol4.scala 215:50 216:21]
  wire [31:0] _GEN_385 = _GEN_268 == 32'h3 ? _T_91[31:0] : _GEN_383; // @[ivncontrol4.scala 215:50 217:21]
  wire [31:0] _GEN_386 = _GEN_268 == 32'h3 ? _T_91[31:0] : 32'h11; // @[ivncontrol4.scala 125:17 215:50 218:21]
  wire [31:0] _GEN_387 = _GEN_268 == 32'h4 ? _T_91[31:0] : _GEN_384; // @[ivncontrol4.scala 207:50 208:21]
  wire [31:0] _GEN_388 = _GEN_268 == 32'h4 ? _T_91[31:0] : _GEN_385; // @[ivncontrol4.scala 207:50 209:21]
  wire [31:0] _GEN_389 = _GEN_268 == 32'h4 ? _T_91[31:0] : _GEN_386; // @[ivncontrol4.scala 207:50 210:21]
  wire [31:0] _GEN_390 = _GEN_268 == 32'h4 ? _T_91[31:0] : 32'hc; // @[ivncontrol4.scala 125:17 207:50 211:21]
  wire [31:0] _GEN_391 = _GEN_268 == 32'h5 ? _T_91[31:0] : _GEN_387; // @[ivncontrol4.scala 200:50 201:21]
  wire [31:0] _GEN_392 = _GEN_268 == 32'h5 ? _T_91[31:0] : _GEN_388; // @[ivncontrol4.scala 200:50 202:21]
  wire [31:0] _GEN_393 = _GEN_268 == 32'h5 ? _T_91[31:0] : _GEN_389; // @[ivncontrol4.scala 200:50 203:21]
  wire [31:0] _GEN_394 = _GEN_268 == 32'h5 ? _T_91[31:0] : _GEN_390; // @[ivncontrol4.scala 200:50 204:21]
  wire [31:0] _GEN_395 = _GEN_268 == 32'h5 ? _T_91[31:0] : 32'h1b; // @[ivncontrol4.scala 126:18 200:50 205:22]
  wire [31:0] _GEN_396 = _GEN_268 == 32'h6 ? _T_91[31:0] : _GEN_391; // @[ivncontrol4.scala 192:52 193:21]
  wire [31:0] _GEN_397 = _GEN_268 == 32'h6 ? _T_91[31:0] : _GEN_392; // @[ivncontrol4.scala 192:52 194:21]
  wire [31:0] _GEN_398 = _GEN_268 == 32'h6 ? _T_91[31:0] : _GEN_393; // @[ivncontrol4.scala 192:52 195:21]
  wire [31:0] _GEN_399 = _GEN_268 == 32'h6 ? _T_91[31:0] : _GEN_394; // @[ivncontrol4.scala 192:52 196:21]
  wire [31:0] _GEN_400 = _GEN_268 == 32'h6 ? _T_91[31:0] : _GEN_395; // @[ivncontrol4.scala 192:52 197:22]
  wire [31:0] _GEN_401 = _GEN_268 == 32'h6 ? _T_91[31:0] : 32'h4; // @[ivncontrol4.scala 126:18 192:52 198:22]
  wire [31:0] _GEN_402 = _GEN_268 == 32'h7 ? _T_91[31:0] : _GEN_396; // @[ivncontrol4.scala 184:52 185:21]
  wire [31:0] _GEN_403 = _GEN_268 == 32'h7 ? _T_91[31:0] : _GEN_397; // @[ivncontrol4.scala 184:52 186:21]
  wire [31:0] _GEN_404 = _GEN_268 == 32'h7 ? _T_91[31:0] : _GEN_398; // @[ivncontrol4.scala 184:52 187:21]
  wire [31:0] _GEN_405 = _GEN_268 == 32'h7 ? _T_91[31:0] : _GEN_399; // @[ivncontrol4.scala 184:52 188:21]
  wire [31:0] _GEN_406 = _GEN_268 == 32'h7 ? _T_91[31:0] : _GEN_400; // @[ivncontrol4.scala 184:52 189:22]
  wire [31:0] _GEN_407 = _GEN_268 == 32'h7 ? _T_91[31:0] : _GEN_401; // @[ivncontrol4.scala 184:52 190:22]
  wire [31:0] _GEN_408 = _GEN_268 == 32'h7 ? _T_91[31:0] : 32'h10; // @[ivncontrol4.scala 126:18 184:52 191:22]
  wire [31:0] _GEN_409 = _GEN_268 >= 32'h8 ? _T_91[31:0] : _GEN_402; // @[ivncontrol4.scala 174:42 175:21]
  wire [31:0] _GEN_410 = _GEN_268 >= 32'h8 ? _T_91[31:0] : _GEN_403; // @[ivncontrol4.scala 174:42 176:21]
  wire [31:0] _GEN_411 = _GEN_268 >= 32'h8 ? _T_91[31:0] : _GEN_404; // @[ivncontrol4.scala 174:42 177:21]
  wire [31:0] _GEN_412 = _GEN_268 >= 32'h8 ? _T_91[31:0] : _GEN_405; // @[ivncontrol4.scala 174:42 178:21]
  wire [31:0] _GEN_413 = _GEN_268 >= 32'h8 ? _T_91[31:0] : _GEN_406; // @[ivncontrol4.scala 174:42 179:22]
  wire [31:0] _GEN_414 = _GEN_268 >= 32'h8 ? _T_91[31:0] : _GEN_407; // @[ivncontrol4.scala 174:42 180:22]
  wire [31:0] _GEN_415 = _GEN_268 >= 32'h8 ? _T_91[31:0] : _GEN_408; // @[ivncontrol4.scala 174:42 181:22]
  wire [31:0] _GEN_416 = _GEN_268 >= 32'h8 ? _T_91[31:0] : 32'h4; // @[ivncontrol4.scala 126:18 174:42 182:22]
  wire [31:0] _T_127 = 32'h8 - _GEN_268; // @[ivncontrol4.scala 228:18]
  wire [31:0] _i_vn_1_T_15 = 32'h1 + pin; // @[ivncontrol4.scala 229:29]
  wire [31:0] _GEN_529 = _T_127 == 32'h1 ? _i_vn_1_T_15 : _GEN_416; // @[ivncontrol4.scala 269:54 272:22]
  wire [31:0] _GEN_530 = _T_127 == 32'h2 ? _i_vn_1_T_15 : _GEN_415; // @[ivncontrol4.scala 264:54 267:22]
  wire [31:0] _GEN_531 = _T_127 == 32'h2 ? _i_vn_1_T_15 : _GEN_529; // @[ivncontrol4.scala 264:54 268:22]
  wire [31:0] _GEN_532 = _T_127 == 32'h3 ? _i_vn_1_T_15 : _GEN_414; // @[ivncontrol4.scala 257:54 259:22]
  wire [31:0] _GEN_533 = _T_127 == 32'h3 ? _i_vn_1_T_15 : _GEN_530; // @[ivncontrol4.scala 257:54 260:22]
  wire [31:0] _GEN_534 = _T_127 == 32'h3 ? _i_vn_1_T_15 : _GEN_531; // @[ivncontrol4.scala 257:54 261:22]
  wire [31:0] _GEN_535 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_413; // @[ivncontrol4.scala 251:54 253:22]
  wire [31:0] _GEN_536 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_532; // @[ivncontrol4.scala 251:54 254:22]
  wire [31:0] _GEN_537 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_533; // @[ivncontrol4.scala 251:54 255:22]
  wire [31:0] _GEN_538 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_534; // @[ivncontrol4.scala 251:54 256:22]
  wire [31:0] _GEN_539 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_412; // @[ivncontrol4.scala 244:54 246:21]
  wire [31:0] _GEN_540 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_535; // @[ivncontrol4.scala 244:54 247:22]
  wire [31:0] _GEN_541 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_536; // @[ivncontrol4.scala 244:54 248:22]
  wire [31:0] _GEN_542 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_537; // @[ivncontrol4.scala 244:54 249:22]
  wire [31:0] _GEN_543 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_538; // @[ivncontrol4.scala 244:54 250:22]
  wire [31:0] _GEN_544 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_411; // @[ivncontrol4.scala 237:54 238:22]
  wire [31:0] _GEN_545 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_539; // @[ivncontrol4.scala 237:54 239:21]
  wire [31:0] _GEN_546 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_540; // @[ivncontrol4.scala 237:54 240:22]
  wire [31:0] _GEN_547 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_541; // @[ivncontrol4.scala 237:54 241:22]
  wire [31:0] _GEN_548 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_542; // @[ivncontrol4.scala 237:54 242:22]
  wire [31:0] _GEN_549 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_543; // @[ivncontrol4.scala 237:54 243:22]
  wire [31:0] _GEN_550 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_410; // @[ivncontrol4.scala 228:49 229:22]
  wire [31:0] _GEN_551 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_544; // @[ivncontrol4.scala 228:49 230:21]
  wire [31:0] _GEN_552 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_545; // @[ivncontrol4.scala 228:49 231:21]
  wire [31:0] _GEN_553 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_546; // @[ivncontrol4.scala 228:49 232:22]
  wire [31:0] _GEN_554 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_547; // @[ivncontrol4.scala 228:49 233:22]
  wire [31:0] _GEN_555 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_548; // @[ivncontrol4.scala 228:49 234:22]
  wire [31:0] _GEN_556 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_549; // @[ivncontrol4.scala 228:49 235:22]
  wire [31:0] _GEN_574 = 4'h1 == _i_vn_1_T_15[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_575 = 4'h2 == _i_vn_1_T_15[3:0] ? rowcount_2 : _GEN_574; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_576 = 4'h3 == _i_vn_1_T_15[3:0] ? rowcount_3 : _GEN_575; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_577 = 4'h4 == _i_vn_1_T_15[3:0] ? rowcount_4 : _GEN_576; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_578 = 4'h5 == _i_vn_1_T_15[3:0] ? rowcount_5 : _GEN_577; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_579 = 4'h6 == _i_vn_1_T_15[3:0] ? rowcount_6 : _GEN_578; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_580 = 4'h7 == _i_vn_1_T_15[3:0] ? rowcount_7 : _GEN_579; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_581 = 4'h8 == _i_vn_1_T_15[3:0] ? rowcount_8 : _GEN_580; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_582 = 4'h9 == _i_vn_1_T_15[3:0] ? rowcount_9 : _GEN_581; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_583 = 4'ha == _i_vn_1_T_15[3:0] ? rowcount_10 : _GEN_582; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_584 = 4'hb == _i_vn_1_T_15[3:0] ? rowcount_11 : _GEN_583; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_585 = 4'hc == _i_vn_1_T_15[3:0] ? rowcount_12 : _GEN_584; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_586 = 4'hd == _i_vn_1_T_15[3:0] ? rowcount_13 : _GEN_585; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_587 = 4'he == _i_vn_1_T_15[3:0] ? rowcount_14 : _GEN_586; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_588 = 4'hf == _i_vn_1_T_15[3:0] ? rowcount_15 : _GEN_587; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _T_172 = _GEN_268 + _GEN_588; // @[ivncontrol4.scala 275:41]
  wire [31:0] _T_174 = 32'h8 - _T_172; // @[ivncontrol4.scala 275:18]
  wire [31:0] _i_vn_1_T_17 = 32'h2 + pin; // @[ivncontrol4.scala 276:29]
  wire [31:0] _GEN_781 = _T_174 == 32'h1 ? _i_vn_1_T_17 : _GEN_556; // @[ivncontrol4.scala 318:78 321:22]
  wire [31:0] _GEN_782 = _T_174 == 32'h2 ? _i_vn_1_T_17 : _GEN_555; // @[ivncontrol4.scala 312:76 315:22]
  wire [31:0] _GEN_783 = _T_174 == 32'h2 ? _i_vn_1_T_17 : _GEN_781; // @[ivncontrol4.scala 312:76 316:22]
  wire [31:0] _GEN_784 = _T_174 == 32'h3 ? _i_vn_1_T_17 : _GEN_554; // @[ivncontrol4.scala 305:78 307:23]
  wire [31:0] _GEN_785 = _T_174 == 32'h3 ? _i_vn_1_T_17 : _GEN_782; // @[ivncontrol4.scala 305:78 308:22]
  wire [31:0] _GEN_786 = _T_174 == 32'h3 ? _i_vn_1_T_17 : _GEN_783; // @[ivncontrol4.scala 305:78 309:22]
  wire [31:0] _GEN_787 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_553; // @[ivncontrol4.scala 299:78 301:22]
  wire [31:0] _GEN_788 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_784; // @[ivncontrol4.scala 299:78 302:22]
  wire [31:0] _GEN_789 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_785; // @[ivncontrol4.scala 299:78 303:22]
  wire [31:0] _GEN_790 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_786; // @[ivncontrol4.scala 299:78 304:22]
  wire [31:0] _GEN_791 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_552; // @[ivncontrol4.scala 292:76 294:23]
  wire [31:0] _GEN_792 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_787; // @[ivncontrol4.scala 292:76 295:22]
  wire [31:0] _GEN_793 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_788; // @[ivncontrol4.scala 292:76 296:22]
  wire [31:0] _GEN_794 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_789; // @[ivncontrol4.scala 292:76 297:22]
  wire [31:0] _GEN_795 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_790; // @[ivncontrol4.scala 292:76 298:22]
  wire [31:0] _GEN_796 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_551; // @[ivncontrol4.scala 284:77 286:22]
  wire [31:0] _GEN_797 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_791; // @[ivncontrol4.scala 284:77 287:21]
  wire [31:0] _GEN_798 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_792; // @[ivncontrol4.scala 284:77 288:22]
  wire [31:0] _GEN_799 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_793; // @[ivncontrol4.scala 284:77 289:22]
  wire [31:0] _GEN_800 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_794; // @[ivncontrol4.scala 284:77 290:22]
  wire [31:0] _GEN_801 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_795; // @[ivncontrol4.scala 284:77 291:22]
  wire [31:0] _GEN_802 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_550; // @[ivncontrol4.scala 275:73 276:22]
  wire [31:0] _GEN_803 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_796; // @[ivncontrol4.scala 275:73 277:21]
  wire [31:0] _GEN_804 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_797; // @[ivncontrol4.scala 275:73 278:21]
  wire [31:0] _GEN_805 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_798; // @[ivncontrol4.scala 275:73 279:22]
  wire [31:0] _GEN_806 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_799; // @[ivncontrol4.scala 275:73 280:22]
  wire [31:0] _GEN_807 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_800; // @[ivncontrol4.scala 275:73 281:22]
  wire [31:0] _GEN_808 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_801; // @[ivncontrol4.scala 275:73 282:22]
  wire [31:0] _GEN_842 = 4'h1 == _i_vn_1_T_17[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_843 = 4'h2 == _i_vn_1_T_17[3:0] ? rowcount_2 : _GEN_842; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_844 = 4'h3 == _i_vn_1_T_17[3:0] ? rowcount_3 : _GEN_843; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_845 = 4'h4 == _i_vn_1_T_17[3:0] ? rowcount_4 : _GEN_844; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_846 = 4'h5 == _i_vn_1_T_17[3:0] ? rowcount_5 : _GEN_845; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_847 = 4'h6 == _i_vn_1_T_17[3:0] ? rowcount_6 : _GEN_846; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_848 = 4'h7 == _i_vn_1_T_17[3:0] ? rowcount_7 : _GEN_847; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_849 = 4'h8 == _i_vn_1_T_17[3:0] ? rowcount_8 : _GEN_848; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_850 = 4'h9 == _i_vn_1_T_17[3:0] ? rowcount_9 : _GEN_849; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_851 = 4'ha == _i_vn_1_T_17[3:0] ? rowcount_10 : _GEN_850; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_852 = 4'hb == _i_vn_1_T_17[3:0] ? rowcount_11 : _GEN_851; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_853 = 4'hc == _i_vn_1_T_17[3:0] ? rowcount_12 : _GEN_852; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_854 = 4'hd == _i_vn_1_T_17[3:0] ? rowcount_13 : _GEN_853; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_855 = 4'he == _i_vn_1_T_17[3:0] ? rowcount_14 : _GEN_854; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_856 = 4'hf == _i_vn_1_T_17[3:0] ? rowcount_15 : _GEN_855; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _T_254 = _T_172 + _GEN_856; // @[ivncontrol4.scala 326:62]
  wire [31:0] _T_256 = 32'h8 - _T_254; // @[ivncontrol4.scala 326:17]
  wire [31:0] _i_vn_1_T_19 = 32'h3 + pin; // @[ivncontrol4.scala 327:29]
  wire [31:0] _GEN_1145 = _T_256 == 32'h1 ? _i_vn_1_T_19 : _GEN_808; // @[ivncontrol4.scala 369:100 372:22]
  wire [31:0] _GEN_1146 = _T_256 == 32'h2 ? _i_vn_1_T_19 : _GEN_807; // @[ivncontrol4.scala 363:98 366:22]
  wire [31:0] _GEN_1147 = _T_256 == 32'h2 ? _i_vn_1_T_19 : _GEN_1145; // @[ivncontrol4.scala 363:98 367:22]
  wire [31:0] _GEN_1148 = _T_256 == 32'h3 ? _i_vn_1_T_19 : _GEN_806; // @[ivncontrol4.scala 356:100 358:23]
  wire [31:0] _GEN_1149 = _T_256 == 32'h3 ? _i_vn_1_T_19 : _GEN_1146; // @[ivncontrol4.scala 356:100 359:22]
  wire [31:0] _GEN_1150 = _T_256 == 32'h3 ? _i_vn_1_T_19 : _GEN_1147; // @[ivncontrol4.scala 356:100 360:22]
  wire [31:0] _GEN_1151 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_805; // @[ivncontrol4.scala 350:100 352:22]
  wire [31:0] _GEN_1152 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_1148; // @[ivncontrol4.scala 350:100 353:22]
  wire [31:0] _GEN_1153 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_1149; // @[ivncontrol4.scala 350:100 354:22]
  wire [31:0] _GEN_1154 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_1150; // @[ivncontrol4.scala 350:100 355:22]
  wire [31:0] _GEN_1155 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_804; // @[ivncontrol4.scala 343:98 345:23]
  wire [31:0] _GEN_1156 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1151; // @[ivncontrol4.scala 343:98 346:22]
  wire [31:0] _GEN_1157 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1152; // @[ivncontrol4.scala 343:98 347:22]
  wire [31:0] _GEN_1158 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1153; // @[ivncontrol4.scala 343:98 348:22]
  wire [31:0] _GEN_1159 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1154; // @[ivncontrol4.scala 343:98 349:22]
  wire [31:0] _GEN_1160 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_803; // @[ivncontrol4.scala 335:99 337:22]
  wire [31:0] _GEN_1161 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1155; // @[ivncontrol4.scala 335:99 338:21]
  wire [31:0] _GEN_1162 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1156; // @[ivncontrol4.scala 335:99 339:22]
  wire [31:0] _GEN_1163 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1157; // @[ivncontrol4.scala 335:99 340:22]
  wire [31:0] _GEN_1164 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1158; // @[ivncontrol4.scala 335:99 341:22]
  wire [31:0] _GEN_1165 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1159; // @[ivncontrol4.scala 335:99 342:22]
  wire [31:0] _GEN_1166 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_802; // @[ivncontrol4.scala 326:94 327:22]
  wire [31:0] _GEN_1167 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1160; // @[ivncontrol4.scala 326:94 328:21]
  wire [31:0] _GEN_1168 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1161; // @[ivncontrol4.scala 326:94 329:21]
  wire [31:0] _GEN_1169 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1162; // @[ivncontrol4.scala 326:94 330:22]
  wire [31:0] _GEN_1170 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1163; // @[ivncontrol4.scala 326:94 331:22]
  wire [31:0] _GEN_1171 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1164; // @[ivncontrol4.scala 326:94 332:22]
  wire [31:0] _GEN_1172 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1165; // @[ivncontrol4.scala 326:94 333:22]
  wire [31:0] _GEN_1222 = 4'h1 == _i_vn_1_T_19[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1223 = 4'h2 == _i_vn_1_T_19[3:0] ? rowcount_2 : _GEN_1222; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1224 = 4'h3 == _i_vn_1_T_19[3:0] ? rowcount_3 : _GEN_1223; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1225 = 4'h4 == _i_vn_1_T_19[3:0] ? rowcount_4 : _GEN_1224; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1226 = 4'h5 == _i_vn_1_T_19[3:0] ? rowcount_5 : _GEN_1225; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1227 = 4'h6 == _i_vn_1_T_19[3:0] ? rowcount_6 : _GEN_1226; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1228 = 4'h7 == _i_vn_1_T_19[3:0] ? rowcount_7 : _GEN_1227; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1229 = 4'h8 == _i_vn_1_T_19[3:0] ? rowcount_8 : _GEN_1228; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1230 = 4'h9 == _i_vn_1_T_19[3:0] ? rowcount_9 : _GEN_1229; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1231 = 4'ha == _i_vn_1_T_19[3:0] ? rowcount_10 : _GEN_1230; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1232 = 4'hb == _i_vn_1_T_19[3:0] ? rowcount_11 : _GEN_1231; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1233 = 4'hc == _i_vn_1_T_19[3:0] ? rowcount_12 : _GEN_1232; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1234 = 4'hd == _i_vn_1_T_19[3:0] ? rowcount_13 : _GEN_1233; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1235 = 4'he == _i_vn_1_T_19[3:0] ? rowcount_14 : _GEN_1234; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1236 = 4'hf == _i_vn_1_T_19[3:0] ? rowcount_15 : _GEN_1235; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _T_371 = _T_254 + _GEN_1236; // @[ivncontrol4.scala 376:86]
  wire [31:0] _T_373 = 32'h8 - _T_371; // @[ivncontrol4.scala 376:19]
  wire [31:0] _i_vn_1_T_21 = 32'h4 + pin; // @[ivncontrol4.scala 377:29]
  wire [31:0] _GEN_1621 = _T_373 == 32'h1 ? _i_vn_1_T_21 : _GEN_1172; // @[ivncontrol4.scala 419:122 422:22]
  wire [31:0] _GEN_1622 = _T_373 == 32'h2 ? _i_vn_1_T_21 : _GEN_1171; // @[ivncontrol4.scala 413:121 416:22]
  wire [31:0] _GEN_1623 = _T_373 == 32'h2 ? _i_vn_1_T_21 : _GEN_1621; // @[ivncontrol4.scala 413:121 417:22]
  wire [31:0] _GEN_1624 = _T_373 == 32'h3 ? _i_vn_1_T_21 : _GEN_1170; // @[ivncontrol4.scala 406:123 408:23]
  wire [31:0] _GEN_1625 = _T_373 == 32'h3 ? _i_vn_1_T_21 : _GEN_1622; // @[ivncontrol4.scala 406:123 409:22]
  wire [31:0] _GEN_1626 = _T_373 == 32'h3 ? _i_vn_1_T_21 : _GEN_1623; // @[ivncontrol4.scala 406:123 410:22]
  wire [31:0] _GEN_1627 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1169; // @[ivncontrol4.scala 400:122 402:22]
  wire [31:0] _GEN_1628 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1624; // @[ivncontrol4.scala 400:122 403:22]
  wire [31:0] _GEN_1629 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1625; // @[ivncontrol4.scala 400:122 404:22]
  wire [31:0] _GEN_1630 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1626; // @[ivncontrol4.scala 400:122 405:22]
  wire [31:0] _GEN_1631 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1168; // @[ivncontrol4.scala 393:121 395:23]
  wire [31:0] _GEN_1632 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1627; // @[ivncontrol4.scala 393:121 396:22]
  wire [31:0] _GEN_1633 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1628; // @[ivncontrol4.scala 393:121 397:22]
  wire [31:0] _GEN_1634 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1629; // @[ivncontrol4.scala 393:121 398:22]
  wire [31:0] _GEN_1635 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1630; // @[ivncontrol4.scala 393:121 399:22]
  wire [31:0] _GEN_1636 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1167; // @[ivncontrol4.scala 385:121 387:22]
  wire [31:0] _GEN_1637 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1631; // @[ivncontrol4.scala 385:121 388:21]
  wire [31:0] _GEN_1638 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1632; // @[ivncontrol4.scala 385:121 389:22]
  wire [31:0] _GEN_1639 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1633; // @[ivncontrol4.scala 385:121 390:22]
  wire [31:0] _GEN_1640 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1634; // @[ivncontrol4.scala 385:121 391:22]
  wire [31:0] _GEN_1641 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1635; // @[ivncontrol4.scala 385:121 392:22]
  wire [31:0] _GEN_1642 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1166; // @[ivncontrol4.scala 376:118 377:22]
  wire [31:0] _GEN_1643 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1636; // @[ivncontrol4.scala 376:118 378:21]
  wire [31:0] _GEN_1644 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1637; // @[ivncontrol4.scala 376:118 379:21]
  wire [31:0] _GEN_1645 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1638; // @[ivncontrol4.scala 376:118 380:22]
  wire [31:0] _GEN_1646 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1639; // @[ivncontrol4.scala 376:118 381:22]
  wire [31:0] _GEN_1647 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1640; // @[ivncontrol4.scala 376:118 382:22]
  wire [31:0] _GEN_1648 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1641; // @[ivncontrol4.scala 376:118 383:22]
  wire [31:0] _GEN_1714 = 4'h1 == _i_vn_1_T_21[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1715 = 4'h2 == _i_vn_1_T_21[3:0] ? rowcount_2 : _GEN_1714; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1716 = 4'h3 == _i_vn_1_T_21[3:0] ? rowcount_3 : _GEN_1715; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1717 = 4'h4 == _i_vn_1_T_21[3:0] ? rowcount_4 : _GEN_1716; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1718 = 4'h5 == _i_vn_1_T_21[3:0] ? rowcount_5 : _GEN_1717; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1719 = 4'h6 == _i_vn_1_T_21[3:0] ? rowcount_6 : _GEN_1718; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1720 = 4'h7 == _i_vn_1_T_21[3:0] ? rowcount_7 : _GEN_1719; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1721 = 4'h8 == _i_vn_1_T_21[3:0] ? rowcount_8 : _GEN_1720; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1722 = 4'h9 == _i_vn_1_T_21[3:0] ? rowcount_9 : _GEN_1721; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1723 = 4'ha == _i_vn_1_T_21[3:0] ? rowcount_10 : _GEN_1722; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1724 = 4'hb == _i_vn_1_T_21[3:0] ? rowcount_11 : _GEN_1723; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1725 = 4'hc == _i_vn_1_T_21[3:0] ? rowcount_12 : _GEN_1724; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1726 = 4'hd == _i_vn_1_T_21[3:0] ? rowcount_13 : _GEN_1725; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1727 = 4'he == _i_vn_1_T_21[3:0] ? rowcount_14 : _GEN_1726; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1728 = 4'hf == _i_vn_1_T_21[3:0] ? rowcount_15 : _GEN_1727; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _T_523 = _T_371 + _GEN_1728; // @[ivncontrol4.scala 426:108]
  wire [31:0] _T_525 = 32'h8 - _T_523; // @[ivncontrol4.scala 426:19]
  wire [31:0] _i_vn_1_T_23 = 32'h5 + pin; // @[ivncontrol4.scala 427:29]
  wire [31:0] _GEN_2209 = _T_525 == 32'h1 ? _i_vn_1_T_23 : _GEN_1648; // @[ivncontrol4.scala 469:144 472:22]
  wire [31:0] _GEN_2210 = _T_525 == 32'h2 ? _i_vn_1_T_23 : _GEN_1647; // @[ivncontrol4.scala 463:143 466:22]
  wire [31:0] _GEN_2211 = _T_525 == 32'h2 ? _i_vn_1_T_23 : _GEN_2209; // @[ivncontrol4.scala 463:143 467:22]
  wire [31:0] _GEN_2212 = _T_525 == 32'h3 ? _i_vn_1_T_23 : _GEN_1646; // @[ivncontrol4.scala 456:145 458:23]
  wire [31:0] _GEN_2213 = _T_525 == 32'h3 ? _i_vn_1_T_23 : _GEN_2210; // @[ivncontrol4.scala 456:145 459:22]
  wire [31:0] _GEN_2214 = _T_525 == 32'h3 ? _i_vn_1_T_23 : _GEN_2211; // @[ivncontrol4.scala 456:145 460:22]
  wire [31:0] _GEN_2215 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_1645; // @[ivncontrol4.scala 450:143 452:22]
  wire [31:0] _GEN_2216 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_2212; // @[ivncontrol4.scala 450:143 453:22]
  wire [31:0] _GEN_2217 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_2213; // @[ivncontrol4.scala 450:143 454:22]
  wire [31:0] _GEN_2218 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_2214; // @[ivncontrol4.scala 450:143 455:22]
  wire [31:0] _GEN_2219 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_1644; // @[ivncontrol4.scala 443:143 445:23]
  wire [31:0] _GEN_2220 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2215; // @[ivncontrol4.scala 443:143 446:22]
  wire [31:0] _GEN_2221 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2216; // @[ivncontrol4.scala 443:143 447:22]
  wire [31:0] _GEN_2222 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2217; // @[ivncontrol4.scala 443:143 448:22]
  wire [31:0] _GEN_2223 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2218; // @[ivncontrol4.scala 443:143 449:22]
  wire [31:0] _GEN_2224 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_1643; // @[ivncontrol4.scala 435:143 437:22]
  wire [31:0] _GEN_2225 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2219; // @[ivncontrol4.scala 435:143 438:21]
  wire [31:0] _GEN_2226 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2220; // @[ivncontrol4.scala 435:143 439:22]
  wire [31:0] _GEN_2227 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2221; // @[ivncontrol4.scala 435:143 440:22]
  wire [31:0] _GEN_2228 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2222; // @[ivncontrol4.scala 435:143 441:22]
  wire [31:0] _GEN_2229 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2223; // @[ivncontrol4.scala 435:143 442:22]
  wire [31:0] _GEN_2230 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_1642; // @[ivncontrol4.scala 426:140 427:22]
  wire [31:0] _GEN_2231 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2224; // @[ivncontrol4.scala 426:140 428:21]
  wire [31:0] _GEN_2232 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2225; // @[ivncontrol4.scala 426:140 429:21]
  wire [31:0] _GEN_2233 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2226; // @[ivncontrol4.scala 426:140 430:22]
  wire [31:0] _GEN_2234 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2227; // @[ivncontrol4.scala 426:140 431:22]
  wire [31:0] _GEN_2235 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2228; // @[ivncontrol4.scala 426:140 432:22]
  wire [31:0] _GEN_2236 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2229; // @[ivncontrol4.scala 426:140 433:22]
  wire [31:0] _GEN_2318 = 4'h1 == _i_vn_1_T_23[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2319 = 4'h2 == _i_vn_1_T_23[3:0] ? rowcount_2 : _GEN_2318; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2320 = 4'h3 == _i_vn_1_T_23[3:0] ? rowcount_3 : _GEN_2319; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2321 = 4'h4 == _i_vn_1_T_23[3:0] ? rowcount_4 : _GEN_2320; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2322 = 4'h5 == _i_vn_1_T_23[3:0] ? rowcount_5 : _GEN_2321; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2323 = 4'h6 == _i_vn_1_T_23[3:0] ? rowcount_6 : _GEN_2322; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2324 = 4'h7 == _i_vn_1_T_23[3:0] ? rowcount_7 : _GEN_2323; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2325 = 4'h8 == _i_vn_1_T_23[3:0] ? rowcount_8 : _GEN_2324; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2326 = 4'h9 == _i_vn_1_T_23[3:0] ? rowcount_9 : _GEN_2325; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2327 = 4'ha == _i_vn_1_T_23[3:0] ? rowcount_10 : _GEN_2326; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2328 = 4'hb == _i_vn_1_T_23[3:0] ? rowcount_11 : _GEN_2327; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2329 = 4'hc == _i_vn_1_T_23[3:0] ? rowcount_12 : _GEN_2328; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2330 = 4'hd == _i_vn_1_T_23[3:0] ? rowcount_13 : _GEN_2329; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2331 = 4'he == _i_vn_1_T_23[3:0] ? rowcount_14 : _GEN_2330; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2332 = 4'hf == _i_vn_1_T_23[3:0] ? rowcount_15 : _GEN_2331; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _T_710 = _T_523 + _GEN_2332; // @[ivncontrol4.scala 477:130]
  wire [31:0] _T_712 = 32'h8 - _T_710; // @[ivncontrol4.scala 477:19]
  wire [31:0] _i_vn_1_T_25 = 32'h6 + pin; // @[ivncontrol4.scala 478:29]
  wire [31:0] _GEN_2909 = _T_712 == 32'h1 ? _i_vn_1_T_25 : _GEN_2236; // @[ivncontrol4.scala 520:166 523:22]
  wire [31:0] _GEN_2910 = _T_712 == 32'h2 ? _i_vn_1_T_25 : _GEN_2235; // @[ivncontrol4.scala 514:166 517:22]
  wire [31:0] _GEN_2911 = _T_712 == 32'h2 ? _i_vn_1_T_25 : _GEN_2909; // @[ivncontrol4.scala 514:166 518:22]
  wire [31:0] _GEN_2912 = _T_712 == 32'h3 ? _i_vn_1_T_25 : _GEN_2234; // @[ivncontrol4.scala 507:168 509:23]
  wire [31:0] _GEN_2913 = _T_712 == 32'h3 ? _i_vn_1_T_25 : _GEN_2910; // @[ivncontrol4.scala 507:168 510:22]
  wire [31:0] _GEN_2914 = _T_712 == 32'h3 ? _i_vn_1_T_25 : _GEN_2911; // @[ivncontrol4.scala 507:168 511:22]
  wire [31:0] _GEN_2915 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2233; // @[ivncontrol4.scala 501:166 503:22]
  wire [31:0] _GEN_2916 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2912; // @[ivncontrol4.scala 501:166 504:22]
  wire [31:0] _GEN_2917 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2913; // @[ivncontrol4.scala 501:166 505:22]
  wire [31:0] _GEN_2918 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2914; // @[ivncontrol4.scala 501:166 506:22]
  wire [31:0] _GEN_2919 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2232; // @[ivncontrol4.scala 494:166 496:23]
  wire [31:0] _GEN_2920 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2915; // @[ivncontrol4.scala 494:166 497:22]
  wire [31:0] _GEN_2921 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2916; // @[ivncontrol4.scala 494:166 498:22]
  wire [31:0] _GEN_2922 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2917; // @[ivncontrol4.scala 494:166 499:22]
  wire [31:0] _GEN_2923 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2918; // @[ivncontrol4.scala 494:166 500:22]
  wire [31:0] _GEN_2924 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2231; // @[ivncontrol4.scala 486:166 488:22]
  wire [31:0] _GEN_2925 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2919; // @[ivncontrol4.scala 486:166 489:21]
  wire [31:0] _GEN_2926 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2920; // @[ivncontrol4.scala 486:166 490:22]
  wire [31:0] _GEN_2927 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2921; // @[ivncontrol4.scala 486:166 491:22]
  wire [31:0] _GEN_2928 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2922; // @[ivncontrol4.scala 486:166 492:22]
  wire [31:0] _GEN_2929 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2923; // @[ivncontrol4.scala 486:166 493:22]
  wire [31:0] _GEN_2930 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2230; // @[ivncontrol4.scala 477:162 478:22]
  wire [31:0] _GEN_2931 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2924; // @[ivncontrol4.scala 477:162 479:21]
  wire [31:0] _GEN_2932 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2925; // @[ivncontrol4.scala 477:162 480:21]
  wire [31:0] _GEN_2933 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2926; // @[ivncontrol4.scala 477:162 481:22]
  wire [31:0] _GEN_2934 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2927; // @[ivncontrol4.scala 477:162 482:22]
  wire [31:0] _GEN_2935 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2928; // @[ivncontrol4.scala 477:162 483:22]
  wire [31:0] _GEN_2936 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2929; // @[ivncontrol4.scala 477:162 484:22]
  wire [31:0] _GEN_3034 = 4'h1 == _i_vn_1_T_25[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3035 = 4'h2 == _i_vn_1_T_25[3:0] ? rowcount_2 : _GEN_3034; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3036 = 4'h3 == _i_vn_1_T_25[3:0] ? rowcount_3 : _GEN_3035; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3037 = 4'h4 == _i_vn_1_T_25[3:0] ? rowcount_4 : _GEN_3036; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3038 = 4'h5 == _i_vn_1_T_25[3:0] ? rowcount_5 : _GEN_3037; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3039 = 4'h6 == _i_vn_1_T_25[3:0] ? rowcount_6 : _GEN_3038; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3040 = 4'h7 == _i_vn_1_T_25[3:0] ? rowcount_7 : _GEN_3039; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3041 = 4'h8 == _i_vn_1_T_25[3:0] ? rowcount_8 : _GEN_3040; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3042 = 4'h9 == _i_vn_1_T_25[3:0] ? rowcount_9 : _GEN_3041; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3043 = 4'ha == _i_vn_1_T_25[3:0] ? rowcount_10 : _GEN_3042; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3044 = 4'hb == _i_vn_1_T_25[3:0] ? rowcount_11 : _GEN_3043; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3045 = 4'hc == _i_vn_1_T_25[3:0] ? rowcount_12 : _GEN_3044; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3046 = 4'hd == _i_vn_1_T_25[3:0] ? rowcount_13 : _GEN_3045; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3047 = 4'he == _i_vn_1_T_25[3:0] ? rowcount_14 : _GEN_3046; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3048 = 4'hf == _i_vn_1_T_25[3:0] ? rowcount_15 : _GEN_3047; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _T_932 = _T_710 + _GEN_3048; // @[ivncontrol4.scala 528:152]
  wire [31:0] _T_934 = 32'h8 - _T_932; // @[ivncontrol4.scala 528:19]
  wire [31:0] _i_vn_1_T_27 = 32'h7 + pin; // @[ivncontrol4.scala 529:29]
  wire [31:0] _GEN_3721 = _T_934 == 32'h1 ? _i_vn_1_T_27 : _GEN_2936; // @[ivncontrol4.scala 571:188 574:22]
  wire [31:0] _GEN_3722 = _T_934 == 32'h2 ? _i_vn_1_T_27 : _GEN_2935; // @[ivncontrol4.scala 565:188 568:22]
  wire [31:0] _GEN_3723 = _T_934 == 32'h2 ? _i_vn_1_T_27 : _GEN_3721; // @[ivncontrol4.scala 565:188 569:22]
  wire [31:0] _GEN_3724 = _T_934 == 32'h3 ? _i_vn_1_T_27 : _GEN_2934; // @[ivncontrol4.scala 558:190 560:23]
  wire [31:0] _GEN_3725 = _T_934 == 32'h3 ? _i_vn_1_T_27 : _GEN_3722; // @[ivncontrol4.scala 558:190 561:22]
  wire [31:0] _GEN_3726 = _T_934 == 32'h3 ? _i_vn_1_T_27 : _GEN_3723; // @[ivncontrol4.scala 558:190 562:22]
  wire [31:0] _GEN_3727 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_2933; // @[ivncontrol4.scala 552:188 554:22]
  wire [31:0] _GEN_3728 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_3724; // @[ivncontrol4.scala 552:188 555:22]
  wire [31:0] _GEN_3729 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_3725; // @[ivncontrol4.scala 552:188 556:22]
  wire [31:0] _GEN_3730 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_3726; // @[ivncontrol4.scala 552:188 557:22]
  wire [31:0] _GEN_3731 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_2932; // @[ivncontrol4.scala 545:188 547:23]
  wire [31:0] _GEN_3732 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3727; // @[ivncontrol4.scala 545:188 548:22]
  wire [31:0] _GEN_3733 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3728; // @[ivncontrol4.scala 545:188 549:22]
  wire [31:0] _GEN_3734 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3729; // @[ivncontrol4.scala 545:188 550:22]
  wire [31:0] _GEN_3735 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3730; // @[ivncontrol4.scala 545:188 551:22]
  wire [31:0] _GEN_3736 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_2931; // @[ivncontrol4.scala 537:188 539:22]
  wire [31:0] _GEN_3737 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3731; // @[ivncontrol4.scala 537:188 540:21]
  wire [31:0] _GEN_3738 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3732; // @[ivncontrol4.scala 537:188 541:22]
  wire [31:0] _GEN_3739 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3733; // @[ivncontrol4.scala 537:188 542:22]
  wire [31:0] _GEN_3740 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3734; // @[ivncontrol4.scala 537:188 543:22]
  wire [31:0] _GEN_3741 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3735; // @[ivncontrol4.scala 537:188 544:22]
  wire [31:0] _GEN_3742 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_2930; // @[ivncontrol4.scala 528:184 529:22]
  wire [31:0] _GEN_3743 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3736; // @[ivncontrol4.scala 528:184 530:21]
  wire [31:0] _GEN_3744 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3737; // @[ivncontrol4.scala 528:184 531:21]
  wire [31:0] _GEN_3745 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3738; // @[ivncontrol4.scala 528:184 532:22]
  wire [31:0] _GEN_3746 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3739; // @[ivncontrol4.scala 528:184 533:22]
  wire [31:0] _GEN_3747 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3740; // @[ivncontrol4.scala 528:184 534:22]
  wire [31:0] _GEN_3748 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3741; // @[ivncontrol4.scala 528:184 535:22]
  wire [31:0] _GEN_3749 = _GEN_244 ? _GEN_409 : 32'h10; // @[ivncontrol4.scala 125:17 172:28]
  wire [31:0] _GEN_3750 = _GEN_244 ? _GEN_3742 : 32'h16; // @[ivncontrol4.scala 125:17 172:28]
  wire [31:0] _GEN_3751 = _GEN_244 ? _GEN_3743 : 32'h11; // @[ivncontrol4.scala 125:17 172:28]
  wire [31:0] _GEN_3752 = _GEN_244 ? _GEN_3744 : 32'hc; // @[ivncontrol4.scala 125:17 172:28]
  wire [31:0] _GEN_3753 = _GEN_244 ? _GEN_3745 : 32'h1b; // @[ivncontrol4.scala 126:18 172:28]
  wire [31:0] _GEN_3754 = _GEN_244 ? _GEN_3746 : 32'h4; // @[ivncontrol4.scala 126:18 172:28]
  wire [31:0] _GEN_3755 = _GEN_244 ? _GEN_3747 : 32'h10; // @[ivncontrol4.scala 126:18 172:28]
  wire [31:0] _GEN_3756 = _GEN_244 ? _GEN_3748 : 32'h4; // @[ivncontrol4.scala 126:18 172:28]
  wire [31:0] _GEN_4137 = reset ? 32'h0 : _GEN_3749; // @[ivncontrol4.scala 16:{23,23}]
  wire [31:0] _GEN_4138 = reset ? 32'h0 : _GEN_3750; // @[ivncontrol4.scala 16:{23,23}]
  wire [31:0] _GEN_4139 = reset ? 32'h0 : _GEN_3751; // @[ivncontrol4.scala 16:{23,23}]
  wire [31:0] _GEN_4140 = reset ? 32'h0 : _GEN_3752; // @[ivncontrol4.scala 16:{23,23}]
  wire [31:0] _GEN_4141 = reset ? 32'h0 : _GEN_3753; // @[ivncontrol4.scala 17:{24,24}]
  wire [31:0] _GEN_4142 = reset ? 32'h0 : _GEN_3754; // @[ivncontrol4.scala 17:{24,24}]
  wire [31:0] _GEN_4143 = reset ? 32'h0 : _GEN_3755; // @[ivncontrol4.scala 17:{24,24}]
  wire [31:0] _GEN_4144 = reset ? 32'h0 : _GEN_3756; // @[ivncontrol4.scala 17:{24,24}]
  assign io_o_vn_0 = i_vn_0; // @[ivncontrol4.scala 121:13]
  assign io_o_vn_1 = i_vn_1; // @[ivncontrol4.scala 121:13]
  assign io_o_vn_2 = i_vn_2; // @[ivncontrol4.scala 121:13]
  assign io_o_vn_3 = i_vn_3; // @[ivncontrol4.scala 121:13]
  assign io_o_vn2_0 = i_vn2_0; // @[ivncontrol4.scala 122:14]
  assign io_o_vn2_1 = i_vn2_1; // @[ivncontrol4.scala 122:14]
  assign io_o_vn2_2 = i_vn2_2; // @[ivncontrol4.scala 122:14]
  assign io_o_vn2_3 = i_vn2_3; // @[ivncontrol4.scala 122:14]
  always @(posedge clock) begin
    i_vn_0 <= _GEN_4137[4:0]; // @[ivncontrol4.scala 16:{23,23}]
    i_vn_1 <= _GEN_4138[4:0]; // @[ivncontrol4.scala 16:{23,23}]
    i_vn_2 <= _GEN_4139[4:0]; // @[ivncontrol4.scala 16:{23,23}]
    i_vn_3 <= _GEN_4140[4:0]; // @[ivncontrol4.scala 16:{23,23}]
    i_vn2_0 <= _GEN_4141[4:0]; // @[ivncontrol4.scala 17:{24,24}]
    i_vn2_1 <= _GEN_4142[4:0]; // @[ivncontrol4.scala 17:{24,24}]
    i_vn2_2 <= _GEN_4143[4:0]; // @[ivncontrol4.scala 17:{24,24}]
    i_vn2_3 <= _GEN_4144[4:0]; // @[ivncontrol4.scala 17:{24,24}]
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_0 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_0 <= count_0; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_1 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_1 <= count_1; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_2 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_2 <= count_2; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_3 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_3 <= count_3; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_4 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_4 <= count_4; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_5 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_5 <= count_5; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_6 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_6 <= count_6; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_7 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_7 <= count_7; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_8 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_8 <= 32'h0; // @[ivncontrol4.scala 81:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_9 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_9 <= 32'h0; // @[ivncontrol4.scala 81:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_10 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_10 <= 32'h0; // @[ivncontrol4.scala 81:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_11 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_11 <= 32'h0; // @[ivncontrol4.scala 81:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_12 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_12 <= 32'h0; // @[ivncontrol4.scala 81:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_13 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_13 <= 32'h0; // @[ivncontrol4.scala 81:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_14 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_14 <= 32'h0; // @[ivncontrol4.scala 81:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_15 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end
    if (reset) begin // @[ivncontrol4.scala 31:22]
      pin <= 32'h0; // @[ivncontrol4.scala 31:22]
    end else if (_T_72 & rowcount_6 == 32'h0 & rowcount_7 != 32'h0) begin // @[ivncontrol4.scala 166:192]
      pin <= 32'h7; // @[ivncontrol4.scala 167:13]
    end else if (_T_59 & rowcount_5 == 32'h0 & rowcount_6 != 32'h0) begin // @[ivncontrol4.scala 163:169]
      pin <= 32'h6; // @[ivncontrol4.scala 164:13]
    end else if (_T_48 & rowcount_4 == 32'h0 & rowcount_5 != 32'h0) begin // @[ivncontrol4.scala 160:146]
      pin <= 32'h5; // @[ivncontrol4.scala 161:13]
    end else begin
      pin <= _GEN_249;
    end
    if (reset) begin // @[ivncontrol4.scala 35:20]
      i <= 32'h0; // @[ivncontrol4.scala 35:20]
    end else if (i < 32'h7 & _k_T_1) begin // @[ivncontrol4.scala 103:74]
      i <= _i_T_1; // @[ivncontrol4.scala 104:11]
    end
    if (reset) begin // @[ivncontrol4.scala 36:20]
      j <= 32'h0; // @[ivncontrol4.scala 36:20]
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 107:71]
      j <= _j_T_1; // @[ivncontrol4.scala 108:11]
    end else if (!(_k_T_2)) begin // @[ivncontrol4.scala 110:81]
      j <= 32'h0; // @[ivncontrol4.scala 114:11]
    end
    if (3'h0 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h0 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h0 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h0 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h0 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h0 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h0 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h0 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h0 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_0 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h1 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_1 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h2 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_2 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h3 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_3 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h4 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_4 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h5 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_5 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h6 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_6 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h7 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_7 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  i_vn_0 = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  i_vn_1 = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  i_vn_2 = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  i_vn_3 = _RAND_3[4:0];
  _RAND_4 = {1{`RANDOM}};
  i_vn2_0 = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  i_vn2_1 = _RAND_5[4:0];
  _RAND_6 = {1{`RANDOM}};
  i_vn2_2 = _RAND_6[4:0];
  _RAND_7 = {1{`RANDOM}};
  i_vn2_3 = _RAND_7[4:0];
  _RAND_8 = {1{`RANDOM}};
  rowcount_0 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  rowcount_1 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  rowcount_2 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  rowcount_3 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  rowcount_4 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  rowcount_5 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  rowcount_6 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  rowcount_7 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  rowcount_8 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  rowcount_9 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  rowcount_10 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  rowcount_11 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  rowcount_12 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  rowcount_13 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  rowcount_14 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  rowcount_15 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  pin = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  i = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  j = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  mat_0_0 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  mat_0_1 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  mat_0_2 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  mat_0_3 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  mat_0_4 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  mat_0_5 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  mat_0_6 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  mat_0_7 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  mat_1_0 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  mat_1_1 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  mat_1_2 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  mat_1_3 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  mat_1_4 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  mat_1_5 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  mat_1_6 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  mat_1_7 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  mat_2_0 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  mat_2_1 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  mat_2_2 = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  mat_2_3 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  mat_2_4 = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  mat_2_5 = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  mat_2_6 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  mat_2_7 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  mat_3_0 = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  mat_3_1 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  mat_3_2 = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  mat_3_3 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  mat_3_4 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  mat_3_5 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  mat_3_6 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  mat_3_7 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  mat_4_0 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  mat_4_1 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  mat_4_2 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  mat_4_3 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  mat_4_4 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  mat_4_5 = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  mat_4_6 = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  mat_4_7 = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  mat_5_0 = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  mat_5_1 = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  mat_5_2 = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  mat_5_3 = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  mat_5_4 = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  mat_5_5 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  mat_5_6 = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  mat_5_7 = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  mat_6_0 = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  mat_6_1 = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  mat_6_2 = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  mat_6_3 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  mat_6_4 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  mat_6_5 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  mat_6_6 = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  mat_6_7 = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  mat_7_0 = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  mat_7_1 = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  mat_7_2 = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  mat_7_3 = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  mat_7_4 = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  mat_7_5 = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  mat_7_6 = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  mat_7_7 = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  count_0 = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  count_1 = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  count_2 = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  count_3 = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  count_4 = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  count_5 = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  count_6 = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  count_7 = _RAND_98[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ivncontrol4_7(
  input         clock,
  input         reset,
  input  [15:0] io_Stationary_matrix_0_0,
  input  [15:0] io_Stationary_matrix_0_1,
  input  [15:0] io_Stationary_matrix_0_2,
  input  [15:0] io_Stationary_matrix_0_3,
  input  [15:0] io_Stationary_matrix_0_4,
  input  [15:0] io_Stationary_matrix_0_5,
  input  [15:0] io_Stationary_matrix_0_6,
  input  [15:0] io_Stationary_matrix_0_7,
  input  [15:0] io_Stationary_matrix_1_0,
  input  [15:0] io_Stationary_matrix_1_1,
  input  [15:0] io_Stationary_matrix_1_2,
  input  [15:0] io_Stationary_matrix_1_3,
  input  [15:0] io_Stationary_matrix_1_4,
  input  [15:0] io_Stationary_matrix_1_5,
  input  [15:0] io_Stationary_matrix_1_6,
  input  [15:0] io_Stationary_matrix_1_7,
  input  [15:0] io_Stationary_matrix_2_0,
  input  [15:0] io_Stationary_matrix_2_1,
  input  [15:0] io_Stationary_matrix_2_2,
  input  [15:0] io_Stationary_matrix_2_3,
  input  [15:0] io_Stationary_matrix_2_4,
  input  [15:0] io_Stationary_matrix_2_5,
  input  [15:0] io_Stationary_matrix_2_6,
  input  [15:0] io_Stationary_matrix_2_7,
  input  [15:0] io_Stationary_matrix_3_0,
  input  [15:0] io_Stationary_matrix_3_1,
  input  [15:0] io_Stationary_matrix_3_2,
  input  [15:0] io_Stationary_matrix_3_3,
  input  [15:0] io_Stationary_matrix_3_4,
  input  [15:0] io_Stationary_matrix_3_5,
  input  [15:0] io_Stationary_matrix_3_6,
  input  [15:0] io_Stationary_matrix_3_7,
  input  [15:0] io_Stationary_matrix_4_0,
  input  [15:0] io_Stationary_matrix_4_1,
  input  [15:0] io_Stationary_matrix_4_2,
  input  [15:0] io_Stationary_matrix_4_3,
  input  [15:0] io_Stationary_matrix_4_4,
  input  [15:0] io_Stationary_matrix_4_5,
  input  [15:0] io_Stationary_matrix_4_6,
  input  [15:0] io_Stationary_matrix_4_7,
  input  [15:0] io_Stationary_matrix_5_0,
  input  [15:0] io_Stationary_matrix_5_1,
  input  [15:0] io_Stationary_matrix_5_2,
  input  [15:0] io_Stationary_matrix_5_3,
  input  [15:0] io_Stationary_matrix_5_4,
  input  [15:0] io_Stationary_matrix_5_5,
  input  [15:0] io_Stationary_matrix_5_6,
  input  [15:0] io_Stationary_matrix_5_7,
  input  [15:0] io_Stationary_matrix_6_0,
  input  [15:0] io_Stationary_matrix_6_1,
  input  [15:0] io_Stationary_matrix_6_2,
  input  [15:0] io_Stationary_matrix_6_3,
  input  [15:0] io_Stationary_matrix_6_4,
  input  [15:0] io_Stationary_matrix_6_5,
  input  [15:0] io_Stationary_matrix_6_6,
  input  [15:0] io_Stationary_matrix_6_7,
  input  [15:0] io_Stationary_matrix_7_0,
  input  [15:0] io_Stationary_matrix_7_1,
  input  [15:0] io_Stationary_matrix_7_2,
  input  [15:0] io_Stationary_matrix_7_3,
  input  [15:0] io_Stationary_matrix_7_4,
  input  [15:0] io_Stationary_matrix_7_5,
  input  [15:0] io_Stationary_matrix_7_6,
  input  [15:0] io_Stationary_matrix_7_7,
  output [4:0]  io_o_vn_0,
  output [4:0]  io_o_vn_1,
  output [4:0]  io_o_vn_2,
  output [4:0]  io_o_vn_3,
  output [4:0]  io_o_vn2_0,
  output [4:0]  io_o_vn2_1,
  output [4:0]  io_o_vn2_2,
  output [4:0]  io_o_vn2_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
`endif // RANDOMIZE_REG_INIT
  reg [4:0] i_vn_0; // @[ivncontrol4.scala 16:23]
  reg [4:0] i_vn_1; // @[ivncontrol4.scala 16:23]
  reg [4:0] i_vn_2; // @[ivncontrol4.scala 16:23]
  reg [4:0] i_vn_3; // @[ivncontrol4.scala 16:23]
  reg [4:0] i_vn2_0; // @[ivncontrol4.scala 17:24]
  reg [4:0] i_vn2_1; // @[ivncontrol4.scala 17:24]
  reg [4:0] i_vn2_2; // @[ivncontrol4.scala 17:24]
  reg [4:0] i_vn2_3; // @[ivncontrol4.scala 17:24]
  reg [31:0] rowcount_0; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_1; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_2; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_3; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_4; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_5; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_6; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_7; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_8; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_9; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_10; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_11; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_12; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_13; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_14; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_15; // @[ivncontrol4.scala 21:27]
  reg [31:0] pin; // @[ivncontrol4.scala 31:22]
  reg [31:0] i; // @[ivncontrol4.scala 35:20]
  reg [31:0] j; // @[ivncontrol4.scala 36:20]
  wire  _k_T_1 = j == 32'h7; // @[ivncontrol4.scala 38:37]
  wire  _k_T_2 = i == 32'h7 & j == 32'h7; // @[ivncontrol4.scala 38:31]
  reg [31:0] mat_0_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_0_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_0_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_0_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_0_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_0_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_0_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_0_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_1_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_2_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_3_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_4_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_5_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_6_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_0; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_1; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_2; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_3; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_4; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_5; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_6; // @[ivncontrol4.scala 48:18]
  reg [31:0] mat_7_7; // @[ivncontrol4.scala 48:18]
  reg [31:0] count_0; // @[ivncontrol4.scala 52:20]
  reg [31:0] count_1; // @[ivncontrol4.scala 52:20]
  reg [31:0] count_2; // @[ivncontrol4.scala 52:20]
  reg [31:0] count_3; // @[ivncontrol4.scala 52:20]
  reg [31:0] count_4; // @[ivncontrol4.scala 52:20]
  reg [31:0] count_5; // @[ivncontrol4.scala 52:20]
  reg [31:0] count_6; // @[ivncontrol4.scala 52:20]
  reg [31:0] count_7; // @[ivncontrol4.scala 52:20]
  wire [15:0] _GEN_66 = 3'h0 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_0_1 : io_Stationary_matrix_0_0; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_67 = 3'h0 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_0_2 : _GEN_66; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_68 = 3'h0 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_0_3 : _GEN_67; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_69 = 3'h0 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_0_4 : _GEN_68; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_70 = 3'h0 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_0_5 : _GEN_69; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_71 = 3'h0 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_0_6 : _GEN_70; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_72 = 3'h0 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_0_7 : _GEN_71; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_73 = 3'h1 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_1_0 : _GEN_72; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_74 = 3'h1 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_1_1 : _GEN_73; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_75 = 3'h1 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_1_2 : _GEN_74; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_76 = 3'h1 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_1_3 : _GEN_75; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_77 = 3'h1 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_1_4 : _GEN_76; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_78 = 3'h1 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_1_5 : _GEN_77; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_79 = 3'h1 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_1_6 : _GEN_78; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_80 = 3'h1 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_1_7 : _GEN_79; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_81 = 3'h2 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_2_0 : _GEN_80; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_82 = 3'h2 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_2_1 : _GEN_81; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_83 = 3'h2 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_2_2 : _GEN_82; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_84 = 3'h2 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_2_3 : _GEN_83; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_85 = 3'h2 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_2_4 : _GEN_84; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_86 = 3'h2 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_2_5 : _GEN_85; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_87 = 3'h2 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_2_6 : _GEN_86; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_88 = 3'h2 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_2_7 : _GEN_87; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_89 = 3'h3 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_3_0 : _GEN_88; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_90 = 3'h3 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_3_1 : _GEN_89; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_91 = 3'h3 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_3_2 : _GEN_90; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_92 = 3'h3 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_3_3 : _GEN_91; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_93 = 3'h3 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_3_4 : _GEN_92; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_94 = 3'h3 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_3_5 : _GEN_93; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_95 = 3'h3 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_3_6 : _GEN_94; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_96 = 3'h3 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_3_7 : _GEN_95; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_97 = 3'h4 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_4_0 : _GEN_96; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_98 = 3'h4 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_4_1 : _GEN_97; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_99 = 3'h4 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_4_2 : _GEN_98; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_100 = 3'h4 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_4_3 : _GEN_99; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_101 = 3'h4 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_4_4 : _GEN_100; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_102 = 3'h4 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_4_5 : _GEN_101; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_103 = 3'h4 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_4_6 : _GEN_102; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_104 = 3'h4 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_4_7 : _GEN_103; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_105 = 3'h5 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_5_0 : _GEN_104; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_106 = 3'h5 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_5_1 : _GEN_105; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_107 = 3'h5 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_5_2 : _GEN_106; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_108 = 3'h5 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_5_3 : _GEN_107; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_109 = 3'h5 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_5_4 : _GEN_108; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_110 = 3'h5 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_5_5 : _GEN_109; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_111 = 3'h5 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_5_6 : _GEN_110; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_112 = 3'h5 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_5_7 : _GEN_111; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_113 = 3'h6 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_6_0 : _GEN_112; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_114 = 3'h6 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_6_1 : _GEN_113; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_115 = 3'h6 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_6_2 : _GEN_114; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_116 = 3'h6 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_6_3 : _GEN_115; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_117 = 3'h6 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_6_4 : _GEN_116; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_118 = 3'h6 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_6_5 : _GEN_117; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_119 = 3'h6 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_6_6 : _GEN_118; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_120 = 3'h6 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_6_7 : _GEN_119; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_121 = 3'h7 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_7_0 : _GEN_120; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_122 = 3'h7 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_7_1 : _GEN_121; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_123 = 3'h7 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_7_2 : _GEN_122; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_124 = 3'h7 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_7_3 : _GEN_123; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_125 = 3'h7 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_7_4 : _GEN_124; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_126 = 3'h7 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_7_5 : _GEN_125; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_127 = 3'h7 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_7_6 : _GEN_126; // @[ivncontrol4.scala 57:{15,15}]
  wire [15:0] _GEN_128 = 3'h7 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_7_7 : _GEN_127; // @[ivncontrol4.scala 57:{15,15}]
  wire [31:0] _mat_T_3_T_4 = {{16'd0}, _GEN_128}; // @[ivncontrol4.scala 57:{15,15}]
  wire  _GEN_225 = count_7 >= 32'h8; // @[ivncontrol4.scala 66:28 67:16]
  wire  valid1 = count_7 >= 32'h8; // @[ivncontrol4.scala 66:28 67:16]
  wire [31:0] _GEN_194 = 3'h1 == i[2:0] ? count_1 : count_0; // @[ivncontrol4.scala 60:{33,33}]
  wire [31:0] _GEN_195 = 3'h2 == i[2:0] ? count_2 : _GEN_194; // @[ivncontrol4.scala 60:{33,33}]
  wire [31:0] _GEN_196 = 3'h3 == i[2:0] ? count_3 : _GEN_195; // @[ivncontrol4.scala 60:{33,33}]
  wire [31:0] _GEN_197 = 3'h4 == i[2:0] ? count_4 : _GEN_196; // @[ivncontrol4.scala 60:{33,33}]
  wire [31:0] _GEN_198 = 3'h5 == i[2:0] ? count_5 : _GEN_197; // @[ivncontrol4.scala 60:{33,33}]
  wire [31:0] _GEN_199 = 3'h6 == i[2:0] ? count_6 : _GEN_198; // @[ivncontrol4.scala 60:{33,33}]
  wire [31:0] _GEN_200 = 3'h7 == i[2:0] ? count_7 : _GEN_199; // @[ivncontrol4.scala 60:{33,33}]
  wire [31:0] _count_T_2 = _GEN_200 + 32'h1; // @[ivncontrol4.scala 60:33]
  wire [31:0] _i_T_1 = i + 32'h1; // @[ivncontrol4.scala 104:16]
  wire [31:0] _j_T_1 = j + 32'h1; // @[ivncontrol4.scala 108:16]
  wire  _GEN_244 = _k_T_2; // @[ivncontrol4.scala 136:75 137:14 139:14]
  wire [31:0] _GEN_245 = rowcount_0 != 32'h0 ? 32'h0 : pin; // @[ivncontrol4.scala 145:30 146:13 31:22]
  wire  _T_27 = rowcount_0 == 32'h0; // @[ivncontrol4.scala 148:23]
  wire [31:0] _GEN_246 = rowcount_0 == 32'h0 & rowcount_1 != 32'h0 ? 32'h1 : _GEN_245; // @[ivncontrol4.scala 148:54 149:13]
  wire  _T_32 = _T_27 & rowcount_1 == 32'h0; // @[ivncontrol4.scala 151:31]
  wire [31:0] _GEN_247 = _T_27 & rowcount_1 == 32'h0 & rowcount_2 != 32'h0 ? 32'h2 : _GEN_246; // @[ivncontrol4.scala 151:77 152:13]
  wire  _T_39 = _T_32 & rowcount_2 == 32'h0; // @[ivncontrol4.scala 154:54]
  wire [31:0] _GEN_248 = _T_32 & rowcount_2 == 32'h0 & rowcount_3 != 32'h0 ? 32'h3 : _GEN_247; // @[ivncontrol4.scala 154:100 155:13]
  wire  _T_48 = _T_39 & rowcount_3 == 32'h0; // @[ivncontrol4.scala 157:77]
  wire [31:0] _GEN_249 = _T_39 & rowcount_3 == 32'h0 & rowcount_4 != 32'h0 ? 32'h4 : _GEN_248; // @[ivncontrol4.scala 157:123 158:13]
  wire  _T_59 = _T_48 & rowcount_4 == 32'h0; // @[ivncontrol4.scala 160:100]
  wire  _T_72 = _T_59 & rowcount_5 == 32'h0; // @[ivncontrol4.scala 163:123]
  wire  valid = _k_T_2; // @[ivncontrol4.scala 136:75 137:14 139:14]
  wire [32:0] _T_91 = {{1'd0}, pin}; // @[ivncontrol4.scala 174:27]
  wire [31:0] _GEN_254 = 4'h1 == _T_91[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_255 = 4'h2 == _T_91[3:0] ? rowcount_2 : _GEN_254; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_256 = 4'h3 == _T_91[3:0] ? rowcount_3 : _GEN_255; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_257 = 4'h4 == _T_91[3:0] ? rowcount_4 : _GEN_256; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_258 = 4'h5 == _T_91[3:0] ? rowcount_5 : _GEN_257; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_259 = 4'h6 == _T_91[3:0] ? rowcount_6 : _GEN_258; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_260 = 4'h7 == _T_91[3:0] ? rowcount_7 : _GEN_259; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_261 = 4'h8 == _T_91[3:0] ? rowcount_8 : _GEN_260; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_262 = 4'h9 == _T_91[3:0] ? rowcount_9 : _GEN_261; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_263 = 4'ha == _T_91[3:0] ? rowcount_10 : _GEN_262; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_264 = 4'hb == _T_91[3:0] ? rowcount_11 : _GEN_263; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_265 = 4'hc == _T_91[3:0] ? rowcount_12 : _GEN_264; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_266 = 4'hd == _T_91[3:0] ? rowcount_13 : _GEN_265; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_267 = 4'he == _T_91[3:0] ? rowcount_14 : _GEN_266; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_268 = 4'hf == _T_91[3:0] ? rowcount_15 : _GEN_267; // @[ivncontrol4.scala 174:{35,35}]
  wire [31:0] _GEN_381 = _GEN_268 == 32'h1 ? _T_91[31:0] : 32'h1d; // @[ivncontrol4.scala 125:17 224:50 225:21]
  wire [31:0] _GEN_382 = _GEN_268 == 32'h2 ? _T_91[31:0] : _GEN_381; // @[ivncontrol4.scala 220:51 221:21]
  wire [31:0] _GEN_383 = _GEN_268 == 32'h2 ? _T_91[31:0] : 32'h0; // @[ivncontrol4.scala 125:17 220:51 222:21]
  wire [31:0] _GEN_384 = _GEN_268 == 32'h3 ? _T_91[31:0] : _GEN_382; // @[ivncontrol4.scala 215:50 216:21]
  wire [31:0] _GEN_385 = _GEN_268 == 32'h3 ? _T_91[31:0] : _GEN_383; // @[ivncontrol4.scala 215:50 217:21]
  wire [31:0] _GEN_386 = _GEN_268 == 32'h3 ? _T_91[31:0] : 32'h17; // @[ivncontrol4.scala 125:17 215:50 218:21]
  wire [31:0] _GEN_387 = _GEN_268 == 32'h4 ? _T_91[31:0] : _GEN_384; // @[ivncontrol4.scala 207:50 208:21]
  wire [31:0] _GEN_388 = _GEN_268 == 32'h4 ? _T_91[31:0] : _GEN_385; // @[ivncontrol4.scala 207:50 209:21]
  wire [31:0] _GEN_389 = _GEN_268 == 32'h4 ? _T_91[31:0] : _GEN_386; // @[ivncontrol4.scala 207:50 210:21]
  wire [31:0] _GEN_390 = _GEN_268 == 32'h4 ? _T_91[31:0] : 32'h11; // @[ivncontrol4.scala 125:17 207:50 211:21]
  wire [31:0] _GEN_391 = _GEN_268 == 32'h5 ? _T_91[31:0] : _GEN_387; // @[ivncontrol4.scala 200:50 201:21]
  wire [31:0] _GEN_392 = _GEN_268 == 32'h5 ? _T_91[31:0] : _GEN_388; // @[ivncontrol4.scala 200:50 202:21]
  wire [31:0] _GEN_393 = _GEN_268 == 32'h5 ? _T_91[31:0] : _GEN_389; // @[ivncontrol4.scala 200:50 203:21]
  wire [31:0] _GEN_394 = _GEN_268 == 32'h5 ? _T_91[31:0] : _GEN_390; // @[ivncontrol4.scala 200:50 204:21]
  wire [31:0] _GEN_395 = _GEN_268 == 32'h5 ? _T_91[31:0] : 32'h3; // @[ivncontrol4.scala 126:18 200:50 205:22]
  wire [31:0] _GEN_396 = _GEN_268 == 32'h6 ? _T_91[31:0] : _GEN_391; // @[ivncontrol4.scala 192:52 193:21]
  wire [31:0] _GEN_397 = _GEN_268 == 32'h6 ? _T_91[31:0] : _GEN_392; // @[ivncontrol4.scala 192:52 194:21]
  wire [31:0] _GEN_398 = _GEN_268 == 32'h6 ? _T_91[31:0] : _GEN_393; // @[ivncontrol4.scala 192:52 195:21]
  wire [31:0] _GEN_399 = _GEN_268 == 32'h6 ? _T_91[31:0] : _GEN_394; // @[ivncontrol4.scala 192:52 196:21]
  wire [31:0] _GEN_400 = _GEN_268 == 32'h6 ? _T_91[31:0] : _GEN_395; // @[ivncontrol4.scala 192:52 197:22]
  wire [31:0] _GEN_401 = _GEN_268 == 32'h6 ? _T_91[31:0] : 32'h17; // @[ivncontrol4.scala 126:18 192:52 198:22]
  wire [31:0] _GEN_402 = _GEN_268 == 32'h7 ? _T_91[31:0] : _GEN_396; // @[ivncontrol4.scala 184:52 185:21]
  wire [31:0] _GEN_403 = _GEN_268 == 32'h7 ? _T_91[31:0] : _GEN_397; // @[ivncontrol4.scala 184:52 186:21]
  wire [31:0] _GEN_404 = _GEN_268 == 32'h7 ? _T_91[31:0] : _GEN_398; // @[ivncontrol4.scala 184:52 187:21]
  wire [31:0] _GEN_405 = _GEN_268 == 32'h7 ? _T_91[31:0] : _GEN_399; // @[ivncontrol4.scala 184:52 188:21]
  wire [31:0] _GEN_406 = _GEN_268 == 32'h7 ? _T_91[31:0] : _GEN_400; // @[ivncontrol4.scala 184:52 189:22]
  wire [31:0] _GEN_407 = _GEN_268 == 32'h7 ? _T_91[31:0] : _GEN_401; // @[ivncontrol4.scala 184:52 190:22]
  wire [31:0] _GEN_408 = _GEN_268 == 32'h7 ? _T_91[31:0] : 32'hb; // @[ivncontrol4.scala 126:18 184:52 191:22]
  wire [31:0] _GEN_409 = _GEN_268 >= 32'h8 ? _T_91[31:0] : _GEN_402; // @[ivncontrol4.scala 174:42 175:21]
  wire [31:0] _GEN_410 = _GEN_268 >= 32'h8 ? _T_91[31:0] : _GEN_403; // @[ivncontrol4.scala 174:42 176:21]
  wire [31:0] _GEN_411 = _GEN_268 >= 32'h8 ? _T_91[31:0] : _GEN_404; // @[ivncontrol4.scala 174:42 177:21]
  wire [31:0] _GEN_412 = _GEN_268 >= 32'h8 ? _T_91[31:0] : _GEN_405; // @[ivncontrol4.scala 174:42 178:21]
  wire [31:0] _GEN_413 = _GEN_268 >= 32'h8 ? _T_91[31:0] : _GEN_406; // @[ivncontrol4.scala 174:42 179:22]
  wire [31:0] _GEN_414 = _GEN_268 >= 32'h8 ? _T_91[31:0] : _GEN_407; // @[ivncontrol4.scala 174:42 180:22]
  wire [31:0] _GEN_415 = _GEN_268 >= 32'h8 ? _T_91[31:0] : _GEN_408; // @[ivncontrol4.scala 174:42 181:22]
  wire [31:0] _GEN_416 = _GEN_268 >= 32'h8 ? _T_91[31:0] : 32'h18; // @[ivncontrol4.scala 126:18 174:42 182:22]
  wire [31:0] _T_127 = 32'h8 - _GEN_268; // @[ivncontrol4.scala 228:18]
  wire [31:0] _i_vn_1_T_15 = 32'h1 + pin; // @[ivncontrol4.scala 229:29]
  wire [31:0] _GEN_529 = _T_127 == 32'h1 ? _i_vn_1_T_15 : _GEN_416; // @[ivncontrol4.scala 269:54 272:22]
  wire [31:0] _GEN_530 = _T_127 == 32'h2 ? _i_vn_1_T_15 : _GEN_415; // @[ivncontrol4.scala 264:54 267:22]
  wire [31:0] _GEN_531 = _T_127 == 32'h2 ? _i_vn_1_T_15 : _GEN_529; // @[ivncontrol4.scala 264:54 268:22]
  wire [31:0] _GEN_532 = _T_127 == 32'h3 ? _i_vn_1_T_15 : _GEN_414; // @[ivncontrol4.scala 257:54 259:22]
  wire [31:0] _GEN_533 = _T_127 == 32'h3 ? _i_vn_1_T_15 : _GEN_530; // @[ivncontrol4.scala 257:54 260:22]
  wire [31:0] _GEN_534 = _T_127 == 32'h3 ? _i_vn_1_T_15 : _GEN_531; // @[ivncontrol4.scala 257:54 261:22]
  wire [31:0] _GEN_535 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_413; // @[ivncontrol4.scala 251:54 253:22]
  wire [31:0] _GEN_536 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_532; // @[ivncontrol4.scala 251:54 254:22]
  wire [31:0] _GEN_537 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_533; // @[ivncontrol4.scala 251:54 255:22]
  wire [31:0] _GEN_538 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_534; // @[ivncontrol4.scala 251:54 256:22]
  wire [31:0] _GEN_539 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_412; // @[ivncontrol4.scala 244:54 246:21]
  wire [31:0] _GEN_540 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_535; // @[ivncontrol4.scala 244:54 247:22]
  wire [31:0] _GEN_541 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_536; // @[ivncontrol4.scala 244:54 248:22]
  wire [31:0] _GEN_542 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_537; // @[ivncontrol4.scala 244:54 249:22]
  wire [31:0] _GEN_543 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_538; // @[ivncontrol4.scala 244:54 250:22]
  wire [31:0] _GEN_544 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_411; // @[ivncontrol4.scala 237:54 238:22]
  wire [31:0] _GEN_545 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_539; // @[ivncontrol4.scala 237:54 239:21]
  wire [31:0] _GEN_546 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_540; // @[ivncontrol4.scala 237:54 240:22]
  wire [31:0] _GEN_547 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_541; // @[ivncontrol4.scala 237:54 241:22]
  wire [31:0] _GEN_548 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_542; // @[ivncontrol4.scala 237:54 242:22]
  wire [31:0] _GEN_549 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_543; // @[ivncontrol4.scala 237:54 243:22]
  wire [31:0] _GEN_550 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_410; // @[ivncontrol4.scala 228:49 229:22]
  wire [31:0] _GEN_551 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_544; // @[ivncontrol4.scala 228:49 230:21]
  wire [31:0] _GEN_552 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_545; // @[ivncontrol4.scala 228:49 231:21]
  wire [31:0] _GEN_553 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_546; // @[ivncontrol4.scala 228:49 232:22]
  wire [31:0] _GEN_554 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_547; // @[ivncontrol4.scala 228:49 233:22]
  wire [31:0] _GEN_555 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_548; // @[ivncontrol4.scala 228:49 234:22]
  wire [31:0] _GEN_556 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_549; // @[ivncontrol4.scala 228:49 235:22]
  wire [31:0] _GEN_574 = 4'h1 == _i_vn_1_T_15[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_575 = 4'h2 == _i_vn_1_T_15[3:0] ? rowcount_2 : _GEN_574; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_576 = 4'h3 == _i_vn_1_T_15[3:0] ? rowcount_3 : _GEN_575; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_577 = 4'h4 == _i_vn_1_T_15[3:0] ? rowcount_4 : _GEN_576; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_578 = 4'h5 == _i_vn_1_T_15[3:0] ? rowcount_5 : _GEN_577; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_579 = 4'h6 == _i_vn_1_T_15[3:0] ? rowcount_6 : _GEN_578; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_580 = 4'h7 == _i_vn_1_T_15[3:0] ? rowcount_7 : _GEN_579; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_581 = 4'h8 == _i_vn_1_T_15[3:0] ? rowcount_8 : _GEN_580; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_582 = 4'h9 == _i_vn_1_T_15[3:0] ? rowcount_9 : _GEN_581; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_583 = 4'ha == _i_vn_1_T_15[3:0] ? rowcount_10 : _GEN_582; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_584 = 4'hb == _i_vn_1_T_15[3:0] ? rowcount_11 : _GEN_583; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_585 = 4'hc == _i_vn_1_T_15[3:0] ? rowcount_12 : _GEN_584; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_586 = 4'hd == _i_vn_1_T_15[3:0] ? rowcount_13 : _GEN_585; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_587 = 4'he == _i_vn_1_T_15[3:0] ? rowcount_14 : _GEN_586; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _GEN_588 = 4'hf == _i_vn_1_T_15[3:0] ? rowcount_15 : _GEN_587; // @[ivncontrol4.scala 275:{41,41}]
  wire [31:0] _T_172 = _GEN_268 + _GEN_588; // @[ivncontrol4.scala 275:41]
  wire [31:0] _T_174 = 32'h8 - _T_172; // @[ivncontrol4.scala 275:18]
  wire [31:0] _i_vn_1_T_17 = 32'h2 + pin; // @[ivncontrol4.scala 276:29]
  wire [31:0] _GEN_781 = _T_174 == 32'h1 ? _i_vn_1_T_17 : _GEN_556; // @[ivncontrol4.scala 318:78 321:22]
  wire [31:0] _GEN_782 = _T_174 == 32'h2 ? _i_vn_1_T_17 : _GEN_555; // @[ivncontrol4.scala 312:76 315:22]
  wire [31:0] _GEN_783 = _T_174 == 32'h2 ? _i_vn_1_T_17 : _GEN_781; // @[ivncontrol4.scala 312:76 316:22]
  wire [31:0] _GEN_784 = _T_174 == 32'h3 ? _i_vn_1_T_17 : _GEN_554; // @[ivncontrol4.scala 305:78 307:23]
  wire [31:0] _GEN_785 = _T_174 == 32'h3 ? _i_vn_1_T_17 : _GEN_782; // @[ivncontrol4.scala 305:78 308:22]
  wire [31:0] _GEN_786 = _T_174 == 32'h3 ? _i_vn_1_T_17 : _GEN_783; // @[ivncontrol4.scala 305:78 309:22]
  wire [31:0] _GEN_787 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_553; // @[ivncontrol4.scala 299:78 301:22]
  wire [31:0] _GEN_788 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_784; // @[ivncontrol4.scala 299:78 302:22]
  wire [31:0] _GEN_789 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_785; // @[ivncontrol4.scala 299:78 303:22]
  wire [31:0] _GEN_790 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_786; // @[ivncontrol4.scala 299:78 304:22]
  wire [31:0] _GEN_791 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_552; // @[ivncontrol4.scala 292:76 294:23]
  wire [31:0] _GEN_792 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_787; // @[ivncontrol4.scala 292:76 295:22]
  wire [31:0] _GEN_793 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_788; // @[ivncontrol4.scala 292:76 296:22]
  wire [31:0] _GEN_794 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_789; // @[ivncontrol4.scala 292:76 297:22]
  wire [31:0] _GEN_795 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_790; // @[ivncontrol4.scala 292:76 298:22]
  wire [31:0] _GEN_796 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_551; // @[ivncontrol4.scala 284:77 286:22]
  wire [31:0] _GEN_797 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_791; // @[ivncontrol4.scala 284:77 287:21]
  wire [31:0] _GEN_798 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_792; // @[ivncontrol4.scala 284:77 288:22]
  wire [31:0] _GEN_799 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_793; // @[ivncontrol4.scala 284:77 289:22]
  wire [31:0] _GEN_800 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_794; // @[ivncontrol4.scala 284:77 290:22]
  wire [31:0] _GEN_801 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_795; // @[ivncontrol4.scala 284:77 291:22]
  wire [31:0] _GEN_802 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_550; // @[ivncontrol4.scala 275:73 276:22]
  wire [31:0] _GEN_803 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_796; // @[ivncontrol4.scala 275:73 277:21]
  wire [31:0] _GEN_804 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_797; // @[ivncontrol4.scala 275:73 278:21]
  wire [31:0] _GEN_805 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_798; // @[ivncontrol4.scala 275:73 279:22]
  wire [31:0] _GEN_806 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_799; // @[ivncontrol4.scala 275:73 280:22]
  wire [31:0] _GEN_807 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_800; // @[ivncontrol4.scala 275:73 281:22]
  wire [31:0] _GEN_808 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_801; // @[ivncontrol4.scala 275:73 282:22]
  wire [31:0] _GEN_842 = 4'h1 == _i_vn_1_T_17[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_843 = 4'h2 == _i_vn_1_T_17[3:0] ? rowcount_2 : _GEN_842; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_844 = 4'h3 == _i_vn_1_T_17[3:0] ? rowcount_3 : _GEN_843; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_845 = 4'h4 == _i_vn_1_T_17[3:0] ? rowcount_4 : _GEN_844; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_846 = 4'h5 == _i_vn_1_T_17[3:0] ? rowcount_5 : _GEN_845; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_847 = 4'h6 == _i_vn_1_T_17[3:0] ? rowcount_6 : _GEN_846; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_848 = 4'h7 == _i_vn_1_T_17[3:0] ? rowcount_7 : _GEN_847; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_849 = 4'h8 == _i_vn_1_T_17[3:0] ? rowcount_8 : _GEN_848; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_850 = 4'h9 == _i_vn_1_T_17[3:0] ? rowcount_9 : _GEN_849; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_851 = 4'ha == _i_vn_1_T_17[3:0] ? rowcount_10 : _GEN_850; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_852 = 4'hb == _i_vn_1_T_17[3:0] ? rowcount_11 : _GEN_851; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_853 = 4'hc == _i_vn_1_T_17[3:0] ? rowcount_12 : _GEN_852; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_854 = 4'hd == _i_vn_1_T_17[3:0] ? rowcount_13 : _GEN_853; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_855 = 4'he == _i_vn_1_T_17[3:0] ? rowcount_14 : _GEN_854; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _GEN_856 = 4'hf == _i_vn_1_T_17[3:0] ? rowcount_15 : _GEN_855; // @[ivncontrol4.scala 326:{62,62}]
  wire [31:0] _T_254 = _T_172 + _GEN_856; // @[ivncontrol4.scala 326:62]
  wire [31:0] _T_256 = 32'h8 - _T_254; // @[ivncontrol4.scala 326:17]
  wire [31:0] _i_vn_1_T_19 = 32'h3 + pin; // @[ivncontrol4.scala 327:29]
  wire [31:0] _GEN_1145 = _T_256 == 32'h1 ? _i_vn_1_T_19 : _GEN_808; // @[ivncontrol4.scala 369:100 372:22]
  wire [31:0] _GEN_1146 = _T_256 == 32'h2 ? _i_vn_1_T_19 : _GEN_807; // @[ivncontrol4.scala 363:98 366:22]
  wire [31:0] _GEN_1147 = _T_256 == 32'h2 ? _i_vn_1_T_19 : _GEN_1145; // @[ivncontrol4.scala 363:98 367:22]
  wire [31:0] _GEN_1148 = _T_256 == 32'h3 ? _i_vn_1_T_19 : _GEN_806; // @[ivncontrol4.scala 356:100 358:23]
  wire [31:0] _GEN_1149 = _T_256 == 32'h3 ? _i_vn_1_T_19 : _GEN_1146; // @[ivncontrol4.scala 356:100 359:22]
  wire [31:0] _GEN_1150 = _T_256 == 32'h3 ? _i_vn_1_T_19 : _GEN_1147; // @[ivncontrol4.scala 356:100 360:22]
  wire [31:0] _GEN_1151 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_805; // @[ivncontrol4.scala 350:100 352:22]
  wire [31:0] _GEN_1152 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_1148; // @[ivncontrol4.scala 350:100 353:22]
  wire [31:0] _GEN_1153 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_1149; // @[ivncontrol4.scala 350:100 354:22]
  wire [31:0] _GEN_1154 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_1150; // @[ivncontrol4.scala 350:100 355:22]
  wire [31:0] _GEN_1155 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_804; // @[ivncontrol4.scala 343:98 345:23]
  wire [31:0] _GEN_1156 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1151; // @[ivncontrol4.scala 343:98 346:22]
  wire [31:0] _GEN_1157 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1152; // @[ivncontrol4.scala 343:98 347:22]
  wire [31:0] _GEN_1158 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1153; // @[ivncontrol4.scala 343:98 348:22]
  wire [31:0] _GEN_1159 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1154; // @[ivncontrol4.scala 343:98 349:22]
  wire [31:0] _GEN_1160 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_803; // @[ivncontrol4.scala 335:99 337:22]
  wire [31:0] _GEN_1161 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1155; // @[ivncontrol4.scala 335:99 338:21]
  wire [31:0] _GEN_1162 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1156; // @[ivncontrol4.scala 335:99 339:22]
  wire [31:0] _GEN_1163 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1157; // @[ivncontrol4.scala 335:99 340:22]
  wire [31:0] _GEN_1164 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1158; // @[ivncontrol4.scala 335:99 341:22]
  wire [31:0] _GEN_1165 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1159; // @[ivncontrol4.scala 335:99 342:22]
  wire [31:0] _GEN_1166 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_802; // @[ivncontrol4.scala 326:94 327:22]
  wire [31:0] _GEN_1167 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1160; // @[ivncontrol4.scala 326:94 328:21]
  wire [31:0] _GEN_1168 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1161; // @[ivncontrol4.scala 326:94 329:21]
  wire [31:0] _GEN_1169 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1162; // @[ivncontrol4.scala 326:94 330:22]
  wire [31:0] _GEN_1170 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1163; // @[ivncontrol4.scala 326:94 331:22]
  wire [31:0] _GEN_1171 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1164; // @[ivncontrol4.scala 326:94 332:22]
  wire [31:0] _GEN_1172 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1165; // @[ivncontrol4.scala 326:94 333:22]
  wire [31:0] _GEN_1222 = 4'h1 == _i_vn_1_T_19[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1223 = 4'h2 == _i_vn_1_T_19[3:0] ? rowcount_2 : _GEN_1222; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1224 = 4'h3 == _i_vn_1_T_19[3:0] ? rowcount_3 : _GEN_1223; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1225 = 4'h4 == _i_vn_1_T_19[3:0] ? rowcount_4 : _GEN_1224; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1226 = 4'h5 == _i_vn_1_T_19[3:0] ? rowcount_5 : _GEN_1225; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1227 = 4'h6 == _i_vn_1_T_19[3:0] ? rowcount_6 : _GEN_1226; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1228 = 4'h7 == _i_vn_1_T_19[3:0] ? rowcount_7 : _GEN_1227; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1229 = 4'h8 == _i_vn_1_T_19[3:0] ? rowcount_8 : _GEN_1228; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1230 = 4'h9 == _i_vn_1_T_19[3:0] ? rowcount_9 : _GEN_1229; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1231 = 4'ha == _i_vn_1_T_19[3:0] ? rowcount_10 : _GEN_1230; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1232 = 4'hb == _i_vn_1_T_19[3:0] ? rowcount_11 : _GEN_1231; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1233 = 4'hc == _i_vn_1_T_19[3:0] ? rowcount_12 : _GEN_1232; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1234 = 4'hd == _i_vn_1_T_19[3:0] ? rowcount_13 : _GEN_1233; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1235 = 4'he == _i_vn_1_T_19[3:0] ? rowcount_14 : _GEN_1234; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _GEN_1236 = 4'hf == _i_vn_1_T_19[3:0] ? rowcount_15 : _GEN_1235; // @[ivncontrol4.scala 376:{86,86}]
  wire [31:0] _T_371 = _T_254 + _GEN_1236; // @[ivncontrol4.scala 376:86]
  wire [31:0] _T_373 = 32'h8 - _T_371; // @[ivncontrol4.scala 376:19]
  wire [31:0] _i_vn_1_T_21 = 32'h4 + pin; // @[ivncontrol4.scala 377:29]
  wire [31:0] _GEN_1621 = _T_373 == 32'h1 ? _i_vn_1_T_21 : _GEN_1172; // @[ivncontrol4.scala 419:122 422:22]
  wire [31:0] _GEN_1622 = _T_373 == 32'h2 ? _i_vn_1_T_21 : _GEN_1171; // @[ivncontrol4.scala 413:121 416:22]
  wire [31:0] _GEN_1623 = _T_373 == 32'h2 ? _i_vn_1_T_21 : _GEN_1621; // @[ivncontrol4.scala 413:121 417:22]
  wire [31:0] _GEN_1624 = _T_373 == 32'h3 ? _i_vn_1_T_21 : _GEN_1170; // @[ivncontrol4.scala 406:123 408:23]
  wire [31:0] _GEN_1625 = _T_373 == 32'h3 ? _i_vn_1_T_21 : _GEN_1622; // @[ivncontrol4.scala 406:123 409:22]
  wire [31:0] _GEN_1626 = _T_373 == 32'h3 ? _i_vn_1_T_21 : _GEN_1623; // @[ivncontrol4.scala 406:123 410:22]
  wire [31:0] _GEN_1627 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1169; // @[ivncontrol4.scala 400:122 402:22]
  wire [31:0] _GEN_1628 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1624; // @[ivncontrol4.scala 400:122 403:22]
  wire [31:0] _GEN_1629 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1625; // @[ivncontrol4.scala 400:122 404:22]
  wire [31:0] _GEN_1630 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1626; // @[ivncontrol4.scala 400:122 405:22]
  wire [31:0] _GEN_1631 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1168; // @[ivncontrol4.scala 393:121 395:23]
  wire [31:0] _GEN_1632 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1627; // @[ivncontrol4.scala 393:121 396:22]
  wire [31:0] _GEN_1633 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1628; // @[ivncontrol4.scala 393:121 397:22]
  wire [31:0] _GEN_1634 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1629; // @[ivncontrol4.scala 393:121 398:22]
  wire [31:0] _GEN_1635 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1630; // @[ivncontrol4.scala 393:121 399:22]
  wire [31:0] _GEN_1636 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1167; // @[ivncontrol4.scala 385:121 387:22]
  wire [31:0] _GEN_1637 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1631; // @[ivncontrol4.scala 385:121 388:21]
  wire [31:0] _GEN_1638 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1632; // @[ivncontrol4.scala 385:121 389:22]
  wire [31:0] _GEN_1639 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1633; // @[ivncontrol4.scala 385:121 390:22]
  wire [31:0] _GEN_1640 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1634; // @[ivncontrol4.scala 385:121 391:22]
  wire [31:0] _GEN_1641 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1635; // @[ivncontrol4.scala 385:121 392:22]
  wire [31:0] _GEN_1642 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1166; // @[ivncontrol4.scala 376:118 377:22]
  wire [31:0] _GEN_1643 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1636; // @[ivncontrol4.scala 376:118 378:21]
  wire [31:0] _GEN_1644 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1637; // @[ivncontrol4.scala 376:118 379:21]
  wire [31:0] _GEN_1645 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1638; // @[ivncontrol4.scala 376:118 380:22]
  wire [31:0] _GEN_1646 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1639; // @[ivncontrol4.scala 376:118 381:22]
  wire [31:0] _GEN_1647 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1640; // @[ivncontrol4.scala 376:118 382:22]
  wire [31:0] _GEN_1648 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1641; // @[ivncontrol4.scala 376:118 383:22]
  wire [31:0] _GEN_1714 = 4'h1 == _i_vn_1_T_21[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1715 = 4'h2 == _i_vn_1_T_21[3:0] ? rowcount_2 : _GEN_1714; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1716 = 4'h3 == _i_vn_1_T_21[3:0] ? rowcount_3 : _GEN_1715; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1717 = 4'h4 == _i_vn_1_T_21[3:0] ? rowcount_4 : _GEN_1716; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1718 = 4'h5 == _i_vn_1_T_21[3:0] ? rowcount_5 : _GEN_1717; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1719 = 4'h6 == _i_vn_1_T_21[3:0] ? rowcount_6 : _GEN_1718; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1720 = 4'h7 == _i_vn_1_T_21[3:0] ? rowcount_7 : _GEN_1719; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1721 = 4'h8 == _i_vn_1_T_21[3:0] ? rowcount_8 : _GEN_1720; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1722 = 4'h9 == _i_vn_1_T_21[3:0] ? rowcount_9 : _GEN_1721; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1723 = 4'ha == _i_vn_1_T_21[3:0] ? rowcount_10 : _GEN_1722; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1724 = 4'hb == _i_vn_1_T_21[3:0] ? rowcount_11 : _GEN_1723; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1725 = 4'hc == _i_vn_1_T_21[3:0] ? rowcount_12 : _GEN_1724; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1726 = 4'hd == _i_vn_1_T_21[3:0] ? rowcount_13 : _GEN_1725; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1727 = 4'he == _i_vn_1_T_21[3:0] ? rowcount_14 : _GEN_1726; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _GEN_1728 = 4'hf == _i_vn_1_T_21[3:0] ? rowcount_15 : _GEN_1727; // @[ivncontrol4.scala 426:{108,108}]
  wire [31:0] _T_523 = _T_371 + _GEN_1728; // @[ivncontrol4.scala 426:108]
  wire [31:0] _T_525 = 32'h8 - _T_523; // @[ivncontrol4.scala 426:19]
  wire [31:0] _i_vn_1_T_23 = 32'h5 + pin; // @[ivncontrol4.scala 427:29]
  wire [31:0] _GEN_2209 = _T_525 == 32'h1 ? _i_vn_1_T_23 : _GEN_1648; // @[ivncontrol4.scala 469:144 472:22]
  wire [31:0] _GEN_2210 = _T_525 == 32'h2 ? _i_vn_1_T_23 : _GEN_1647; // @[ivncontrol4.scala 463:143 466:22]
  wire [31:0] _GEN_2211 = _T_525 == 32'h2 ? _i_vn_1_T_23 : _GEN_2209; // @[ivncontrol4.scala 463:143 467:22]
  wire [31:0] _GEN_2212 = _T_525 == 32'h3 ? _i_vn_1_T_23 : _GEN_1646; // @[ivncontrol4.scala 456:145 458:23]
  wire [31:0] _GEN_2213 = _T_525 == 32'h3 ? _i_vn_1_T_23 : _GEN_2210; // @[ivncontrol4.scala 456:145 459:22]
  wire [31:0] _GEN_2214 = _T_525 == 32'h3 ? _i_vn_1_T_23 : _GEN_2211; // @[ivncontrol4.scala 456:145 460:22]
  wire [31:0] _GEN_2215 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_1645; // @[ivncontrol4.scala 450:143 452:22]
  wire [31:0] _GEN_2216 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_2212; // @[ivncontrol4.scala 450:143 453:22]
  wire [31:0] _GEN_2217 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_2213; // @[ivncontrol4.scala 450:143 454:22]
  wire [31:0] _GEN_2218 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_2214; // @[ivncontrol4.scala 450:143 455:22]
  wire [31:0] _GEN_2219 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_1644; // @[ivncontrol4.scala 443:143 445:23]
  wire [31:0] _GEN_2220 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2215; // @[ivncontrol4.scala 443:143 446:22]
  wire [31:0] _GEN_2221 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2216; // @[ivncontrol4.scala 443:143 447:22]
  wire [31:0] _GEN_2222 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2217; // @[ivncontrol4.scala 443:143 448:22]
  wire [31:0] _GEN_2223 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2218; // @[ivncontrol4.scala 443:143 449:22]
  wire [31:0] _GEN_2224 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_1643; // @[ivncontrol4.scala 435:143 437:22]
  wire [31:0] _GEN_2225 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2219; // @[ivncontrol4.scala 435:143 438:21]
  wire [31:0] _GEN_2226 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2220; // @[ivncontrol4.scala 435:143 439:22]
  wire [31:0] _GEN_2227 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2221; // @[ivncontrol4.scala 435:143 440:22]
  wire [31:0] _GEN_2228 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2222; // @[ivncontrol4.scala 435:143 441:22]
  wire [31:0] _GEN_2229 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2223; // @[ivncontrol4.scala 435:143 442:22]
  wire [31:0] _GEN_2230 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_1642; // @[ivncontrol4.scala 426:140 427:22]
  wire [31:0] _GEN_2231 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2224; // @[ivncontrol4.scala 426:140 428:21]
  wire [31:0] _GEN_2232 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2225; // @[ivncontrol4.scala 426:140 429:21]
  wire [31:0] _GEN_2233 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2226; // @[ivncontrol4.scala 426:140 430:22]
  wire [31:0] _GEN_2234 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2227; // @[ivncontrol4.scala 426:140 431:22]
  wire [31:0] _GEN_2235 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2228; // @[ivncontrol4.scala 426:140 432:22]
  wire [31:0] _GEN_2236 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2229; // @[ivncontrol4.scala 426:140 433:22]
  wire [31:0] _GEN_2318 = 4'h1 == _i_vn_1_T_23[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2319 = 4'h2 == _i_vn_1_T_23[3:0] ? rowcount_2 : _GEN_2318; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2320 = 4'h3 == _i_vn_1_T_23[3:0] ? rowcount_3 : _GEN_2319; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2321 = 4'h4 == _i_vn_1_T_23[3:0] ? rowcount_4 : _GEN_2320; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2322 = 4'h5 == _i_vn_1_T_23[3:0] ? rowcount_5 : _GEN_2321; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2323 = 4'h6 == _i_vn_1_T_23[3:0] ? rowcount_6 : _GEN_2322; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2324 = 4'h7 == _i_vn_1_T_23[3:0] ? rowcount_7 : _GEN_2323; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2325 = 4'h8 == _i_vn_1_T_23[3:0] ? rowcount_8 : _GEN_2324; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2326 = 4'h9 == _i_vn_1_T_23[3:0] ? rowcount_9 : _GEN_2325; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2327 = 4'ha == _i_vn_1_T_23[3:0] ? rowcount_10 : _GEN_2326; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2328 = 4'hb == _i_vn_1_T_23[3:0] ? rowcount_11 : _GEN_2327; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2329 = 4'hc == _i_vn_1_T_23[3:0] ? rowcount_12 : _GEN_2328; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2330 = 4'hd == _i_vn_1_T_23[3:0] ? rowcount_13 : _GEN_2329; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2331 = 4'he == _i_vn_1_T_23[3:0] ? rowcount_14 : _GEN_2330; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _GEN_2332 = 4'hf == _i_vn_1_T_23[3:0] ? rowcount_15 : _GEN_2331; // @[ivncontrol4.scala 477:{130,130}]
  wire [31:0] _T_710 = _T_523 + _GEN_2332; // @[ivncontrol4.scala 477:130]
  wire [31:0] _T_712 = 32'h8 - _T_710; // @[ivncontrol4.scala 477:19]
  wire [31:0] _i_vn_1_T_25 = 32'h6 + pin; // @[ivncontrol4.scala 478:29]
  wire [31:0] _GEN_2909 = _T_712 == 32'h1 ? _i_vn_1_T_25 : _GEN_2236; // @[ivncontrol4.scala 520:166 523:22]
  wire [31:0] _GEN_2910 = _T_712 == 32'h2 ? _i_vn_1_T_25 : _GEN_2235; // @[ivncontrol4.scala 514:166 517:22]
  wire [31:0] _GEN_2911 = _T_712 == 32'h2 ? _i_vn_1_T_25 : _GEN_2909; // @[ivncontrol4.scala 514:166 518:22]
  wire [31:0] _GEN_2912 = _T_712 == 32'h3 ? _i_vn_1_T_25 : _GEN_2234; // @[ivncontrol4.scala 507:168 509:23]
  wire [31:0] _GEN_2913 = _T_712 == 32'h3 ? _i_vn_1_T_25 : _GEN_2910; // @[ivncontrol4.scala 507:168 510:22]
  wire [31:0] _GEN_2914 = _T_712 == 32'h3 ? _i_vn_1_T_25 : _GEN_2911; // @[ivncontrol4.scala 507:168 511:22]
  wire [31:0] _GEN_2915 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2233; // @[ivncontrol4.scala 501:166 503:22]
  wire [31:0] _GEN_2916 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2912; // @[ivncontrol4.scala 501:166 504:22]
  wire [31:0] _GEN_2917 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2913; // @[ivncontrol4.scala 501:166 505:22]
  wire [31:0] _GEN_2918 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2914; // @[ivncontrol4.scala 501:166 506:22]
  wire [31:0] _GEN_2919 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2232; // @[ivncontrol4.scala 494:166 496:23]
  wire [31:0] _GEN_2920 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2915; // @[ivncontrol4.scala 494:166 497:22]
  wire [31:0] _GEN_2921 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2916; // @[ivncontrol4.scala 494:166 498:22]
  wire [31:0] _GEN_2922 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2917; // @[ivncontrol4.scala 494:166 499:22]
  wire [31:0] _GEN_2923 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2918; // @[ivncontrol4.scala 494:166 500:22]
  wire [31:0] _GEN_2924 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2231; // @[ivncontrol4.scala 486:166 488:22]
  wire [31:0] _GEN_2925 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2919; // @[ivncontrol4.scala 486:166 489:21]
  wire [31:0] _GEN_2926 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2920; // @[ivncontrol4.scala 486:166 490:22]
  wire [31:0] _GEN_2927 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2921; // @[ivncontrol4.scala 486:166 491:22]
  wire [31:0] _GEN_2928 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2922; // @[ivncontrol4.scala 486:166 492:22]
  wire [31:0] _GEN_2929 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2923; // @[ivncontrol4.scala 486:166 493:22]
  wire [31:0] _GEN_2930 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2230; // @[ivncontrol4.scala 477:162 478:22]
  wire [31:0] _GEN_2931 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2924; // @[ivncontrol4.scala 477:162 479:21]
  wire [31:0] _GEN_2932 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2925; // @[ivncontrol4.scala 477:162 480:21]
  wire [31:0] _GEN_2933 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2926; // @[ivncontrol4.scala 477:162 481:22]
  wire [31:0] _GEN_2934 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2927; // @[ivncontrol4.scala 477:162 482:22]
  wire [31:0] _GEN_2935 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2928; // @[ivncontrol4.scala 477:162 483:22]
  wire [31:0] _GEN_2936 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2929; // @[ivncontrol4.scala 477:162 484:22]
  wire [31:0] _GEN_3034 = 4'h1 == _i_vn_1_T_25[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3035 = 4'h2 == _i_vn_1_T_25[3:0] ? rowcount_2 : _GEN_3034; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3036 = 4'h3 == _i_vn_1_T_25[3:0] ? rowcount_3 : _GEN_3035; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3037 = 4'h4 == _i_vn_1_T_25[3:0] ? rowcount_4 : _GEN_3036; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3038 = 4'h5 == _i_vn_1_T_25[3:0] ? rowcount_5 : _GEN_3037; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3039 = 4'h6 == _i_vn_1_T_25[3:0] ? rowcount_6 : _GEN_3038; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3040 = 4'h7 == _i_vn_1_T_25[3:0] ? rowcount_7 : _GEN_3039; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3041 = 4'h8 == _i_vn_1_T_25[3:0] ? rowcount_8 : _GEN_3040; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3042 = 4'h9 == _i_vn_1_T_25[3:0] ? rowcount_9 : _GEN_3041; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3043 = 4'ha == _i_vn_1_T_25[3:0] ? rowcount_10 : _GEN_3042; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3044 = 4'hb == _i_vn_1_T_25[3:0] ? rowcount_11 : _GEN_3043; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3045 = 4'hc == _i_vn_1_T_25[3:0] ? rowcount_12 : _GEN_3044; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3046 = 4'hd == _i_vn_1_T_25[3:0] ? rowcount_13 : _GEN_3045; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3047 = 4'he == _i_vn_1_T_25[3:0] ? rowcount_14 : _GEN_3046; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _GEN_3048 = 4'hf == _i_vn_1_T_25[3:0] ? rowcount_15 : _GEN_3047; // @[ivncontrol4.scala 528:{152,152}]
  wire [31:0] _T_932 = _T_710 + _GEN_3048; // @[ivncontrol4.scala 528:152]
  wire [31:0] _T_934 = 32'h8 - _T_932; // @[ivncontrol4.scala 528:19]
  wire [31:0] _i_vn_1_T_27 = 32'h7 + pin; // @[ivncontrol4.scala 529:29]
  wire [31:0] _GEN_3721 = _T_934 == 32'h1 ? _i_vn_1_T_27 : _GEN_2936; // @[ivncontrol4.scala 571:188 574:22]
  wire [31:0] _GEN_3722 = _T_934 == 32'h2 ? _i_vn_1_T_27 : _GEN_2935; // @[ivncontrol4.scala 565:188 568:22]
  wire [31:0] _GEN_3723 = _T_934 == 32'h2 ? _i_vn_1_T_27 : _GEN_3721; // @[ivncontrol4.scala 565:188 569:22]
  wire [31:0] _GEN_3724 = _T_934 == 32'h3 ? _i_vn_1_T_27 : _GEN_2934; // @[ivncontrol4.scala 558:190 560:23]
  wire [31:0] _GEN_3725 = _T_934 == 32'h3 ? _i_vn_1_T_27 : _GEN_3722; // @[ivncontrol4.scala 558:190 561:22]
  wire [31:0] _GEN_3726 = _T_934 == 32'h3 ? _i_vn_1_T_27 : _GEN_3723; // @[ivncontrol4.scala 558:190 562:22]
  wire [31:0] _GEN_3727 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_2933; // @[ivncontrol4.scala 552:188 554:22]
  wire [31:0] _GEN_3728 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_3724; // @[ivncontrol4.scala 552:188 555:22]
  wire [31:0] _GEN_3729 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_3725; // @[ivncontrol4.scala 552:188 556:22]
  wire [31:0] _GEN_3730 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_3726; // @[ivncontrol4.scala 552:188 557:22]
  wire [31:0] _GEN_3731 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_2932; // @[ivncontrol4.scala 545:188 547:23]
  wire [31:0] _GEN_3732 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3727; // @[ivncontrol4.scala 545:188 548:22]
  wire [31:0] _GEN_3733 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3728; // @[ivncontrol4.scala 545:188 549:22]
  wire [31:0] _GEN_3734 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3729; // @[ivncontrol4.scala 545:188 550:22]
  wire [31:0] _GEN_3735 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3730; // @[ivncontrol4.scala 545:188 551:22]
  wire [31:0] _GEN_3736 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_2931; // @[ivncontrol4.scala 537:188 539:22]
  wire [31:0] _GEN_3737 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3731; // @[ivncontrol4.scala 537:188 540:21]
  wire [31:0] _GEN_3738 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3732; // @[ivncontrol4.scala 537:188 541:22]
  wire [31:0] _GEN_3739 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3733; // @[ivncontrol4.scala 537:188 542:22]
  wire [31:0] _GEN_3740 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3734; // @[ivncontrol4.scala 537:188 543:22]
  wire [31:0] _GEN_3741 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3735; // @[ivncontrol4.scala 537:188 544:22]
  wire [31:0] _GEN_3742 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_2930; // @[ivncontrol4.scala 528:184 529:22]
  wire [31:0] _GEN_3743 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3736; // @[ivncontrol4.scala 528:184 530:21]
  wire [31:0] _GEN_3744 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3737; // @[ivncontrol4.scala 528:184 531:21]
  wire [31:0] _GEN_3745 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3738; // @[ivncontrol4.scala 528:184 532:22]
  wire [31:0] _GEN_3746 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3739; // @[ivncontrol4.scala 528:184 533:22]
  wire [31:0] _GEN_3747 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3740; // @[ivncontrol4.scala 528:184 534:22]
  wire [31:0] _GEN_3748 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3741; // @[ivncontrol4.scala 528:184 535:22]
  wire [31:0] _GEN_3749 = _GEN_244 ? _GEN_409 : 32'h1d; // @[ivncontrol4.scala 125:17 172:28]
  wire [31:0] _GEN_3750 = _GEN_244 ? _GEN_3742 : 32'h0; // @[ivncontrol4.scala 125:17 172:28]
  wire [31:0] _GEN_3751 = _GEN_244 ? _GEN_3743 : 32'h17; // @[ivncontrol4.scala 125:17 172:28]
  wire [31:0] _GEN_3752 = _GEN_244 ? _GEN_3744 : 32'h11; // @[ivncontrol4.scala 125:17 172:28]
  wire [31:0] _GEN_3753 = _GEN_244 ? _GEN_3745 : 32'h3; // @[ivncontrol4.scala 126:18 172:28]
  wire [31:0] _GEN_3754 = _GEN_244 ? _GEN_3746 : 32'h17; // @[ivncontrol4.scala 126:18 172:28]
  wire [31:0] _GEN_3755 = _GEN_244 ? _GEN_3747 : 32'hb; // @[ivncontrol4.scala 126:18 172:28]
  wire [31:0] _GEN_3756 = _GEN_244 ? _GEN_3748 : 32'h18; // @[ivncontrol4.scala 126:18 172:28]
  wire [31:0] _GEN_4137 = reset ? 32'h0 : _GEN_3749; // @[ivncontrol4.scala 16:{23,23}]
  wire [31:0] _GEN_4138 = reset ? 32'h0 : _GEN_3750; // @[ivncontrol4.scala 16:{23,23}]
  wire [31:0] _GEN_4139 = reset ? 32'h0 : _GEN_3751; // @[ivncontrol4.scala 16:{23,23}]
  wire [31:0] _GEN_4140 = reset ? 32'h0 : _GEN_3752; // @[ivncontrol4.scala 16:{23,23}]
  wire [31:0] _GEN_4141 = reset ? 32'h0 : _GEN_3753; // @[ivncontrol4.scala 17:{24,24}]
  wire [31:0] _GEN_4142 = reset ? 32'h0 : _GEN_3754; // @[ivncontrol4.scala 17:{24,24}]
  wire [31:0] _GEN_4143 = reset ? 32'h0 : _GEN_3755; // @[ivncontrol4.scala 17:{24,24}]
  wire [31:0] _GEN_4144 = reset ? 32'h0 : _GEN_3756; // @[ivncontrol4.scala 17:{24,24}]
  assign io_o_vn_0 = i_vn_0; // @[ivncontrol4.scala 121:13]
  assign io_o_vn_1 = i_vn_1; // @[ivncontrol4.scala 121:13]
  assign io_o_vn_2 = i_vn_2; // @[ivncontrol4.scala 121:13]
  assign io_o_vn_3 = i_vn_3; // @[ivncontrol4.scala 121:13]
  assign io_o_vn2_0 = i_vn2_0; // @[ivncontrol4.scala 122:14]
  assign io_o_vn2_1 = i_vn2_1; // @[ivncontrol4.scala 122:14]
  assign io_o_vn2_2 = i_vn2_2; // @[ivncontrol4.scala 122:14]
  assign io_o_vn2_3 = i_vn2_3; // @[ivncontrol4.scala 122:14]
  always @(posedge clock) begin
    i_vn_0 <= _GEN_4137[4:0]; // @[ivncontrol4.scala 16:{23,23}]
    i_vn_1 <= _GEN_4138[4:0]; // @[ivncontrol4.scala 16:{23,23}]
    i_vn_2 <= _GEN_4139[4:0]; // @[ivncontrol4.scala 16:{23,23}]
    i_vn_3 <= _GEN_4140[4:0]; // @[ivncontrol4.scala 16:{23,23}]
    i_vn2_0 <= _GEN_4141[4:0]; // @[ivncontrol4.scala 17:{24,24}]
    i_vn2_1 <= _GEN_4142[4:0]; // @[ivncontrol4.scala 17:{24,24}]
    i_vn2_2 <= _GEN_4143[4:0]; // @[ivncontrol4.scala 17:{24,24}]
    i_vn2_3 <= _GEN_4144[4:0]; // @[ivncontrol4.scala 17:{24,24}]
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_0 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_0 <= count_0; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_1 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_1 <= count_1; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_2 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_2 <= count_2; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_3 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_3 <= count_3; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_4 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_4 <= count_4; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_5 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_5 <= count_5; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_6 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_6 <= count_6; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_7 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_7 <= count_7; // @[ivncontrol4.scala 79:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_8 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_8 <= 32'h0; // @[ivncontrol4.scala 81:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_9 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_9 <= 32'h0; // @[ivncontrol4.scala 81:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_10 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_10 <= 32'h0; // @[ivncontrol4.scala 81:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_11 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_11 <= 32'h0; // @[ivncontrol4.scala 81:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_12 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_12 <= 32'h0; // @[ivncontrol4.scala 81:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_13 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_13 <= 32'h0; // @[ivncontrol4.scala 81:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_14 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end else if (_k_T_2) begin // @[ivncontrol4.scala 72:75]
      rowcount_14 <= 32'h0; // @[ivncontrol4.scala 81:19]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      rowcount_15 <= 32'h0; // @[ivncontrol4.scala 21:27]
    end
    if (reset) begin // @[ivncontrol4.scala 31:22]
      pin <= 32'h0; // @[ivncontrol4.scala 31:22]
    end else if (_T_72 & rowcount_6 == 32'h0 & rowcount_7 != 32'h0) begin // @[ivncontrol4.scala 166:192]
      pin <= 32'h7; // @[ivncontrol4.scala 167:13]
    end else if (_T_59 & rowcount_5 == 32'h0 & rowcount_6 != 32'h0) begin // @[ivncontrol4.scala 163:169]
      pin <= 32'h6; // @[ivncontrol4.scala 164:13]
    end else if (_T_48 & rowcount_4 == 32'h0 & rowcount_5 != 32'h0) begin // @[ivncontrol4.scala 160:146]
      pin <= 32'h5; // @[ivncontrol4.scala 161:13]
    end else begin
      pin <= _GEN_249;
    end
    if (reset) begin // @[ivncontrol4.scala 35:20]
      i <= 32'h0; // @[ivncontrol4.scala 35:20]
    end else if (i < 32'h7 & _k_T_1) begin // @[ivncontrol4.scala 103:74]
      i <= _i_T_1; // @[ivncontrol4.scala 104:11]
    end
    if (reset) begin // @[ivncontrol4.scala 36:20]
      j <= 32'h0; // @[ivncontrol4.scala 36:20]
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 107:71]
      j <= _j_T_1; // @[ivncontrol4.scala 108:11]
    end else if (!(_k_T_2)) begin // @[ivncontrol4.scala 110:81]
      j <= 32'h0; // @[ivncontrol4.scala 114:11]
    end
    if (3'h0 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h0 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h0 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h0 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h0 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h0 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h0 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h0 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_0_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h1 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_1_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h2 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_2_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h3 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_3_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h4 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_4_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h5 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_5_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h6 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_6_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_0 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_1 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_2 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_3 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_4 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_5 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_6 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 57:15]
      mat_7_7 <= _mat_T_3_T_4; // @[ivncontrol4.scala 57:15]
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h0 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_0 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h1 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_1 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h2 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_2 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h3 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_3 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h4 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_4 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h5 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_5 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h6 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_6 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
    if (~_GEN_225) begin // @[ivncontrol4.scala 58:28]
      if (_GEN_128 != 16'h0) begin // @[ivncontrol4.scala 59:51]
        if (3'h7 == i[2:0]) begin // @[ivncontrol4.scala 60:22]
          count_7 <= _count_T_2; // @[ivncontrol4.scala 60:22]
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  i_vn_0 = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  i_vn_1 = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  i_vn_2 = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  i_vn_3 = _RAND_3[4:0];
  _RAND_4 = {1{`RANDOM}};
  i_vn2_0 = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  i_vn2_1 = _RAND_5[4:0];
  _RAND_6 = {1{`RANDOM}};
  i_vn2_2 = _RAND_6[4:0];
  _RAND_7 = {1{`RANDOM}};
  i_vn2_3 = _RAND_7[4:0];
  _RAND_8 = {1{`RANDOM}};
  rowcount_0 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  rowcount_1 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  rowcount_2 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  rowcount_3 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  rowcount_4 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  rowcount_5 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  rowcount_6 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  rowcount_7 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  rowcount_8 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  rowcount_9 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  rowcount_10 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  rowcount_11 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  rowcount_12 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  rowcount_13 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  rowcount_14 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  rowcount_15 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  pin = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  i = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  j = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  mat_0_0 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  mat_0_1 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  mat_0_2 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  mat_0_3 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  mat_0_4 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  mat_0_5 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  mat_0_6 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  mat_0_7 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  mat_1_0 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  mat_1_1 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  mat_1_2 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  mat_1_3 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  mat_1_4 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  mat_1_5 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  mat_1_6 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  mat_1_7 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  mat_2_0 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  mat_2_1 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  mat_2_2 = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  mat_2_3 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  mat_2_4 = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  mat_2_5 = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  mat_2_6 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  mat_2_7 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  mat_3_0 = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  mat_3_1 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  mat_3_2 = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  mat_3_3 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  mat_3_4 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  mat_3_5 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  mat_3_6 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  mat_3_7 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  mat_4_0 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  mat_4_1 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  mat_4_2 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  mat_4_3 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  mat_4_4 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  mat_4_5 = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  mat_4_6 = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  mat_4_7 = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  mat_5_0 = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  mat_5_1 = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  mat_5_2 = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  mat_5_3 = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  mat_5_4 = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  mat_5_5 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  mat_5_6 = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  mat_5_7 = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  mat_6_0 = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  mat_6_1 = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  mat_6_2 = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  mat_6_3 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  mat_6_4 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  mat_6_5 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  mat_6_6 = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  mat_6_7 = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  mat_7_0 = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  mat_7_1 = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  mat_7_2 = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  mat_7_3 = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  mat_7_4 = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  mat_7_5 = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  mat_7_6 = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  mat_7_7 = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  count_0 = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  count_1 = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  count_2 = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  count_3 = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  count_4 = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  count_5 = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  count_6 = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  count_7 = _RAND_98[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ivntop(
  input         clock,
  input         reset,
  output        io_ProcessValid,
  input  [15:0] io_Stationary_matrix_0_0,
  input  [15:0] io_Stationary_matrix_0_1,
  input  [15:0] io_Stationary_matrix_0_2,
  input  [15:0] io_Stationary_matrix_0_3,
  input  [15:0] io_Stationary_matrix_0_4,
  input  [15:0] io_Stationary_matrix_0_5,
  input  [15:0] io_Stationary_matrix_0_6,
  input  [15:0] io_Stationary_matrix_0_7,
  input  [15:0] io_Stationary_matrix_1_0,
  input  [15:0] io_Stationary_matrix_1_1,
  input  [15:0] io_Stationary_matrix_1_2,
  input  [15:0] io_Stationary_matrix_1_3,
  input  [15:0] io_Stationary_matrix_1_4,
  input  [15:0] io_Stationary_matrix_1_5,
  input  [15:0] io_Stationary_matrix_1_6,
  input  [15:0] io_Stationary_matrix_1_7,
  input  [15:0] io_Stationary_matrix_2_0,
  input  [15:0] io_Stationary_matrix_2_1,
  input  [15:0] io_Stationary_matrix_2_2,
  input  [15:0] io_Stationary_matrix_2_3,
  input  [15:0] io_Stationary_matrix_2_4,
  input  [15:0] io_Stationary_matrix_2_5,
  input  [15:0] io_Stationary_matrix_2_6,
  input  [15:0] io_Stationary_matrix_2_7,
  input  [15:0] io_Stationary_matrix_3_0,
  input  [15:0] io_Stationary_matrix_3_1,
  input  [15:0] io_Stationary_matrix_3_2,
  input  [15:0] io_Stationary_matrix_3_3,
  input  [15:0] io_Stationary_matrix_3_4,
  input  [15:0] io_Stationary_matrix_3_5,
  input  [15:0] io_Stationary_matrix_3_6,
  input  [15:0] io_Stationary_matrix_3_7,
  input  [15:0] io_Stationary_matrix_4_0,
  input  [15:0] io_Stationary_matrix_4_1,
  input  [15:0] io_Stationary_matrix_4_2,
  input  [15:0] io_Stationary_matrix_4_3,
  input  [15:0] io_Stationary_matrix_4_4,
  input  [15:0] io_Stationary_matrix_4_5,
  input  [15:0] io_Stationary_matrix_4_6,
  input  [15:0] io_Stationary_matrix_4_7,
  input  [15:0] io_Stationary_matrix_5_0,
  input  [15:0] io_Stationary_matrix_5_1,
  input  [15:0] io_Stationary_matrix_5_2,
  input  [15:0] io_Stationary_matrix_5_3,
  input  [15:0] io_Stationary_matrix_5_4,
  input  [15:0] io_Stationary_matrix_5_5,
  input  [15:0] io_Stationary_matrix_5_6,
  input  [15:0] io_Stationary_matrix_5_7,
  input  [15:0] io_Stationary_matrix_6_0,
  input  [15:0] io_Stationary_matrix_6_1,
  input  [15:0] io_Stationary_matrix_6_2,
  input  [15:0] io_Stationary_matrix_6_3,
  input  [15:0] io_Stationary_matrix_6_4,
  input  [15:0] io_Stationary_matrix_6_5,
  input  [15:0] io_Stationary_matrix_6_6,
  input  [15:0] io_Stationary_matrix_6_7,
  input  [15:0] io_Stationary_matrix_7_0,
  input  [15:0] io_Stationary_matrix_7_1,
  input  [15:0] io_Stationary_matrix_7_2,
  input  [15:0] io_Stationary_matrix_7_3,
  input  [15:0] io_Stationary_matrix_7_4,
  input  [15:0] io_Stationary_matrix_7_5,
  input  [15:0] io_Stationary_matrix_7_6,
  input  [15:0] io_Stationary_matrix_7_7,
  output [4:0]  io_o_vn_0_0,
  output [4:0]  io_o_vn_0_1,
  output [4:0]  io_o_vn_0_2,
  output [4:0]  io_o_vn_0_3,
  output [4:0]  io_o_vn_1_0,
  output [4:0]  io_o_vn_1_1,
  output [4:0]  io_o_vn_1_2,
  output [4:0]  io_o_vn_1_3,
  output [4:0]  io_o_vn_2_0,
  output [4:0]  io_o_vn_2_1,
  output [4:0]  io_o_vn_2_2,
  output [4:0]  io_o_vn_2_3,
  output [4:0]  io_o_vn_3_0,
  output [4:0]  io_o_vn_3_1,
  output [4:0]  io_o_vn_3_2,
  output [4:0]  io_o_vn_3_3,
  output [4:0]  io_o_vn_4_0,
  output [4:0]  io_o_vn_4_1,
  output [4:0]  io_o_vn_4_2,
  output [4:0]  io_o_vn_4_3,
  output [4:0]  io_o_vn_5_0,
  output [4:0]  io_o_vn_5_1,
  output [4:0]  io_o_vn_5_2,
  output [4:0]  io_o_vn_5_3,
  output [4:0]  io_o_vn_6_0,
  output [4:0]  io_o_vn_6_1,
  output [4:0]  io_o_vn_6_2,
  output [4:0]  io_o_vn_6_3,
  output [4:0]  io_o_vn_7_0,
  output [4:0]  io_o_vn_7_1,
  output [4:0]  io_o_vn_7_2,
  output [4:0]  io_o_vn_7_3,
  output [4:0]  io_o_vn_8_0,
  output [4:0]  io_o_vn_8_1,
  output [4:0]  io_o_vn_8_2,
  output [4:0]  io_o_vn_8_3,
  output [4:0]  io_o_vn_9_0,
  output [4:0]  io_o_vn_9_1,
  output [4:0]  io_o_vn_9_2,
  output [4:0]  io_o_vn_9_3,
  output [4:0]  io_o_vn_10_0,
  output [4:0]  io_o_vn_10_1,
  output [4:0]  io_o_vn_10_2,
  output [4:0]  io_o_vn_10_3,
  output [4:0]  io_o_vn_11_0,
  output [4:0]  io_o_vn_11_1,
  output [4:0]  io_o_vn_11_2,
  output [4:0]  io_o_vn_11_3,
  output [4:0]  io_o_vn_12_0,
  output [4:0]  io_o_vn_12_1,
  output [4:0]  io_o_vn_12_2,
  output [4:0]  io_o_vn_12_3,
  output [4:0]  io_o_vn_13_0,
  output [4:0]  io_o_vn_13_1,
  output [4:0]  io_o_vn_13_2,
  output [4:0]  io_o_vn_13_3,
  output [4:0]  io_o_vn_14_0,
  output [4:0]  io_o_vn_14_1,
  output [4:0]  io_o_vn_14_2,
  output [4:0]  io_o_vn_14_3,
  output [4:0]  io_o_vn_15_0,
  output [4:0]  io_o_vn_15_1,
  output [4:0]  io_o_vn_15_2,
  output [4:0]  io_o_vn_15_3
);
  wire  my_stationary_clock; // @[ivntop.scala 19:31]
  wire  my_stationary_reset; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_0_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_0_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_0_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_0_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_0_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_0_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_0_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_0_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_1_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_1_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_1_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_1_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_1_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_1_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_1_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_1_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_2_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_2_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_2_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_2_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_2_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_2_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_2_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_2_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_3_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_3_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_3_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_3_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_3_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_3_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_3_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_3_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_4_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_4_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_4_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_4_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_4_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_4_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_4_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_4_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_5_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_5_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_5_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_5_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_5_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_5_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_5_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_5_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_6_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_6_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_6_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_6_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_6_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_6_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_6_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_6_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_7_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_7_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_7_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_7_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_7_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_7_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_7_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_Stationary_matrix_7_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_0_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_0_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_0_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_0_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_0_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_0_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_0_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_0_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_1_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_1_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_1_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_1_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_1_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_1_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_1_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_1_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_2_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_2_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_2_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_2_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_2_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_2_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_2_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_2_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_3_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_3_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_3_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_3_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_3_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_3_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_3_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_3_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_4_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_4_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_4_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_4_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_4_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_4_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_4_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_4_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_5_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_5_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_5_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_5_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_5_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_5_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_5_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_5_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_6_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_6_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_6_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_6_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_6_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_6_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_6_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_6_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_7_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_7_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_7_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_7_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_7_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_7_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_7_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_7_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_0_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_0_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_0_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_0_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_0_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_0_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_0_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_0_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_1_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_1_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_1_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_1_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_1_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_1_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_1_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_1_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_2_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_2_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_2_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_2_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_2_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_2_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_2_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_2_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_3_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_3_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_3_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_3_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_3_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_3_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_3_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_3_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_4_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_4_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_4_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_4_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_4_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_4_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_4_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_4_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_5_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_5_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_5_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_5_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_5_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_5_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_5_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_5_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_6_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_6_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_6_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_6_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_6_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_6_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_6_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_6_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_7_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_7_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_7_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_7_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_7_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_7_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_7_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_7_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_0_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_0_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_0_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_0_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_0_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_0_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_0_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_0_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_1_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_1_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_1_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_1_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_1_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_1_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_1_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_1_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_2_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_2_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_2_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_2_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_2_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_2_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_2_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_2_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_3_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_3_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_3_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_3_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_3_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_3_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_3_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_3_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_4_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_4_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_4_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_4_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_4_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_4_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_4_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_4_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_5_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_5_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_5_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_5_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_5_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_5_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_5_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_5_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_6_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_6_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_6_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_6_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_6_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_6_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_6_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_6_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_7_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_7_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_7_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_7_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_7_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_7_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_7_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_7_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_0_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_0_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_0_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_0_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_0_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_0_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_0_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_0_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_1_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_1_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_1_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_1_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_1_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_1_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_1_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_1_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_2_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_2_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_2_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_2_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_2_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_2_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_2_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_2_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_3_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_3_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_3_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_3_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_3_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_3_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_3_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_3_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_4_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_4_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_4_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_4_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_4_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_4_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_4_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_4_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_5_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_5_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_5_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_5_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_5_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_5_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_5_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_5_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_6_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_6_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_6_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_6_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_6_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_6_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_6_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_6_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_7_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_7_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_7_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_7_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_7_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_7_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_7_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_7_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_0_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_0_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_0_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_0_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_0_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_0_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_0_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_0_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_1_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_1_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_1_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_1_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_1_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_1_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_1_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_1_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_2_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_2_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_2_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_2_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_2_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_2_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_2_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_2_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_3_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_3_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_3_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_3_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_3_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_3_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_3_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_3_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_4_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_4_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_4_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_4_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_4_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_4_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_4_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_4_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_5_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_5_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_5_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_5_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_5_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_5_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_5_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_5_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_6_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_6_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_6_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_6_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_6_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_6_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_6_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_6_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_7_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_7_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_7_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_7_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_7_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_7_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_7_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_7_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_0_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_0_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_0_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_0_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_0_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_0_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_0_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_0_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_1_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_1_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_1_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_1_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_1_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_1_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_1_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_1_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_2_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_2_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_2_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_2_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_2_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_2_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_2_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_2_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_3_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_3_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_3_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_3_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_3_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_3_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_3_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_3_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_4_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_4_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_4_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_4_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_4_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_4_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_4_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_4_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_5_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_5_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_5_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_5_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_5_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_5_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_5_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_5_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_6_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_6_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_6_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_6_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_6_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_6_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_6_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_6_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_7_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_7_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_7_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_7_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_7_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_7_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_7_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_7_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_0_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_0_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_0_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_0_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_0_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_0_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_0_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_0_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_1_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_1_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_1_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_1_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_1_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_1_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_1_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_1_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_2_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_2_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_2_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_2_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_2_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_2_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_2_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_2_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_3_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_3_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_3_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_3_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_3_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_3_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_3_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_3_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_4_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_4_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_4_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_4_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_4_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_4_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_4_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_4_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_5_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_5_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_5_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_5_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_5_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_5_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_5_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_5_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_6_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_6_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_6_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_6_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_6_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_6_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_6_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_6_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_7_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_7_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_7_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_7_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_7_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_7_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_7_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_7_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_0_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_0_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_0_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_0_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_0_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_0_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_0_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_0_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_1_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_1_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_1_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_1_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_1_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_1_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_1_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_1_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_2_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_2_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_2_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_2_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_2_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_2_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_2_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_2_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_3_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_3_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_3_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_3_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_3_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_3_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_3_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_3_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_4_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_4_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_4_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_4_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_4_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_4_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_4_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_4_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_5_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_5_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_5_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_5_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_5_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_5_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_5_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_5_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_6_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_6_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_6_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_6_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_6_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_6_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_6_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_6_7; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_7_0; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_7_1; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_7_2; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_7_3; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_7_4; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_7_5; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_7_6; // @[ivntop.scala 19:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_7_7; // @[ivntop.scala 19:31]
  wire  my_ivn1_clock; // @[ivntop.scala 32:24]
  wire  my_ivn1_reset; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_0_0; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_0_1; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_0_2; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_0_3; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_0_4; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_0_5; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_0_6; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_0_7; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_1_0; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_1_1; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_1_2; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_1_3; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_1_4; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_1_5; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_1_6; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_1_7; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_2_0; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_2_1; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_2_2; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_2_3; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_2_4; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_2_5; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_2_6; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_2_7; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_3_0; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_3_1; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_3_2; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_3_3; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_3_4; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_3_5; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_3_6; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_3_7; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_4_0; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_4_1; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_4_2; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_4_3; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_4_4; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_4_5; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_4_6; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_4_7; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_5_0; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_5_1; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_5_2; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_5_3; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_5_4; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_5_5; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_5_6; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_5_7; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_6_0; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_6_1; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_6_2; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_6_3; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_6_4; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_6_5; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_6_6; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_6_7; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_7_0; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_7_1; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_7_2; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_7_3; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_7_4; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_7_5; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_7_6; // @[ivntop.scala 32:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_7_7; // @[ivntop.scala 32:24]
  wire [4:0] my_ivn1_io_o_vn_0; // @[ivntop.scala 32:24]
  wire [4:0] my_ivn1_io_o_vn_1; // @[ivntop.scala 32:24]
  wire [4:0] my_ivn1_io_o_vn_2; // @[ivntop.scala 32:24]
  wire [4:0] my_ivn1_io_o_vn_3; // @[ivntop.scala 32:24]
  wire [4:0] my_ivn1_io_o_vn2_0; // @[ivntop.scala 32:24]
  wire [4:0] my_ivn1_io_o_vn2_1; // @[ivntop.scala 32:24]
  wire [4:0] my_ivn1_io_o_vn2_2; // @[ivntop.scala 32:24]
  wire [4:0] my_ivn1_io_o_vn2_3; // @[ivntop.scala 32:24]
  wire  my_ivn1_io_ProcessValid; // @[ivntop.scala 32:24]
  wire  my_ivn2_clock; // @[ivntop.scala 40:24]
  wire  my_ivn2_reset; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_0_0; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_0_1; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_0_2; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_0_3; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_0_4; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_0_5; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_0_6; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_0_7; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_1_0; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_1_1; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_1_2; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_1_3; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_1_4; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_1_5; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_1_6; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_1_7; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_2_0; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_2_1; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_2_2; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_2_3; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_2_4; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_2_5; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_2_6; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_2_7; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_3_0; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_3_1; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_3_2; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_3_3; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_3_4; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_3_5; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_3_6; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_3_7; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_4_0; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_4_1; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_4_2; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_4_3; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_4_4; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_4_5; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_4_6; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_4_7; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_5_0; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_5_1; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_5_2; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_5_3; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_5_4; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_5_5; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_5_6; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_5_7; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_6_0; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_6_1; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_6_2; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_6_3; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_6_4; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_6_5; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_6_6; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_6_7; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_7_0; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_7_1; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_7_2; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_7_3; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_7_4; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_7_5; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_7_6; // @[ivntop.scala 40:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_7_7; // @[ivntop.scala 40:24]
  wire [4:0] my_ivn2_io_o_vn_0; // @[ivntop.scala 40:24]
  wire [4:0] my_ivn2_io_o_vn_1; // @[ivntop.scala 40:24]
  wire [4:0] my_ivn2_io_o_vn_2; // @[ivntop.scala 40:24]
  wire [4:0] my_ivn2_io_o_vn_3; // @[ivntop.scala 40:24]
  wire [4:0] my_ivn2_io_o_vn2_0; // @[ivntop.scala 40:24]
  wire [4:0] my_ivn2_io_o_vn2_1; // @[ivntop.scala 40:24]
  wire [4:0] my_ivn2_io_o_vn2_2; // @[ivntop.scala 40:24]
  wire [4:0] my_ivn2_io_o_vn2_3; // @[ivntop.scala 40:24]
  wire  my_ivn3_clock; // @[ivntop.scala 47:25]
  wire  my_ivn3_reset; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_0_0; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_0_1; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_0_2; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_0_3; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_0_4; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_0_5; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_0_6; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_0_7; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_1_0; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_1_1; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_1_2; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_1_3; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_1_4; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_1_5; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_1_6; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_1_7; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_2_0; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_2_1; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_2_2; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_2_3; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_2_4; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_2_5; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_2_6; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_2_7; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_3_0; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_3_1; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_3_2; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_3_3; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_3_4; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_3_5; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_3_6; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_3_7; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_4_0; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_4_1; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_4_2; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_4_3; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_4_4; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_4_5; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_4_6; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_4_7; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_5_0; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_5_1; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_5_2; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_5_3; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_5_4; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_5_5; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_5_6; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_5_7; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_6_0; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_6_1; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_6_2; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_6_3; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_6_4; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_6_5; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_6_6; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_6_7; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_7_0; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_7_1; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_7_2; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_7_3; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_7_4; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_7_5; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_7_6; // @[ivntop.scala 47:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_7_7; // @[ivntop.scala 47:25]
  wire [4:0] my_ivn3_io_o_vn_0; // @[ivntop.scala 47:25]
  wire [4:0] my_ivn3_io_o_vn_1; // @[ivntop.scala 47:25]
  wire [4:0] my_ivn3_io_o_vn_2; // @[ivntop.scala 47:25]
  wire [4:0] my_ivn3_io_o_vn_3; // @[ivntop.scala 47:25]
  wire [4:0] my_ivn3_io_o_vn2_0; // @[ivntop.scala 47:25]
  wire [4:0] my_ivn3_io_o_vn2_1; // @[ivntop.scala 47:25]
  wire [4:0] my_ivn3_io_o_vn2_2; // @[ivntop.scala 47:25]
  wire [4:0] my_ivn3_io_o_vn2_3; // @[ivntop.scala 47:25]
  wire  my_ivn4_clock; // @[ivntop.scala 54:25]
  wire  my_ivn4_reset; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_0_0; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_0_1; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_0_2; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_0_3; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_0_4; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_0_5; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_0_6; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_0_7; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_1_0; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_1_1; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_1_2; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_1_3; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_1_4; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_1_5; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_1_6; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_1_7; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_2_0; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_2_1; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_2_2; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_2_3; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_2_4; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_2_5; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_2_6; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_2_7; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_3_0; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_3_1; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_3_2; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_3_3; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_3_4; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_3_5; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_3_6; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_3_7; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_4_0; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_4_1; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_4_2; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_4_3; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_4_4; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_4_5; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_4_6; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_4_7; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_5_0; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_5_1; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_5_2; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_5_3; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_5_4; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_5_5; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_5_6; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_5_7; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_6_0; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_6_1; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_6_2; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_6_3; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_6_4; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_6_5; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_6_6; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_6_7; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_7_0; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_7_1; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_7_2; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_7_3; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_7_4; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_7_5; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_7_6; // @[ivntop.scala 54:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_7_7; // @[ivntop.scala 54:25]
  wire [4:0] my_ivn4_io_o_vn_0; // @[ivntop.scala 54:25]
  wire [4:0] my_ivn4_io_o_vn_1; // @[ivntop.scala 54:25]
  wire [4:0] my_ivn4_io_o_vn_2; // @[ivntop.scala 54:25]
  wire [4:0] my_ivn4_io_o_vn_3; // @[ivntop.scala 54:25]
  wire [4:0] my_ivn4_io_o_vn2_0; // @[ivntop.scala 54:25]
  wire [4:0] my_ivn4_io_o_vn2_1; // @[ivntop.scala 54:25]
  wire [4:0] my_ivn4_io_o_vn2_2; // @[ivntop.scala 54:25]
  wire [4:0] my_ivn4_io_o_vn2_3; // @[ivntop.scala 54:25]
  wire  my_ivn5_clock; // @[ivntop.scala 61:25]
  wire  my_ivn5_reset; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_0_0; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_0_1; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_0_2; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_0_3; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_0_4; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_0_5; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_0_6; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_0_7; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_1_0; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_1_1; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_1_2; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_1_3; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_1_4; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_1_5; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_1_6; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_1_7; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_2_0; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_2_1; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_2_2; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_2_3; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_2_4; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_2_5; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_2_6; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_2_7; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_3_0; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_3_1; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_3_2; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_3_3; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_3_4; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_3_5; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_3_6; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_3_7; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_4_0; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_4_1; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_4_2; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_4_3; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_4_4; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_4_5; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_4_6; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_4_7; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_5_0; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_5_1; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_5_2; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_5_3; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_5_4; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_5_5; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_5_6; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_5_7; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_6_0; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_6_1; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_6_2; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_6_3; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_6_4; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_6_5; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_6_6; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_6_7; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_7_0; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_7_1; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_7_2; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_7_3; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_7_4; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_7_5; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_7_6; // @[ivntop.scala 61:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_7_7; // @[ivntop.scala 61:25]
  wire [4:0] my_ivn5_io_o_vn_0; // @[ivntop.scala 61:25]
  wire [4:0] my_ivn5_io_o_vn_1; // @[ivntop.scala 61:25]
  wire [4:0] my_ivn5_io_o_vn_2; // @[ivntop.scala 61:25]
  wire [4:0] my_ivn5_io_o_vn_3; // @[ivntop.scala 61:25]
  wire [4:0] my_ivn5_io_o_vn2_0; // @[ivntop.scala 61:25]
  wire [4:0] my_ivn5_io_o_vn2_1; // @[ivntop.scala 61:25]
  wire [4:0] my_ivn5_io_o_vn2_2; // @[ivntop.scala 61:25]
  wire [4:0] my_ivn5_io_o_vn2_3; // @[ivntop.scala 61:25]
  wire  my_ivn6_clock; // @[ivntop.scala 68:25]
  wire  my_ivn6_reset; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_0_0; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_0_1; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_0_2; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_0_3; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_0_4; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_0_5; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_0_6; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_0_7; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_1_0; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_1_1; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_1_2; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_1_3; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_1_4; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_1_5; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_1_6; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_1_7; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_2_0; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_2_1; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_2_2; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_2_3; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_2_4; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_2_5; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_2_6; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_2_7; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_3_0; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_3_1; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_3_2; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_3_3; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_3_4; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_3_5; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_3_6; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_3_7; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_4_0; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_4_1; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_4_2; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_4_3; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_4_4; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_4_5; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_4_6; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_4_7; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_5_0; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_5_1; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_5_2; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_5_3; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_5_4; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_5_5; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_5_6; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_5_7; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_6_0; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_6_1; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_6_2; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_6_3; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_6_4; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_6_5; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_6_6; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_6_7; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_7_0; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_7_1; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_7_2; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_7_3; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_7_4; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_7_5; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_7_6; // @[ivntop.scala 68:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_7_7; // @[ivntop.scala 68:25]
  wire [4:0] my_ivn6_io_o_vn_0; // @[ivntop.scala 68:25]
  wire [4:0] my_ivn6_io_o_vn_1; // @[ivntop.scala 68:25]
  wire [4:0] my_ivn6_io_o_vn_2; // @[ivntop.scala 68:25]
  wire [4:0] my_ivn6_io_o_vn_3; // @[ivntop.scala 68:25]
  wire [4:0] my_ivn6_io_o_vn2_0; // @[ivntop.scala 68:25]
  wire [4:0] my_ivn6_io_o_vn2_1; // @[ivntop.scala 68:25]
  wire [4:0] my_ivn6_io_o_vn2_2; // @[ivntop.scala 68:25]
  wire [4:0] my_ivn6_io_o_vn2_3; // @[ivntop.scala 68:25]
  wire  my_ivn7_clock; // @[ivntop.scala 75:25]
  wire  my_ivn7_reset; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_0_0; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_0_1; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_0_2; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_0_3; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_0_4; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_0_5; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_0_6; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_0_7; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_1_0; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_1_1; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_1_2; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_1_3; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_1_4; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_1_5; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_1_6; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_1_7; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_2_0; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_2_1; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_2_2; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_2_3; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_2_4; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_2_5; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_2_6; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_2_7; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_3_0; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_3_1; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_3_2; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_3_3; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_3_4; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_3_5; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_3_6; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_3_7; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_4_0; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_4_1; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_4_2; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_4_3; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_4_4; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_4_5; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_4_6; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_4_7; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_5_0; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_5_1; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_5_2; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_5_3; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_5_4; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_5_5; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_5_6; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_5_7; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_6_0; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_6_1; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_6_2; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_6_3; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_6_4; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_6_5; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_6_6; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_6_7; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_7_0; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_7_1; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_7_2; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_7_3; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_7_4; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_7_5; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_7_6; // @[ivntop.scala 75:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_7_7; // @[ivntop.scala 75:25]
  wire [4:0] my_ivn7_io_o_vn_0; // @[ivntop.scala 75:25]
  wire [4:0] my_ivn7_io_o_vn_1; // @[ivntop.scala 75:25]
  wire [4:0] my_ivn7_io_o_vn_2; // @[ivntop.scala 75:25]
  wire [4:0] my_ivn7_io_o_vn_3; // @[ivntop.scala 75:25]
  wire [4:0] my_ivn7_io_o_vn2_0; // @[ivntop.scala 75:25]
  wire [4:0] my_ivn7_io_o_vn2_1; // @[ivntop.scala 75:25]
  wire [4:0] my_ivn7_io_o_vn2_2; // @[ivntop.scala 75:25]
  wire [4:0] my_ivn7_io_o_vn2_3; // @[ivntop.scala 75:25]
  wire  my_ivn8_clock; // @[ivntop.scala 82:25]
  wire  my_ivn8_reset; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_0_0; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_0_1; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_0_2; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_0_3; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_0_4; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_0_5; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_0_6; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_0_7; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_1_0; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_1_1; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_1_2; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_1_3; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_1_4; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_1_5; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_1_6; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_1_7; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_2_0; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_2_1; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_2_2; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_2_3; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_2_4; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_2_5; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_2_6; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_2_7; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_3_0; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_3_1; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_3_2; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_3_3; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_3_4; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_3_5; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_3_6; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_3_7; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_4_0; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_4_1; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_4_2; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_4_3; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_4_4; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_4_5; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_4_6; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_4_7; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_5_0; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_5_1; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_5_2; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_5_3; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_5_4; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_5_5; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_5_6; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_5_7; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_6_0; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_6_1; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_6_2; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_6_3; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_6_4; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_6_5; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_6_6; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_6_7; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_7_0; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_7_1; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_7_2; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_7_3; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_7_4; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_7_5; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_7_6; // @[ivntop.scala 82:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_7_7; // @[ivntop.scala 82:25]
  wire [4:0] my_ivn8_io_o_vn_0; // @[ivntop.scala 82:25]
  wire [4:0] my_ivn8_io_o_vn_1; // @[ivntop.scala 82:25]
  wire [4:0] my_ivn8_io_o_vn_2; // @[ivntop.scala 82:25]
  wire [4:0] my_ivn8_io_o_vn_3; // @[ivntop.scala 82:25]
  wire [4:0] my_ivn8_io_o_vn2_0; // @[ivntop.scala 82:25]
  wire [4:0] my_ivn8_io_o_vn2_1; // @[ivntop.scala 82:25]
  wire [4:0] my_ivn8_io_o_vn2_2; // @[ivntop.scala 82:25]
  wire [4:0] my_ivn8_io_o_vn2_3; // @[ivntop.scala 82:25]
  stationary my_stationary ( // @[ivntop.scala 19:31]
    .clock(my_stationary_clock),
    .reset(my_stationary_reset),
    .io_Stationary_matrix_0_0(my_stationary_io_Stationary_matrix_0_0),
    .io_Stationary_matrix_0_1(my_stationary_io_Stationary_matrix_0_1),
    .io_Stationary_matrix_0_2(my_stationary_io_Stationary_matrix_0_2),
    .io_Stationary_matrix_0_3(my_stationary_io_Stationary_matrix_0_3),
    .io_Stationary_matrix_0_4(my_stationary_io_Stationary_matrix_0_4),
    .io_Stationary_matrix_0_5(my_stationary_io_Stationary_matrix_0_5),
    .io_Stationary_matrix_0_6(my_stationary_io_Stationary_matrix_0_6),
    .io_Stationary_matrix_0_7(my_stationary_io_Stationary_matrix_0_7),
    .io_Stationary_matrix_1_0(my_stationary_io_Stationary_matrix_1_0),
    .io_Stationary_matrix_1_1(my_stationary_io_Stationary_matrix_1_1),
    .io_Stationary_matrix_1_2(my_stationary_io_Stationary_matrix_1_2),
    .io_Stationary_matrix_1_3(my_stationary_io_Stationary_matrix_1_3),
    .io_Stationary_matrix_1_4(my_stationary_io_Stationary_matrix_1_4),
    .io_Stationary_matrix_1_5(my_stationary_io_Stationary_matrix_1_5),
    .io_Stationary_matrix_1_6(my_stationary_io_Stationary_matrix_1_6),
    .io_Stationary_matrix_1_7(my_stationary_io_Stationary_matrix_1_7),
    .io_Stationary_matrix_2_0(my_stationary_io_Stationary_matrix_2_0),
    .io_Stationary_matrix_2_1(my_stationary_io_Stationary_matrix_2_1),
    .io_Stationary_matrix_2_2(my_stationary_io_Stationary_matrix_2_2),
    .io_Stationary_matrix_2_3(my_stationary_io_Stationary_matrix_2_3),
    .io_Stationary_matrix_2_4(my_stationary_io_Stationary_matrix_2_4),
    .io_Stationary_matrix_2_5(my_stationary_io_Stationary_matrix_2_5),
    .io_Stationary_matrix_2_6(my_stationary_io_Stationary_matrix_2_6),
    .io_Stationary_matrix_2_7(my_stationary_io_Stationary_matrix_2_7),
    .io_Stationary_matrix_3_0(my_stationary_io_Stationary_matrix_3_0),
    .io_Stationary_matrix_3_1(my_stationary_io_Stationary_matrix_3_1),
    .io_Stationary_matrix_3_2(my_stationary_io_Stationary_matrix_3_2),
    .io_Stationary_matrix_3_3(my_stationary_io_Stationary_matrix_3_3),
    .io_Stationary_matrix_3_4(my_stationary_io_Stationary_matrix_3_4),
    .io_Stationary_matrix_3_5(my_stationary_io_Stationary_matrix_3_5),
    .io_Stationary_matrix_3_6(my_stationary_io_Stationary_matrix_3_6),
    .io_Stationary_matrix_3_7(my_stationary_io_Stationary_matrix_3_7),
    .io_Stationary_matrix_4_0(my_stationary_io_Stationary_matrix_4_0),
    .io_Stationary_matrix_4_1(my_stationary_io_Stationary_matrix_4_1),
    .io_Stationary_matrix_4_2(my_stationary_io_Stationary_matrix_4_2),
    .io_Stationary_matrix_4_3(my_stationary_io_Stationary_matrix_4_3),
    .io_Stationary_matrix_4_4(my_stationary_io_Stationary_matrix_4_4),
    .io_Stationary_matrix_4_5(my_stationary_io_Stationary_matrix_4_5),
    .io_Stationary_matrix_4_6(my_stationary_io_Stationary_matrix_4_6),
    .io_Stationary_matrix_4_7(my_stationary_io_Stationary_matrix_4_7),
    .io_Stationary_matrix_5_0(my_stationary_io_Stationary_matrix_5_0),
    .io_Stationary_matrix_5_1(my_stationary_io_Stationary_matrix_5_1),
    .io_Stationary_matrix_5_2(my_stationary_io_Stationary_matrix_5_2),
    .io_Stationary_matrix_5_3(my_stationary_io_Stationary_matrix_5_3),
    .io_Stationary_matrix_5_4(my_stationary_io_Stationary_matrix_5_4),
    .io_Stationary_matrix_5_5(my_stationary_io_Stationary_matrix_5_5),
    .io_Stationary_matrix_5_6(my_stationary_io_Stationary_matrix_5_6),
    .io_Stationary_matrix_5_7(my_stationary_io_Stationary_matrix_5_7),
    .io_Stationary_matrix_6_0(my_stationary_io_Stationary_matrix_6_0),
    .io_Stationary_matrix_6_1(my_stationary_io_Stationary_matrix_6_1),
    .io_Stationary_matrix_6_2(my_stationary_io_Stationary_matrix_6_2),
    .io_Stationary_matrix_6_3(my_stationary_io_Stationary_matrix_6_3),
    .io_Stationary_matrix_6_4(my_stationary_io_Stationary_matrix_6_4),
    .io_Stationary_matrix_6_5(my_stationary_io_Stationary_matrix_6_5),
    .io_Stationary_matrix_6_6(my_stationary_io_Stationary_matrix_6_6),
    .io_Stationary_matrix_6_7(my_stationary_io_Stationary_matrix_6_7),
    .io_Stationary_matrix_7_0(my_stationary_io_Stationary_matrix_7_0),
    .io_Stationary_matrix_7_1(my_stationary_io_Stationary_matrix_7_1),
    .io_Stationary_matrix_7_2(my_stationary_io_Stationary_matrix_7_2),
    .io_Stationary_matrix_7_3(my_stationary_io_Stationary_matrix_7_3),
    .io_Stationary_matrix_7_4(my_stationary_io_Stationary_matrix_7_4),
    .io_Stationary_matrix_7_5(my_stationary_io_Stationary_matrix_7_5),
    .io_Stationary_matrix_7_6(my_stationary_io_Stationary_matrix_7_6),
    .io_Stationary_matrix_7_7(my_stationary_io_Stationary_matrix_7_7),
    .io_o_Stationary_matrix1_0_0(my_stationary_io_o_Stationary_matrix1_0_0),
    .io_o_Stationary_matrix1_0_1(my_stationary_io_o_Stationary_matrix1_0_1),
    .io_o_Stationary_matrix1_0_2(my_stationary_io_o_Stationary_matrix1_0_2),
    .io_o_Stationary_matrix1_0_3(my_stationary_io_o_Stationary_matrix1_0_3),
    .io_o_Stationary_matrix1_0_4(my_stationary_io_o_Stationary_matrix1_0_4),
    .io_o_Stationary_matrix1_0_5(my_stationary_io_o_Stationary_matrix1_0_5),
    .io_o_Stationary_matrix1_0_6(my_stationary_io_o_Stationary_matrix1_0_6),
    .io_o_Stationary_matrix1_0_7(my_stationary_io_o_Stationary_matrix1_0_7),
    .io_o_Stationary_matrix1_1_0(my_stationary_io_o_Stationary_matrix1_1_0),
    .io_o_Stationary_matrix1_1_1(my_stationary_io_o_Stationary_matrix1_1_1),
    .io_o_Stationary_matrix1_1_2(my_stationary_io_o_Stationary_matrix1_1_2),
    .io_o_Stationary_matrix1_1_3(my_stationary_io_o_Stationary_matrix1_1_3),
    .io_o_Stationary_matrix1_1_4(my_stationary_io_o_Stationary_matrix1_1_4),
    .io_o_Stationary_matrix1_1_5(my_stationary_io_o_Stationary_matrix1_1_5),
    .io_o_Stationary_matrix1_1_6(my_stationary_io_o_Stationary_matrix1_1_6),
    .io_o_Stationary_matrix1_1_7(my_stationary_io_o_Stationary_matrix1_1_7),
    .io_o_Stationary_matrix1_2_0(my_stationary_io_o_Stationary_matrix1_2_0),
    .io_o_Stationary_matrix1_2_1(my_stationary_io_o_Stationary_matrix1_2_1),
    .io_o_Stationary_matrix1_2_2(my_stationary_io_o_Stationary_matrix1_2_2),
    .io_o_Stationary_matrix1_2_3(my_stationary_io_o_Stationary_matrix1_2_3),
    .io_o_Stationary_matrix1_2_4(my_stationary_io_o_Stationary_matrix1_2_4),
    .io_o_Stationary_matrix1_2_5(my_stationary_io_o_Stationary_matrix1_2_5),
    .io_o_Stationary_matrix1_2_6(my_stationary_io_o_Stationary_matrix1_2_6),
    .io_o_Stationary_matrix1_2_7(my_stationary_io_o_Stationary_matrix1_2_7),
    .io_o_Stationary_matrix1_3_0(my_stationary_io_o_Stationary_matrix1_3_0),
    .io_o_Stationary_matrix1_3_1(my_stationary_io_o_Stationary_matrix1_3_1),
    .io_o_Stationary_matrix1_3_2(my_stationary_io_o_Stationary_matrix1_3_2),
    .io_o_Stationary_matrix1_3_3(my_stationary_io_o_Stationary_matrix1_3_3),
    .io_o_Stationary_matrix1_3_4(my_stationary_io_o_Stationary_matrix1_3_4),
    .io_o_Stationary_matrix1_3_5(my_stationary_io_o_Stationary_matrix1_3_5),
    .io_o_Stationary_matrix1_3_6(my_stationary_io_o_Stationary_matrix1_3_6),
    .io_o_Stationary_matrix1_3_7(my_stationary_io_o_Stationary_matrix1_3_7),
    .io_o_Stationary_matrix1_4_0(my_stationary_io_o_Stationary_matrix1_4_0),
    .io_o_Stationary_matrix1_4_1(my_stationary_io_o_Stationary_matrix1_4_1),
    .io_o_Stationary_matrix1_4_2(my_stationary_io_o_Stationary_matrix1_4_2),
    .io_o_Stationary_matrix1_4_3(my_stationary_io_o_Stationary_matrix1_4_3),
    .io_o_Stationary_matrix1_4_4(my_stationary_io_o_Stationary_matrix1_4_4),
    .io_o_Stationary_matrix1_4_5(my_stationary_io_o_Stationary_matrix1_4_5),
    .io_o_Stationary_matrix1_4_6(my_stationary_io_o_Stationary_matrix1_4_6),
    .io_o_Stationary_matrix1_4_7(my_stationary_io_o_Stationary_matrix1_4_7),
    .io_o_Stationary_matrix1_5_0(my_stationary_io_o_Stationary_matrix1_5_0),
    .io_o_Stationary_matrix1_5_1(my_stationary_io_o_Stationary_matrix1_5_1),
    .io_o_Stationary_matrix1_5_2(my_stationary_io_o_Stationary_matrix1_5_2),
    .io_o_Stationary_matrix1_5_3(my_stationary_io_o_Stationary_matrix1_5_3),
    .io_o_Stationary_matrix1_5_4(my_stationary_io_o_Stationary_matrix1_5_4),
    .io_o_Stationary_matrix1_5_5(my_stationary_io_o_Stationary_matrix1_5_5),
    .io_o_Stationary_matrix1_5_6(my_stationary_io_o_Stationary_matrix1_5_6),
    .io_o_Stationary_matrix1_5_7(my_stationary_io_o_Stationary_matrix1_5_7),
    .io_o_Stationary_matrix1_6_0(my_stationary_io_o_Stationary_matrix1_6_0),
    .io_o_Stationary_matrix1_6_1(my_stationary_io_o_Stationary_matrix1_6_1),
    .io_o_Stationary_matrix1_6_2(my_stationary_io_o_Stationary_matrix1_6_2),
    .io_o_Stationary_matrix1_6_3(my_stationary_io_o_Stationary_matrix1_6_3),
    .io_o_Stationary_matrix1_6_4(my_stationary_io_o_Stationary_matrix1_6_4),
    .io_o_Stationary_matrix1_6_5(my_stationary_io_o_Stationary_matrix1_6_5),
    .io_o_Stationary_matrix1_6_6(my_stationary_io_o_Stationary_matrix1_6_6),
    .io_o_Stationary_matrix1_6_7(my_stationary_io_o_Stationary_matrix1_6_7),
    .io_o_Stationary_matrix1_7_0(my_stationary_io_o_Stationary_matrix1_7_0),
    .io_o_Stationary_matrix1_7_1(my_stationary_io_o_Stationary_matrix1_7_1),
    .io_o_Stationary_matrix1_7_2(my_stationary_io_o_Stationary_matrix1_7_2),
    .io_o_Stationary_matrix1_7_3(my_stationary_io_o_Stationary_matrix1_7_3),
    .io_o_Stationary_matrix1_7_4(my_stationary_io_o_Stationary_matrix1_7_4),
    .io_o_Stationary_matrix1_7_5(my_stationary_io_o_Stationary_matrix1_7_5),
    .io_o_Stationary_matrix1_7_6(my_stationary_io_o_Stationary_matrix1_7_6),
    .io_o_Stationary_matrix1_7_7(my_stationary_io_o_Stationary_matrix1_7_7),
    .io_o_Stationary_matrix2_0_0(my_stationary_io_o_Stationary_matrix2_0_0),
    .io_o_Stationary_matrix2_0_1(my_stationary_io_o_Stationary_matrix2_0_1),
    .io_o_Stationary_matrix2_0_2(my_stationary_io_o_Stationary_matrix2_0_2),
    .io_o_Stationary_matrix2_0_3(my_stationary_io_o_Stationary_matrix2_0_3),
    .io_o_Stationary_matrix2_0_4(my_stationary_io_o_Stationary_matrix2_0_4),
    .io_o_Stationary_matrix2_0_5(my_stationary_io_o_Stationary_matrix2_0_5),
    .io_o_Stationary_matrix2_0_6(my_stationary_io_o_Stationary_matrix2_0_6),
    .io_o_Stationary_matrix2_0_7(my_stationary_io_o_Stationary_matrix2_0_7),
    .io_o_Stationary_matrix2_1_0(my_stationary_io_o_Stationary_matrix2_1_0),
    .io_o_Stationary_matrix2_1_1(my_stationary_io_o_Stationary_matrix2_1_1),
    .io_o_Stationary_matrix2_1_2(my_stationary_io_o_Stationary_matrix2_1_2),
    .io_o_Stationary_matrix2_1_3(my_stationary_io_o_Stationary_matrix2_1_3),
    .io_o_Stationary_matrix2_1_4(my_stationary_io_o_Stationary_matrix2_1_4),
    .io_o_Stationary_matrix2_1_5(my_stationary_io_o_Stationary_matrix2_1_5),
    .io_o_Stationary_matrix2_1_6(my_stationary_io_o_Stationary_matrix2_1_6),
    .io_o_Stationary_matrix2_1_7(my_stationary_io_o_Stationary_matrix2_1_7),
    .io_o_Stationary_matrix2_2_0(my_stationary_io_o_Stationary_matrix2_2_0),
    .io_o_Stationary_matrix2_2_1(my_stationary_io_o_Stationary_matrix2_2_1),
    .io_o_Stationary_matrix2_2_2(my_stationary_io_o_Stationary_matrix2_2_2),
    .io_o_Stationary_matrix2_2_3(my_stationary_io_o_Stationary_matrix2_2_3),
    .io_o_Stationary_matrix2_2_4(my_stationary_io_o_Stationary_matrix2_2_4),
    .io_o_Stationary_matrix2_2_5(my_stationary_io_o_Stationary_matrix2_2_5),
    .io_o_Stationary_matrix2_2_6(my_stationary_io_o_Stationary_matrix2_2_6),
    .io_o_Stationary_matrix2_2_7(my_stationary_io_o_Stationary_matrix2_2_7),
    .io_o_Stationary_matrix2_3_0(my_stationary_io_o_Stationary_matrix2_3_0),
    .io_o_Stationary_matrix2_3_1(my_stationary_io_o_Stationary_matrix2_3_1),
    .io_o_Stationary_matrix2_3_2(my_stationary_io_o_Stationary_matrix2_3_2),
    .io_o_Stationary_matrix2_3_3(my_stationary_io_o_Stationary_matrix2_3_3),
    .io_o_Stationary_matrix2_3_4(my_stationary_io_o_Stationary_matrix2_3_4),
    .io_o_Stationary_matrix2_3_5(my_stationary_io_o_Stationary_matrix2_3_5),
    .io_o_Stationary_matrix2_3_6(my_stationary_io_o_Stationary_matrix2_3_6),
    .io_o_Stationary_matrix2_3_7(my_stationary_io_o_Stationary_matrix2_3_7),
    .io_o_Stationary_matrix2_4_0(my_stationary_io_o_Stationary_matrix2_4_0),
    .io_o_Stationary_matrix2_4_1(my_stationary_io_o_Stationary_matrix2_4_1),
    .io_o_Stationary_matrix2_4_2(my_stationary_io_o_Stationary_matrix2_4_2),
    .io_o_Stationary_matrix2_4_3(my_stationary_io_o_Stationary_matrix2_4_3),
    .io_o_Stationary_matrix2_4_4(my_stationary_io_o_Stationary_matrix2_4_4),
    .io_o_Stationary_matrix2_4_5(my_stationary_io_o_Stationary_matrix2_4_5),
    .io_o_Stationary_matrix2_4_6(my_stationary_io_o_Stationary_matrix2_4_6),
    .io_o_Stationary_matrix2_4_7(my_stationary_io_o_Stationary_matrix2_4_7),
    .io_o_Stationary_matrix2_5_0(my_stationary_io_o_Stationary_matrix2_5_0),
    .io_o_Stationary_matrix2_5_1(my_stationary_io_o_Stationary_matrix2_5_1),
    .io_o_Stationary_matrix2_5_2(my_stationary_io_o_Stationary_matrix2_5_2),
    .io_o_Stationary_matrix2_5_3(my_stationary_io_o_Stationary_matrix2_5_3),
    .io_o_Stationary_matrix2_5_4(my_stationary_io_o_Stationary_matrix2_5_4),
    .io_o_Stationary_matrix2_5_5(my_stationary_io_o_Stationary_matrix2_5_5),
    .io_o_Stationary_matrix2_5_6(my_stationary_io_o_Stationary_matrix2_5_6),
    .io_o_Stationary_matrix2_5_7(my_stationary_io_o_Stationary_matrix2_5_7),
    .io_o_Stationary_matrix2_6_0(my_stationary_io_o_Stationary_matrix2_6_0),
    .io_o_Stationary_matrix2_6_1(my_stationary_io_o_Stationary_matrix2_6_1),
    .io_o_Stationary_matrix2_6_2(my_stationary_io_o_Stationary_matrix2_6_2),
    .io_o_Stationary_matrix2_6_3(my_stationary_io_o_Stationary_matrix2_6_3),
    .io_o_Stationary_matrix2_6_4(my_stationary_io_o_Stationary_matrix2_6_4),
    .io_o_Stationary_matrix2_6_5(my_stationary_io_o_Stationary_matrix2_6_5),
    .io_o_Stationary_matrix2_6_6(my_stationary_io_o_Stationary_matrix2_6_6),
    .io_o_Stationary_matrix2_6_7(my_stationary_io_o_Stationary_matrix2_6_7),
    .io_o_Stationary_matrix2_7_0(my_stationary_io_o_Stationary_matrix2_7_0),
    .io_o_Stationary_matrix2_7_1(my_stationary_io_o_Stationary_matrix2_7_1),
    .io_o_Stationary_matrix2_7_2(my_stationary_io_o_Stationary_matrix2_7_2),
    .io_o_Stationary_matrix2_7_3(my_stationary_io_o_Stationary_matrix2_7_3),
    .io_o_Stationary_matrix2_7_4(my_stationary_io_o_Stationary_matrix2_7_4),
    .io_o_Stationary_matrix2_7_5(my_stationary_io_o_Stationary_matrix2_7_5),
    .io_o_Stationary_matrix2_7_6(my_stationary_io_o_Stationary_matrix2_7_6),
    .io_o_Stationary_matrix2_7_7(my_stationary_io_o_Stationary_matrix2_7_7),
    .io_o_Stationary_matrix3_0_0(my_stationary_io_o_Stationary_matrix3_0_0),
    .io_o_Stationary_matrix3_0_1(my_stationary_io_o_Stationary_matrix3_0_1),
    .io_o_Stationary_matrix3_0_2(my_stationary_io_o_Stationary_matrix3_0_2),
    .io_o_Stationary_matrix3_0_3(my_stationary_io_o_Stationary_matrix3_0_3),
    .io_o_Stationary_matrix3_0_4(my_stationary_io_o_Stationary_matrix3_0_4),
    .io_o_Stationary_matrix3_0_5(my_stationary_io_o_Stationary_matrix3_0_5),
    .io_o_Stationary_matrix3_0_6(my_stationary_io_o_Stationary_matrix3_0_6),
    .io_o_Stationary_matrix3_0_7(my_stationary_io_o_Stationary_matrix3_0_7),
    .io_o_Stationary_matrix3_1_0(my_stationary_io_o_Stationary_matrix3_1_0),
    .io_o_Stationary_matrix3_1_1(my_stationary_io_o_Stationary_matrix3_1_1),
    .io_o_Stationary_matrix3_1_2(my_stationary_io_o_Stationary_matrix3_1_2),
    .io_o_Stationary_matrix3_1_3(my_stationary_io_o_Stationary_matrix3_1_3),
    .io_o_Stationary_matrix3_1_4(my_stationary_io_o_Stationary_matrix3_1_4),
    .io_o_Stationary_matrix3_1_5(my_stationary_io_o_Stationary_matrix3_1_5),
    .io_o_Stationary_matrix3_1_6(my_stationary_io_o_Stationary_matrix3_1_6),
    .io_o_Stationary_matrix3_1_7(my_stationary_io_o_Stationary_matrix3_1_7),
    .io_o_Stationary_matrix3_2_0(my_stationary_io_o_Stationary_matrix3_2_0),
    .io_o_Stationary_matrix3_2_1(my_stationary_io_o_Stationary_matrix3_2_1),
    .io_o_Stationary_matrix3_2_2(my_stationary_io_o_Stationary_matrix3_2_2),
    .io_o_Stationary_matrix3_2_3(my_stationary_io_o_Stationary_matrix3_2_3),
    .io_o_Stationary_matrix3_2_4(my_stationary_io_o_Stationary_matrix3_2_4),
    .io_o_Stationary_matrix3_2_5(my_stationary_io_o_Stationary_matrix3_2_5),
    .io_o_Stationary_matrix3_2_6(my_stationary_io_o_Stationary_matrix3_2_6),
    .io_o_Stationary_matrix3_2_7(my_stationary_io_o_Stationary_matrix3_2_7),
    .io_o_Stationary_matrix3_3_0(my_stationary_io_o_Stationary_matrix3_3_0),
    .io_o_Stationary_matrix3_3_1(my_stationary_io_o_Stationary_matrix3_3_1),
    .io_o_Stationary_matrix3_3_2(my_stationary_io_o_Stationary_matrix3_3_2),
    .io_o_Stationary_matrix3_3_3(my_stationary_io_o_Stationary_matrix3_3_3),
    .io_o_Stationary_matrix3_3_4(my_stationary_io_o_Stationary_matrix3_3_4),
    .io_o_Stationary_matrix3_3_5(my_stationary_io_o_Stationary_matrix3_3_5),
    .io_o_Stationary_matrix3_3_6(my_stationary_io_o_Stationary_matrix3_3_6),
    .io_o_Stationary_matrix3_3_7(my_stationary_io_o_Stationary_matrix3_3_7),
    .io_o_Stationary_matrix3_4_0(my_stationary_io_o_Stationary_matrix3_4_0),
    .io_o_Stationary_matrix3_4_1(my_stationary_io_o_Stationary_matrix3_4_1),
    .io_o_Stationary_matrix3_4_2(my_stationary_io_o_Stationary_matrix3_4_2),
    .io_o_Stationary_matrix3_4_3(my_stationary_io_o_Stationary_matrix3_4_3),
    .io_o_Stationary_matrix3_4_4(my_stationary_io_o_Stationary_matrix3_4_4),
    .io_o_Stationary_matrix3_4_5(my_stationary_io_o_Stationary_matrix3_4_5),
    .io_o_Stationary_matrix3_4_6(my_stationary_io_o_Stationary_matrix3_4_6),
    .io_o_Stationary_matrix3_4_7(my_stationary_io_o_Stationary_matrix3_4_7),
    .io_o_Stationary_matrix3_5_0(my_stationary_io_o_Stationary_matrix3_5_0),
    .io_o_Stationary_matrix3_5_1(my_stationary_io_o_Stationary_matrix3_5_1),
    .io_o_Stationary_matrix3_5_2(my_stationary_io_o_Stationary_matrix3_5_2),
    .io_o_Stationary_matrix3_5_3(my_stationary_io_o_Stationary_matrix3_5_3),
    .io_o_Stationary_matrix3_5_4(my_stationary_io_o_Stationary_matrix3_5_4),
    .io_o_Stationary_matrix3_5_5(my_stationary_io_o_Stationary_matrix3_5_5),
    .io_o_Stationary_matrix3_5_6(my_stationary_io_o_Stationary_matrix3_5_6),
    .io_o_Stationary_matrix3_5_7(my_stationary_io_o_Stationary_matrix3_5_7),
    .io_o_Stationary_matrix3_6_0(my_stationary_io_o_Stationary_matrix3_6_0),
    .io_o_Stationary_matrix3_6_1(my_stationary_io_o_Stationary_matrix3_6_1),
    .io_o_Stationary_matrix3_6_2(my_stationary_io_o_Stationary_matrix3_6_2),
    .io_o_Stationary_matrix3_6_3(my_stationary_io_o_Stationary_matrix3_6_3),
    .io_o_Stationary_matrix3_6_4(my_stationary_io_o_Stationary_matrix3_6_4),
    .io_o_Stationary_matrix3_6_5(my_stationary_io_o_Stationary_matrix3_6_5),
    .io_o_Stationary_matrix3_6_6(my_stationary_io_o_Stationary_matrix3_6_6),
    .io_o_Stationary_matrix3_6_7(my_stationary_io_o_Stationary_matrix3_6_7),
    .io_o_Stationary_matrix3_7_0(my_stationary_io_o_Stationary_matrix3_7_0),
    .io_o_Stationary_matrix3_7_1(my_stationary_io_o_Stationary_matrix3_7_1),
    .io_o_Stationary_matrix3_7_2(my_stationary_io_o_Stationary_matrix3_7_2),
    .io_o_Stationary_matrix3_7_3(my_stationary_io_o_Stationary_matrix3_7_3),
    .io_o_Stationary_matrix3_7_4(my_stationary_io_o_Stationary_matrix3_7_4),
    .io_o_Stationary_matrix3_7_5(my_stationary_io_o_Stationary_matrix3_7_5),
    .io_o_Stationary_matrix3_7_6(my_stationary_io_o_Stationary_matrix3_7_6),
    .io_o_Stationary_matrix3_7_7(my_stationary_io_o_Stationary_matrix3_7_7),
    .io_o_Stationary_matrix4_0_0(my_stationary_io_o_Stationary_matrix4_0_0),
    .io_o_Stationary_matrix4_0_1(my_stationary_io_o_Stationary_matrix4_0_1),
    .io_o_Stationary_matrix4_0_2(my_stationary_io_o_Stationary_matrix4_0_2),
    .io_o_Stationary_matrix4_0_3(my_stationary_io_o_Stationary_matrix4_0_3),
    .io_o_Stationary_matrix4_0_4(my_stationary_io_o_Stationary_matrix4_0_4),
    .io_o_Stationary_matrix4_0_5(my_stationary_io_o_Stationary_matrix4_0_5),
    .io_o_Stationary_matrix4_0_6(my_stationary_io_o_Stationary_matrix4_0_6),
    .io_o_Stationary_matrix4_0_7(my_stationary_io_o_Stationary_matrix4_0_7),
    .io_o_Stationary_matrix4_1_0(my_stationary_io_o_Stationary_matrix4_1_0),
    .io_o_Stationary_matrix4_1_1(my_stationary_io_o_Stationary_matrix4_1_1),
    .io_o_Stationary_matrix4_1_2(my_stationary_io_o_Stationary_matrix4_1_2),
    .io_o_Stationary_matrix4_1_3(my_stationary_io_o_Stationary_matrix4_1_3),
    .io_o_Stationary_matrix4_1_4(my_stationary_io_o_Stationary_matrix4_1_4),
    .io_o_Stationary_matrix4_1_5(my_stationary_io_o_Stationary_matrix4_1_5),
    .io_o_Stationary_matrix4_1_6(my_stationary_io_o_Stationary_matrix4_1_6),
    .io_o_Stationary_matrix4_1_7(my_stationary_io_o_Stationary_matrix4_1_7),
    .io_o_Stationary_matrix4_2_0(my_stationary_io_o_Stationary_matrix4_2_0),
    .io_o_Stationary_matrix4_2_1(my_stationary_io_o_Stationary_matrix4_2_1),
    .io_o_Stationary_matrix4_2_2(my_stationary_io_o_Stationary_matrix4_2_2),
    .io_o_Stationary_matrix4_2_3(my_stationary_io_o_Stationary_matrix4_2_3),
    .io_o_Stationary_matrix4_2_4(my_stationary_io_o_Stationary_matrix4_2_4),
    .io_o_Stationary_matrix4_2_5(my_stationary_io_o_Stationary_matrix4_2_5),
    .io_o_Stationary_matrix4_2_6(my_stationary_io_o_Stationary_matrix4_2_6),
    .io_o_Stationary_matrix4_2_7(my_stationary_io_o_Stationary_matrix4_2_7),
    .io_o_Stationary_matrix4_3_0(my_stationary_io_o_Stationary_matrix4_3_0),
    .io_o_Stationary_matrix4_3_1(my_stationary_io_o_Stationary_matrix4_3_1),
    .io_o_Stationary_matrix4_3_2(my_stationary_io_o_Stationary_matrix4_3_2),
    .io_o_Stationary_matrix4_3_3(my_stationary_io_o_Stationary_matrix4_3_3),
    .io_o_Stationary_matrix4_3_4(my_stationary_io_o_Stationary_matrix4_3_4),
    .io_o_Stationary_matrix4_3_5(my_stationary_io_o_Stationary_matrix4_3_5),
    .io_o_Stationary_matrix4_3_6(my_stationary_io_o_Stationary_matrix4_3_6),
    .io_o_Stationary_matrix4_3_7(my_stationary_io_o_Stationary_matrix4_3_7),
    .io_o_Stationary_matrix4_4_0(my_stationary_io_o_Stationary_matrix4_4_0),
    .io_o_Stationary_matrix4_4_1(my_stationary_io_o_Stationary_matrix4_4_1),
    .io_o_Stationary_matrix4_4_2(my_stationary_io_o_Stationary_matrix4_4_2),
    .io_o_Stationary_matrix4_4_3(my_stationary_io_o_Stationary_matrix4_4_3),
    .io_o_Stationary_matrix4_4_4(my_stationary_io_o_Stationary_matrix4_4_4),
    .io_o_Stationary_matrix4_4_5(my_stationary_io_o_Stationary_matrix4_4_5),
    .io_o_Stationary_matrix4_4_6(my_stationary_io_o_Stationary_matrix4_4_6),
    .io_o_Stationary_matrix4_4_7(my_stationary_io_o_Stationary_matrix4_4_7),
    .io_o_Stationary_matrix4_5_0(my_stationary_io_o_Stationary_matrix4_5_0),
    .io_o_Stationary_matrix4_5_1(my_stationary_io_o_Stationary_matrix4_5_1),
    .io_o_Stationary_matrix4_5_2(my_stationary_io_o_Stationary_matrix4_5_2),
    .io_o_Stationary_matrix4_5_3(my_stationary_io_o_Stationary_matrix4_5_3),
    .io_o_Stationary_matrix4_5_4(my_stationary_io_o_Stationary_matrix4_5_4),
    .io_o_Stationary_matrix4_5_5(my_stationary_io_o_Stationary_matrix4_5_5),
    .io_o_Stationary_matrix4_5_6(my_stationary_io_o_Stationary_matrix4_5_6),
    .io_o_Stationary_matrix4_5_7(my_stationary_io_o_Stationary_matrix4_5_7),
    .io_o_Stationary_matrix4_6_0(my_stationary_io_o_Stationary_matrix4_6_0),
    .io_o_Stationary_matrix4_6_1(my_stationary_io_o_Stationary_matrix4_6_1),
    .io_o_Stationary_matrix4_6_2(my_stationary_io_o_Stationary_matrix4_6_2),
    .io_o_Stationary_matrix4_6_3(my_stationary_io_o_Stationary_matrix4_6_3),
    .io_o_Stationary_matrix4_6_4(my_stationary_io_o_Stationary_matrix4_6_4),
    .io_o_Stationary_matrix4_6_5(my_stationary_io_o_Stationary_matrix4_6_5),
    .io_o_Stationary_matrix4_6_6(my_stationary_io_o_Stationary_matrix4_6_6),
    .io_o_Stationary_matrix4_6_7(my_stationary_io_o_Stationary_matrix4_6_7),
    .io_o_Stationary_matrix4_7_0(my_stationary_io_o_Stationary_matrix4_7_0),
    .io_o_Stationary_matrix4_7_1(my_stationary_io_o_Stationary_matrix4_7_1),
    .io_o_Stationary_matrix4_7_2(my_stationary_io_o_Stationary_matrix4_7_2),
    .io_o_Stationary_matrix4_7_3(my_stationary_io_o_Stationary_matrix4_7_3),
    .io_o_Stationary_matrix4_7_4(my_stationary_io_o_Stationary_matrix4_7_4),
    .io_o_Stationary_matrix4_7_5(my_stationary_io_o_Stationary_matrix4_7_5),
    .io_o_Stationary_matrix4_7_6(my_stationary_io_o_Stationary_matrix4_7_6),
    .io_o_Stationary_matrix4_7_7(my_stationary_io_o_Stationary_matrix4_7_7),
    .io_o_Stationary_matrix5_0_0(my_stationary_io_o_Stationary_matrix5_0_0),
    .io_o_Stationary_matrix5_0_1(my_stationary_io_o_Stationary_matrix5_0_1),
    .io_o_Stationary_matrix5_0_2(my_stationary_io_o_Stationary_matrix5_0_2),
    .io_o_Stationary_matrix5_0_3(my_stationary_io_o_Stationary_matrix5_0_3),
    .io_o_Stationary_matrix5_0_4(my_stationary_io_o_Stationary_matrix5_0_4),
    .io_o_Stationary_matrix5_0_5(my_stationary_io_o_Stationary_matrix5_0_5),
    .io_o_Stationary_matrix5_0_6(my_stationary_io_o_Stationary_matrix5_0_6),
    .io_o_Stationary_matrix5_0_7(my_stationary_io_o_Stationary_matrix5_0_7),
    .io_o_Stationary_matrix5_1_0(my_stationary_io_o_Stationary_matrix5_1_0),
    .io_o_Stationary_matrix5_1_1(my_stationary_io_o_Stationary_matrix5_1_1),
    .io_o_Stationary_matrix5_1_2(my_stationary_io_o_Stationary_matrix5_1_2),
    .io_o_Stationary_matrix5_1_3(my_stationary_io_o_Stationary_matrix5_1_3),
    .io_o_Stationary_matrix5_1_4(my_stationary_io_o_Stationary_matrix5_1_4),
    .io_o_Stationary_matrix5_1_5(my_stationary_io_o_Stationary_matrix5_1_5),
    .io_o_Stationary_matrix5_1_6(my_stationary_io_o_Stationary_matrix5_1_6),
    .io_o_Stationary_matrix5_1_7(my_stationary_io_o_Stationary_matrix5_1_7),
    .io_o_Stationary_matrix5_2_0(my_stationary_io_o_Stationary_matrix5_2_0),
    .io_o_Stationary_matrix5_2_1(my_stationary_io_o_Stationary_matrix5_2_1),
    .io_o_Stationary_matrix5_2_2(my_stationary_io_o_Stationary_matrix5_2_2),
    .io_o_Stationary_matrix5_2_3(my_stationary_io_o_Stationary_matrix5_2_3),
    .io_o_Stationary_matrix5_2_4(my_stationary_io_o_Stationary_matrix5_2_4),
    .io_o_Stationary_matrix5_2_5(my_stationary_io_o_Stationary_matrix5_2_5),
    .io_o_Stationary_matrix5_2_6(my_stationary_io_o_Stationary_matrix5_2_6),
    .io_o_Stationary_matrix5_2_7(my_stationary_io_o_Stationary_matrix5_2_7),
    .io_o_Stationary_matrix5_3_0(my_stationary_io_o_Stationary_matrix5_3_0),
    .io_o_Stationary_matrix5_3_1(my_stationary_io_o_Stationary_matrix5_3_1),
    .io_o_Stationary_matrix5_3_2(my_stationary_io_o_Stationary_matrix5_3_2),
    .io_o_Stationary_matrix5_3_3(my_stationary_io_o_Stationary_matrix5_3_3),
    .io_o_Stationary_matrix5_3_4(my_stationary_io_o_Stationary_matrix5_3_4),
    .io_o_Stationary_matrix5_3_5(my_stationary_io_o_Stationary_matrix5_3_5),
    .io_o_Stationary_matrix5_3_6(my_stationary_io_o_Stationary_matrix5_3_6),
    .io_o_Stationary_matrix5_3_7(my_stationary_io_o_Stationary_matrix5_3_7),
    .io_o_Stationary_matrix5_4_0(my_stationary_io_o_Stationary_matrix5_4_0),
    .io_o_Stationary_matrix5_4_1(my_stationary_io_o_Stationary_matrix5_4_1),
    .io_o_Stationary_matrix5_4_2(my_stationary_io_o_Stationary_matrix5_4_2),
    .io_o_Stationary_matrix5_4_3(my_stationary_io_o_Stationary_matrix5_4_3),
    .io_o_Stationary_matrix5_4_4(my_stationary_io_o_Stationary_matrix5_4_4),
    .io_o_Stationary_matrix5_4_5(my_stationary_io_o_Stationary_matrix5_4_5),
    .io_o_Stationary_matrix5_4_6(my_stationary_io_o_Stationary_matrix5_4_6),
    .io_o_Stationary_matrix5_4_7(my_stationary_io_o_Stationary_matrix5_4_7),
    .io_o_Stationary_matrix5_5_0(my_stationary_io_o_Stationary_matrix5_5_0),
    .io_o_Stationary_matrix5_5_1(my_stationary_io_o_Stationary_matrix5_5_1),
    .io_o_Stationary_matrix5_5_2(my_stationary_io_o_Stationary_matrix5_5_2),
    .io_o_Stationary_matrix5_5_3(my_stationary_io_o_Stationary_matrix5_5_3),
    .io_o_Stationary_matrix5_5_4(my_stationary_io_o_Stationary_matrix5_5_4),
    .io_o_Stationary_matrix5_5_5(my_stationary_io_o_Stationary_matrix5_5_5),
    .io_o_Stationary_matrix5_5_6(my_stationary_io_o_Stationary_matrix5_5_6),
    .io_o_Stationary_matrix5_5_7(my_stationary_io_o_Stationary_matrix5_5_7),
    .io_o_Stationary_matrix5_6_0(my_stationary_io_o_Stationary_matrix5_6_0),
    .io_o_Stationary_matrix5_6_1(my_stationary_io_o_Stationary_matrix5_6_1),
    .io_o_Stationary_matrix5_6_2(my_stationary_io_o_Stationary_matrix5_6_2),
    .io_o_Stationary_matrix5_6_3(my_stationary_io_o_Stationary_matrix5_6_3),
    .io_o_Stationary_matrix5_6_4(my_stationary_io_o_Stationary_matrix5_6_4),
    .io_o_Stationary_matrix5_6_5(my_stationary_io_o_Stationary_matrix5_6_5),
    .io_o_Stationary_matrix5_6_6(my_stationary_io_o_Stationary_matrix5_6_6),
    .io_o_Stationary_matrix5_6_7(my_stationary_io_o_Stationary_matrix5_6_7),
    .io_o_Stationary_matrix5_7_0(my_stationary_io_o_Stationary_matrix5_7_0),
    .io_o_Stationary_matrix5_7_1(my_stationary_io_o_Stationary_matrix5_7_1),
    .io_o_Stationary_matrix5_7_2(my_stationary_io_o_Stationary_matrix5_7_2),
    .io_o_Stationary_matrix5_7_3(my_stationary_io_o_Stationary_matrix5_7_3),
    .io_o_Stationary_matrix5_7_4(my_stationary_io_o_Stationary_matrix5_7_4),
    .io_o_Stationary_matrix5_7_5(my_stationary_io_o_Stationary_matrix5_7_5),
    .io_o_Stationary_matrix5_7_6(my_stationary_io_o_Stationary_matrix5_7_6),
    .io_o_Stationary_matrix5_7_7(my_stationary_io_o_Stationary_matrix5_7_7),
    .io_o_Stationary_matrix6_0_0(my_stationary_io_o_Stationary_matrix6_0_0),
    .io_o_Stationary_matrix6_0_1(my_stationary_io_o_Stationary_matrix6_0_1),
    .io_o_Stationary_matrix6_0_2(my_stationary_io_o_Stationary_matrix6_0_2),
    .io_o_Stationary_matrix6_0_3(my_stationary_io_o_Stationary_matrix6_0_3),
    .io_o_Stationary_matrix6_0_4(my_stationary_io_o_Stationary_matrix6_0_4),
    .io_o_Stationary_matrix6_0_5(my_stationary_io_o_Stationary_matrix6_0_5),
    .io_o_Stationary_matrix6_0_6(my_stationary_io_o_Stationary_matrix6_0_6),
    .io_o_Stationary_matrix6_0_7(my_stationary_io_o_Stationary_matrix6_0_7),
    .io_o_Stationary_matrix6_1_0(my_stationary_io_o_Stationary_matrix6_1_0),
    .io_o_Stationary_matrix6_1_1(my_stationary_io_o_Stationary_matrix6_1_1),
    .io_o_Stationary_matrix6_1_2(my_stationary_io_o_Stationary_matrix6_1_2),
    .io_o_Stationary_matrix6_1_3(my_stationary_io_o_Stationary_matrix6_1_3),
    .io_o_Stationary_matrix6_1_4(my_stationary_io_o_Stationary_matrix6_1_4),
    .io_o_Stationary_matrix6_1_5(my_stationary_io_o_Stationary_matrix6_1_5),
    .io_o_Stationary_matrix6_1_6(my_stationary_io_o_Stationary_matrix6_1_6),
    .io_o_Stationary_matrix6_1_7(my_stationary_io_o_Stationary_matrix6_1_7),
    .io_o_Stationary_matrix6_2_0(my_stationary_io_o_Stationary_matrix6_2_0),
    .io_o_Stationary_matrix6_2_1(my_stationary_io_o_Stationary_matrix6_2_1),
    .io_o_Stationary_matrix6_2_2(my_stationary_io_o_Stationary_matrix6_2_2),
    .io_o_Stationary_matrix6_2_3(my_stationary_io_o_Stationary_matrix6_2_3),
    .io_o_Stationary_matrix6_2_4(my_stationary_io_o_Stationary_matrix6_2_4),
    .io_o_Stationary_matrix6_2_5(my_stationary_io_o_Stationary_matrix6_2_5),
    .io_o_Stationary_matrix6_2_6(my_stationary_io_o_Stationary_matrix6_2_6),
    .io_o_Stationary_matrix6_2_7(my_stationary_io_o_Stationary_matrix6_2_7),
    .io_o_Stationary_matrix6_3_0(my_stationary_io_o_Stationary_matrix6_3_0),
    .io_o_Stationary_matrix6_3_1(my_stationary_io_o_Stationary_matrix6_3_1),
    .io_o_Stationary_matrix6_3_2(my_stationary_io_o_Stationary_matrix6_3_2),
    .io_o_Stationary_matrix6_3_3(my_stationary_io_o_Stationary_matrix6_3_3),
    .io_o_Stationary_matrix6_3_4(my_stationary_io_o_Stationary_matrix6_3_4),
    .io_o_Stationary_matrix6_3_5(my_stationary_io_o_Stationary_matrix6_3_5),
    .io_o_Stationary_matrix6_3_6(my_stationary_io_o_Stationary_matrix6_3_6),
    .io_o_Stationary_matrix6_3_7(my_stationary_io_o_Stationary_matrix6_3_7),
    .io_o_Stationary_matrix6_4_0(my_stationary_io_o_Stationary_matrix6_4_0),
    .io_o_Stationary_matrix6_4_1(my_stationary_io_o_Stationary_matrix6_4_1),
    .io_o_Stationary_matrix6_4_2(my_stationary_io_o_Stationary_matrix6_4_2),
    .io_o_Stationary_matrix6_4_3(my_stationary_io_o_Stationary_matrix6_4_3),
    .io_o_Stationary_matrix6_4_4(my_stationary_io_o_Stationary_matrix6_4_4),
    .io_o_Stationary_matrix6_4_5(my_stationary_io_o_Stationary_matrix6_4_5),
    .io_o_Stationary_matrix6_4_6(my_stationary_io_o_Stationary_matrix6_4_6),
    .io_o_Stationary_matrix6_4_7(my_stationary_io_o_Stationary_matrix6_4_7),
    .io_o_Stationary_matrix6_5_0(my_stationary_io_o_Stationary_matrix6_5_0),
    .io_o_Stationary_matrix6_5_1(my_stationary_io_o_Stationary_matrix6_5_1),
    .io_o_Stationary_matrix6_5_2(my_stationary_io_o_Stationary_matrix6_5_2),
    .io_o_Stationary_matrix6_5_3(my_stationary_io_o_Stationary_matrix6_5_3),
    .io_o_Stationary_matrix6_5_4(my_stationary_io_o_Stationary_matrix6_5_4),
    .io_o_Stationary_matrix6_5_5(my_stationary_io_o_Stationary_matrix6_5_5),
    .io_o_Stationary_matrix6_5_6(my_stationary_io_o_Stationary_matrix6_5_6),
    .io_o_Stationary_matrix6_5_7(my_stationary_io_o_Stationary_matrix6_5_7),
    .io_o_Stationary_matrix6_6_0(my_stationary_io_o_Stationary_matrix6_6_0),
    .io_o_Stationary_matrix6_6_1(my_stationary_io_o_Stationary_matrix6_6_1),
    .io_o_Stationary_matrix6_6_2(my_stationary_io_o_Stationary_matrix6_6_2),
    .io_o_Stationary_matrix6_6_3(my_stationary_io_o_Stationary_matrix6_6_3),
    .io_o_Stationary_matrix6_6_4(my_stationary_io_o_Stationary_matrix6_6_4),
    .io_o_Stationary_matrix6_6_5(my_stationary_io_o_Stationary_matrix6_6_5),
    .io_o_Stationary_matrix6_6_6(my_stationary_io_o_Stationary_matrix6_6_6),
    .io_o_Stationary_matrix6_6_7(my_stationary_io_o_Stationary_matrix6_6_7),
    .io_o_Stationary_matrix6_7_0(my_stationary_io_o_Stationary_matrix6_7_0),
    .io_o_Stationary_matrix6_7_1(my_stationary_io_o_Stationary_matrix6_7_1),
    .io_o_Stationary_matrix6_7_2(my_stationary_io_o_Stationary_matrix6_7_2),
    .io_o_Stationary_matrix6_7_3(my_stationary_io_o_Stationary_matrix6_7_3),
    .io_o_Stationary_matrix6_7_4(my_stationary_io_o_Stationary_matrix6_7_4),
    .io_o_Stationary_matrix6_7_5(my_stationary_io_o_Stationary_matrix6_7_5),
    .io_o_Stationary_matrix6_7_6(my_stationary_io_o_Stationary_matrix6_7_6),
    .io_o_Stationary_matrix6_7_7(my_stationary_io_o_Stationary_matrix6_7_7),
    .io_o_Stationary_matrix7_0_0(my_stationary_io_o_Stationary_matrix7_0_0),
    .io_o_Stationary_matrix7_0_1(my_stationary_io_o_Stationary_matrix7_0_1),
    .io_o_Stationary_matrix7_0_2(my_stationary_io_o_Stationary_matrix7_0_2),
    .io_o_Stationary_matrix7_0_3(my_stationary_io_o_Stationary_matrix7_0_3),
    .io_o_Stationary_matrix7_0_4(my_stationary_io_o_Stationary_matrix7_0_4),
    .io_o_Stationary_matrix7_0_5(my_stationary_io_o_Stationary_matrix7_0_5),
    .io_o_Stationary_matrix7_0_6(my_stationary_io_o_Stationary_matrix7_0_6),
    .io_o_Stationary_matrix7_0_7(my_stationary_io_o_Stationary_matrix7_0_7),
    .io_o_Stationary_matrix7_1_0(my_stationary_io_o_Stationary_matrix7_1_0),
    .io_o_Stationary_matrix7_1_1(my_stationary_io_o_Stationary_matrix7_1_1),
    .io_o_Stationary_matrix7_1_2(my_stationary_io_o_Stationary_matrix7_1_2),
    .io_o_Stationary_matrix7_1_3(my_stationary_io_o_Stationary_matrix7_1_3),
    .io_o_Stationary_matrix7_1_4(my_stationary_io_o_Stationary_matrix7_1_4),
    .io_o_Stationary_matrix7_1_5(my_stationary_io_o_Stationary_matrix7_1_5),
    .io_o_Stationary_matrix7_1_6(my_stationary_io_o_Stationary_matrix7_1_6),
    .io_o_Stationary_matrix7_1_7(my_stationary_io_o_Stationary_matrix7_1_7),
    .io_o_Stationary_matrix7_2_0(my_stationary_io_o_Stationary_matrix7_2_0),
    .io_o_Stationary_matrix7_2_1(my_stationary_io_o_Stationary_matrix7_2_1),
    .io_o_Stationary_matrix7_2_2(my_stationary_io_o_Stationary_matrix7_2_2),
    .io_o_Stationary_matrix7_2_3(my_stationary_io_o_Stationary_matrix7_2_3),
    .io_o_Stationary_matrix7_2_4(my_stationary_io_o_Stationary_matrix7_2_4),
    .io_o_Stationary_matrix7_2_5(my_stationary_io_o_Stationary_matrix7_2_5),
    .io_o_Stationary_matrix7_2_6(my_stationary_io_o_Stationary_matrix7_2_6),
    .io_o_Stationary_matrix7_2_7(my_stationary_io_o_Stationary_matrix7_2_7),
    .io_o_Stationary_matrix7_3_0(my_stationary_io_o_Stationary_matrix7_3_0),
    .io_o_Stationary_matrix7_3_1(my_stationary_io_o_Stationary_matrix7_3_1),
    .io_o_Stationary_matrix7_3_2(my_stationary_io_o_Stationary_matrix7_3_2),
    .io_o_Stationary_matrix7_3_3(my_stationary_io_o_Stationary_matrix7_3_3),
    .io_o_Stationary_matrix7_3_4(my_stationary_io_o_Stationary_matrix7_3_4),
    .io_o_Stationary_matrix7_3_5(my_stationary_io_o_Stationary_matrix7_3_5),
    .io_o_Stationary_matrix7_3_6(my_stationary_io_o_Stationary_matrix7_3_6),
    .io_o_Stationary_matrix7_3_7(my_stationary_io_o_Stationary_matrix7_3_7),
    .io_o_Stationary_matrix7_4_0(my_stationary_io_o_Stationary_matrix7_4_0),
    .io_o_Stationary_matrix7_4_1(my_stationary_io_o_Stationary_matrix7_4_1),
    .io_o_Stationary_matrix7_4_2(my_stationary_io_o_Stationary_matrix7_4_2),
    .io_o_Stationary_matrix7_4_3(my_stationary_io_o_Stationary_matrix7_4_3),
    .io_o_Stationary_matrix7_4_4(my_stationary_io_o_Stationary_matrix7_4_4),
    .io_o_Stationary_matrix7_4_5(my_stationary_io_o_Stationary_matrix7_4_5),
    .io_o_Stationary_matrix7_4_6(my_stationary_io_o_Stationary_matrix7_4_6),
    .io_o_Stationary_matrix7_4_7(my_stationary_io_o_Stationary_matrix7_4_7),
    .io_o_Stationary_matrix7_5_0(my_stationary_io_o_Stationary_matrix7_5_0),
    .io_o_Stationary_matrix7_5_1(my_stationary_io_o_Stationary_matrix7_5_1),
    .io_o_Stationary_matrix7_5_2(my_stationary_io_o_Stationary_matrix7_5_2),
    .io_o_Stationary_matrix7_5_3(my_stationary_io_o_Stationary_matrix7_5_3),
    .io_o_Stationary_matrix7_5_4(my_stationary_io_o_Stationary_matrix7_5_4),
    .io_o_Stationary_matrix7_5_5(my_stationary_io_o_Stationary_matrix7_5_5),
    .io_o_Stationary_matrix7_5_6(my_stationary_io_o_Stationary_matrix7_5_6),
    .io_o_Stationary_matrix7_5_7(my_stationary_io_o_Stationary_matrix7_5_7),
    .io_o_Stationary_matrix7_6_0(my_stationary_io_o_Stationary_matrix7_6_0),
    .io_o_Stationary_matrix7_6_1(my_stationary_io_o_Stationary_matrix7_6_1),
    .io_o_Stationary_matrix7_6_2(my_stationary_io_o_Stationary_matrix7_6_2),
    .io_o_Stationary_matrix7_6_3(my_stationary_io_o_Stationary_matrix7_6_3),
    .io_o_Stationary_matrix7_6_4(my_stationary_io_o_Stationary_matrix7_6_4),
    .io_o_Stationary_matrix7_6_5(my_stationary_io_o_Stationary_matrix7_6_5),
    .io_o_Stationary_matrix7_6_6(my_stationary_io_o_Stationary_matrix7_6_6),
    .io_o_Stationary_matrix7_6_7(my_stationary_io_o_Stationary_matrix7_6_7),
    .io_o_Stationary_matrix7_7_0(my_stationary_io_o_Stationary_matrix7_7_0),
    .io_o_Stationary_matrix7_7_1(my_stationary_io_o_Stationary_matrix7_7_1),
    .io_o_Stationary_matrix7_7_2(my_stationary_io_o_Stationary_matrix7_7_2),
    .io_o_Stationary_matrix7_7_3(my_stationary_io_o_Stationary_matrix7_7_3),
    .io_o_Stationary_matrix7_7_4(my_stationary_io_o_Stationary_matrix7_7_4),
    .io_o_Stationary_matrix7_7_5(my_stationary_io_o_Stationary_matrix7_7_5),
    .io_o_Stationary_matrix7_7_6(my_stationary_io_o_Stationary_matrix7_7_6),
    .io_o_Stationary_matrix7_7_7(my_stationary_io_o_Stationary_matrix7_7_7),
    .io_o_Stationary_matrix8_0_0(my_stationary_io_o_Stationary_matrix8_0_0),
    .io_o_Stationary_matrix8_0_1(my_stationary_io_o_Stationary_matrix8_0_1),
    .io_o_Stationary_matrix8_0_2(my_stationary_io_o_Stationary_matrix8_0_2),
    .io_o_Stationary_matrix8_0_3(my_stationary_io_o_Stationary_matrix8_0_3),
    .io_o_Stationary_matrix8_0_4(my_stationary_io_o_Stationary_matrix8_0_4),
    .io_o_Stationary_matrix8_0_5(my_stationary_io_o_Stationary_matrix8_0_5),
    .io_o_Stationary_matrix8_0_6(my_stationary_io_o_Stationary_matrix8_0_6),
    .io_o_Stationary_matrix8_0_7(my_stationary_io_o_Stationary_matrix8_0_7),
    .io_o_Stationary_matrix8_1_0(my_stationary_io_o_Stationary_matrix8_1_0),
    .io_o_Stationary_matrix8_1_1(my_stationary_io_o_Stationary_matrix8_1_1),
    .io_o_Stationary_matrix8_1_2(my_stationary_io_o_Stationary_matrix8_1_2),
    .io_o_Stationary_matrix8_1_3(my_stationary_io_o_Stationary_matrix8_1_3),
    .io_o_Stationary_matrix8_1_4(my_stationary_io_o_Stationary_matrix8_1_4),
    .io_o_Stationary_matrix8_1_5(my_stationary_io_o_Stationary_matrix8_1_5),
    .io_o_Stationary_matrix8_1_6(my_stationary_io_o_Stationary_matrix8_1_6),
    .io_o_Stationary_matrix8_1_7(my_stationary_io_o_Stationary_matrix8_1_7),
    .io_o_Stationary_matrix8_2_0(my_stationary_io_o_Stationary_matrix8_2_0),
    .io_o_Stationary_matrix8_2_1(my_stationary_io_o_Stationary_matrix8_2_1),
    .io_o_Stationary_matrix8_2_2(my_stationary_io_o_Stationary_matrix8_2_2),
    .io_o_Stationary_matrix8_2_3(my_stationary_io_o_Stationary_matrix8_2_3),
    .io_o_Stationary_matrix8_2_4(my_stationary_io_o_Stationary_matrix8_2_4),
    .io_o_Stationary_matrix8_2_5(my_stationary_io_o_Stationary_matrix8_2_5),
    .io_o_Stationary_matrix8_2_6(my_stationary_io_o_Stationary_matrix8_2_6),
    .io_o_Stationary_matrix8_2_7(my_stationary_io_o_Stationary_matrix8_2_7),
    .io_o_Stationary_matrix8_3_0(my_stationary_io_o_Stationary_matrix8_3_0),
    .io_o_Stationary_matrix8_3_1(my_stationary_io_o_Stationary_matrix8_3_1),
    .io_o_Stationary_matrix8_3_2(my_stationary_io_o_Stationary_matrix8_3_2),
    .io_o_Stationary_matrix8_3_3(my_stationary_io_o_Stationary_matrix8_3_3),
    .io_o_Stationary_matrix8_3_4(my_stationary_io_o_Stationary_matrix8_3_4),
    .io_o_Stationary_matrix8_3_5(my_stationary_io_o_Stationary_matrix8_3_5),
    .io_o_Stationary_matrix8_3_6(my_stationary_io_o_Stationary_matrix8_3_6),
    .io_o_Stationary_matrix8_3_7(my_stationary_io_o_Stationary_matrix8_3_7),
    .io_o_Stationary_matrix8_4_0(my_stationary_io_o_Stationary_matrix8_4_0),
    .io_o_Stationary_matrix8_4_1(my_stationary_io_o_Stationary_matrix8_4_1),
    .io_o_Stationary_matrix8_4_2(my_stationary_io_o_Stationary_matrix8_4_2),
    .io_o_Stationary_matrix8_4_3(my_stationary_io_o_Stationary_matrix8_4_3),
    .io_o_Stationary_matrix8_4_4(my_stationary_io_o_Stationary_matrix8_4_4),
    .io_o_Stationary_matrix8_4_5(my_stationary_io_o_Stationary_matrix8_4_5),
    .io_o_Stationary_matrix8_4_6(my_stationary_io_o_Stationary_matrix8_4_6),
    .io_o_Stationary_matrix8_4_7(my_stationary_io_o_Stationary_matrix8_4_7),
    .io_o_Stationary_matrix8_5_0(my_stationary_io_o_Stationary_matrix8_5_0),
    .io_o_Stationary_matrix8_5_1(my_stationary_io_o_Stationary_matrix8_5_1),
    .io_o_Stationary_matrix8_5_2(my_stationary_io_o_Stationary_matrix8_5_2),
    .io_o_Stationary_matrix8_5_3(my_stationary_io_o_Stationary_matrix8_5_3),
    .io_o_Stationary_matrix8_5_4(my_stationary_io_o_Stationary_matrix8_5_4),
    .io_o_Stationary_matrix8_5_5(my_stationary_io_o_Stationary_matrix8_5_5),
    .io_o_Stationary_matrix8_5_6(my_stationary_io_o_Stationary_matrix8_5_6),
    .io_o_Stationary_matrix8_5_7(my_stationary_io_o_Stationary_matrix8_5_7),
    .io_o_Stationary_matrix8_6_0(my_stationary_io_o_Stationary_matrix8_6_0),
    .io_o_Stationary_matrix8_6_1(my_stationary_io_o_Stationary_matrix8_6_1),
    .io_o_Stationary_matrix8_6_2(my_stationary_io_o_Stationary_matrix8_6_2),
    .io_o_Stationary_matrix8_6_3(my_stationary_io_o_Stationary_matrix8_6_3),
    .io_o_Stationary_matrix8_6_4(my_stationary_io_o_Stationary_matrix8_6_4),
    .io_o_Stationary_matrix8_6_5(my_stationary_io_o_Stationary_matrix8_6_5),
    .io_o_Stationary_matrix8_6_6(my_stationary_io_o_Stationary_matrix8_6_6),
    .io_o_Stationary_matrix8_6_7(my_stationary_io_o_Stationary_matrix8_6_7),
    .io_o_Stationary_matrix8_7_0(my_stationary_io_o_Stationary_matrix8_7_0),
    .io_o_Stationary_matrix8_7_1(my_stationary_io_o_Stationary_matrix8_7_1),
    .io_o_Stationary_matrix8_7_2(my_stationary_io_o_Stationary_matrix8_7_2),
    .io_o_Stationary_matrix8_7_3(my_stationary_io_o_Stationary_matrix8_7_3),
    .io_o_Stationary_matrix8_7_4(my_stationary_io_o_Stationary_matrix8_7_4),
    .io_o_Stationary_matrix8_7_5(my_stationary_io_o_Stationary_matrix8_7_5),
    .io_o_Stationary_matrix8_7_6(my_stationary_io_o_Stationary_matrix8_7_6),
    .io_o_Stationary_matrix8_7_7(my_stationary_io_o_Stationary_matrix8_7_7)
  );
  ivncontrol4 my_ivn1 ( // @[ivntop.scala 32:24]
    .clock(my_ivn1_clock),
    .reset(my_ivn1_reset),
    .io_Stationary_matrix_0_0(my_ivn1_io_Stationary_matrix_0_0),
    .io_Stationary_matrix_0_1(my_ivn1_io_Stationary_matrix_0_1),
    .io_Stationary_matrix_0_2(my_ivn1_io_Stationary_matrix_0_2),
    .io_Stationary_matrix_0_3(my_ivn1_io_Stationary_matrix_0_3),
    .io_Stationary_matrix_0_4(my_ivn1_io_Stationary_matrix_0_4),
    .io_Stationary_matrix_0_5(my_ivn1_io_Stationary_matrix_0_5),
    .io_Stationary_matrix_0_6(my_ivn1_io_Stationary_matrix_0_6),
    .io_Stationary_matrix_0_7(my_ivn1_io_Stationary_matrix_0_7),
    .io_Stationary_matrix_1_0(my_ivn1_io_Stationary_matrix_1_0),
    .io_Stationary_matrix_1_1(my_ivn1_io_Stationary_matrix_1_1),
    .io_Stationary_matrix_1_2(my_ivn1_io_Stationary_matrix_1_2),
    .io_Stationary_matrix_1_3(my_ivn1_io_Stationary_matrix_1_3),
    .io_Stationary_matrix_1_4(my_ivn1_io_Stationary_matrix_1_4),
    .io_Stationary_matrix_1_5(my_ivn1_io_Stationary_matrix_1_5),
    .io_Stationary_matrix_1_6(my_ivn1_io_Stationary_matrix_1_6),
    .io_Stationary_matrix_1_7(my_ivn1_io_Stationary_matrix_1_7),
    .io_Stationary_matrix_2_0(my_ivn1_io_Stationary_matrix_2_0),
    .io_Stationary_matrix_2_1(my_ivn1_io_Stationary_matrix_2_1),
    .io_Stationary_matrix_2_2(my_ivn1_io_Stationary_matrix_2_2),
    .io_Stationary_matrix_2_3(my_ivn1_io_Stationary_matrix_2_3),
    .io_Stationary_matrix_2_4(my_ivn1_io_Stationary_matrix_2_4),
    .io_Stationary_matrix_2_5(my_ivn1_io_Stationary_matrix_2_5),
    .io_Stationary_matrix_2_6(my_ivn1_io_Stationary_matrix_2_6),
    .io_Stationary_matrix_2_7(my_ivn1_io_Stationary_matrix_2_7),
    .io_Stationary_matrix_3_0(my_ivn1_io_Stationary_matrix_3_0),
    .io_Stationary_matrix_3_1(my_ivn1_io_Stationary_matrix_3_1),
    .io_Stationary_matrix_3_2(my_ivn1_io_Stationary_matrix_3_2),
    .io_Stationary_matrix_3_3(my_ivn1_io_Stationary_matrix_3_3),
    .io_Stationary_matrix_3_4(my_ivn1_io_Stationary_matrix_3_4),
    .io_Stationary_matrix_3_5(my_ivn1_io_Stationary_matrix_3_5),
    .io_Stationary_matrix_3_6(my_ivn1_io_Stationary_matrix_3_6),
    .io_Stationary_matrix_3_7(my_ivn1_io_Stationary_matrix_3_7),
    .io_Stationary_matrix_4_0(my_ivn1_io_Stationary_matrix_4_0),
    .io_Stationary_matrix_4_1(my_ivn1_io_Stationary_matrix_4_1),
    .io_Stationary_matrix_4_2(my_ivn1_io_Stationary_matrix_4_2),
    .io_Stationary_matrix_4_3(my_ivn1_io_Stationary_matrix_4_3),
    .io_Stationary_matrix_4_4(my_ivn1_io_Stationary_matrix_4_4),
    .io_Stationary_matrix_4_5(my_ivn1_io_Stationary_matrix_4_5),
    .io_Stationary_matrix_4_6(my_ivn1_io_Stationary_matrix_4_6),
    .io_Stationary_matrix_4_7(my_ivn1_io_Stationary_matrix_4_7),
    .io_Stationary_matrix_5_0(my_ivn1_io_Stationary_matrix_5_0),
    .io_Stationary_matrix_5_1(my_ivn1_io_Stationary_matrix_5_1),
    .io_Stationary_matrix_5_2(my_ivn1_io_Stationary_matrix_5_2),
    .io_Stationary_matrix_5_3(my_ivn1_io_Stationary_matrix_5_3),
    .io_Stationary_matrix_5_4(my_ivn1_io_Stationary_matrix_5_4),
    .io_Stationary_matrix_5_5(my_ivn1_io_Stationary_matrix_5_5),
    .io_Stationary_matrix_5_6(my_ivn1_io_Stationary_matrix_5_6),
    .io_Stationary_matrix_5_7(my_ivn1_io_Stationary_matrix_5_7),
    .io_Stationary_matrix_6_0(my_ivn1_io_Stationary_matrix_6_0),
    .io_Stationary_matrix_6_1(my_ivn1_io_Stationary_matrix_6_1),
    .io_Stationary_matrix_6_2(my_ivn1_io_Stationary_matrix_6_2),
    .io_Stationary_matrix_6_3(my_ivn1_io_Stationary_matrix_6_3),
    .io_Stationary_matrix_6_4(my_ivn1_io_Stationary_matrix_6_4),
    .io_Stationary_matrix_6_5(my_ivn1_io_Stationary_matrix_6_5),
    .io_Stationary_matrix_6_6(my_ivn1_io_Stationary_matrix_6_6),
    .io_Stationary_matrix_6_7(my_ivn1_io_Stationary_matrix_6_7),
    .io_Stationary_matrix_7_0(my_ivn1_io_Stationary_matrix_7_0),
    .io_Stationary_matrix_7_1(my_ivn1_io_Stationary_matrix_7_1),
    .io_Stationary_matrix_7_2(my_ivn1_io_Stationary_matrix_7_2),
    .io_Stationary_matrix_7_3(my_ivn1_io_Stationary_matrix_7_3),
    .io_Stationary_matrix_7_4(my_ivn1_io_Stationary_matrix_7_4),
    .io_Stationary_matrix_7_5(my_ivn1_io_Stationary_matrix_7_5),
    .io_Stationary_matrix_7_6(my_ivn1_io_Stationary_matrix_7_6),
    .io_Stationary_matrix_7_7(my_ivn1_io_Stationary_matrix_7_7),
    .io_o_vn_0(my_ivn1_io_o_vn_0),
    .io_o_vn_1(my_ivn1_io_o_vn_1),
    .io_o_vn_2(my_ivn1_io_o_vn_2),
    .io_o_vn_3(my_ivn1_io_o_vn_3),
    .io_o_vn2_0(my_ivn1_io_o_vn2_0),
    .io_o_vn2_1(my_ivn1_io_o_vn2_1),
    .io_o_vn2_2(my_ivn1_io_o_vn2_2),
    .io_o_vn2_3(my_ivn1_io_o_vn2_3),
    .io_ProcessValid(my_ivn1_io_ProcessValid)
  );
  ivncontrol4_1 my_ivn2 ( // @[ivntop.scala 40:24]
    .clock(my_ivn2_clock),
    .reset(my_ivn2_reset),
    .io_Stationary_matrix_0_0(my_ivn2_io_Stationary_matrix_0_0),
    .io_Stationary_matrix_0_1(my_ivn2_io_Stationary_matrix_0_1),
    .io_Stationary_matrix_0_2(my_ivn2_io_Stationary_matrix_0_2),
    .io_Stationary_matrix_0_3(my_ivn2_io_Stationary_matrix_0_3),
    .io_Stationary_matrix_0_4(my_ivn2_io_Stationary_matrix_0_4),
    .io_Stationary_matrix_0_5(my_ivn2_io_Stationary_matrix_0_5),
    .io_Stationary_matrix_0_6(my_ivn2_io_Stationary_matrix_0_6),
    .io_Stationary_matrix_0_7(my_ivn2_io_Stationary_matrix_0_7),
    .io_Stationary_matrix_1_0(my_ivn2_io_Stationary_matrix_1_0),
    .io_Stationary_matrix_1_1(my_ivn2_io_Stationary_matrix_1_1),
    .io_Stationary_matrix_1_2(my_ivn2_io_Stationary_matrix_1_2),
    .io_Stationary_matrix_1_3(my_ivn2_io_Stationary_matrix_1_3),
    .io_Stationary_matrix_1_4(my_ivn2_io_Stationary_matrix_1_4),
    .io_Stationary_matrix_1_5(my_ivn2_io_Stationary_matrix_1_5),
    .io_Stationary_matrix_1_6(my_ivn2_io_Stationary_matrix_1_6),
    .io_Stationary_matrix_1_7(my_ivn2_io_Stationary_matrix_1_7),
    .io_Stationary_matrix_2_0(my_ivn2_io_Stationary_matrix_2_0),
    .io_Stationary_matrix_2_1(my_ivn2_io_Stationary_matrix_2_1),
    .io_Stationary_matrix_2_2(my_ivn2_io_Stationary_matrix_2_2),
    .io_Stationary_matrix_2_3(my_ivn2_io_Stationary_matrix_2_3),
    .io_Stationary_matrix_2_4(my_ivn2_io_Stationary_matrix_2_4),
    .io_Stationary_matrix_2_5(my_ivn2_io_Stationary_matrix_2_5),
    .io_Stationary_matrix_2_6(my_ivn2_io_Stationary_matrix_2_6),
    .io_Stationary_matrix_2_7(my_ivn2_io_Stationary_matrix_2_7),
    .io_Stationary_matrix_3_0(my_ivn2_io_Stationary_matrix_3_0),
    .io_Stationary_matrix_3_1(my_ivn2_io_Stationary_matrix_3_1),
    .io_Stationary_matrix_3_2(my_ivn2_io_Stationary_matrix_3_2),
    .io_Stationary_matrix_3_3(my_ivn2_io_Stationary_matrix_3_3),
    .io_Stationary_matrix_3_4(my_ivn2_io_Stationary_matrix_3_4),
    .io_Stationary_matrix_3_5(my_ivn2_io_Stationary_matrix_3_5),
    .io_Stationary_matrix_3_6(my_ivn2_io_Stationary_matrix_3_6),
    .io_Stationary_matrix_3_7(my_ivn2_io_Stationary_matrix_3_7),
    .io_Stationary_matrix_4_0(my_ivn2_io_Stationary_matrix_4_0),
    .io_Stationary_matrix_4_1(my_ivn2_io_Stationary_matrix_4_1),
    .io_Stationary_matrix_4_2(my_ivn2_io_Stationary_matrix_4_2),
    .io_Stationary_matrix_4_3(my_ivn2_io_Stationary_matrix_4_3),
    .io_Stationary_matrix_4_4(my_ivn2_io_Stationary_matrix_4_4),
    .io_Stationary_matrix_4_5(my_ivn2_io_Stationary_matrix_4_5),
    .io_Stationary_matrix_4_6(my_ivn2_io_Stationary_matrix_4_6),
    .io_Stationary_matrix_4_7(my_ivn2_io_Stationary_matrix_4_7),
    .io_Stationary_matrix_5_0(my_ivn2_io_Stationary_matrix_5_0),
    .io_Stationary_matrix_5_1(my_ivn2_io_Stationary_matrix_5_1),
    .io_Stationary_matrix_5_2(my_ivn2_io_Stationary_matrix_5_2),
    .io_Stationary_matrix_5_3(my_ivn2_io_Stationary_matrix_5_3),
    .io_Stationary_matrix_5_4(my_ivn2_io_Stationary_matrix_5_4),
    .io_Stationary_matrix_5_5(my_ivn2_io_Stationary_matrix_5_5),
    .io_Stationary_matrix_5_6(my_ivn2_io_Stationary_matrix_5_6),
    .io_Stationary_matrix_5_7(my_ivn2_io_Stationary_matrix_5_7),
    .io_Stationary_matrix_6_0(my_ivn2_io_Stationary_matrix_6_0),
    .io_Stationary_matrix_6_1(my_ivn2_io_Stationary_matrix_6_1),
    .io_Stationary_matrix_6_2(my_ivn2_io_Stationary_matrix_6_2),
    .io_Stationary_matrix_6_3(my_ivn2_io_Stationary_matrix_6_3),
    .io_Stationary_matrix_6_4(my_ivn2_io_Stationary_matrix_6_4),
    .io_Stationary_matrix_6_5(my_ivn2_io_Stationary_matrix_6_5),
    .io_Stationary_matrix_6_6(my_ivn2_io_Stationary_matrix_6_6),
    .io_Stationary_matrix_6_7(my_ivn2_io_Stationary_matrix_6_7),
    .io_Stationary_matrix_7_0(my_ivn2_io_Stationary_matrix_7_0),
    .io_Stationary_matrix_7_1(my_ivn2_io_Stationary_matrix_7_1),
    .io_Stationary_matrix_7_2(my_ivn2_io_Stationary_matrix_7_2),
    .io_Stationary_matrix_7_3(my_ivn2_io_Stationary_matrix_7_3),
    .io_Stationary_matrix_7_4(my_ivn2_io_Stationary_matrix_7_4),
    .io_Stationary_matrix_7_5(my_ivn2_io_Stationary_matrix_7_5),
    .io_Stationary_matrix_7_6(my_ivn2_io_Stationary_matrix_7_6),
    .io_Stationary_matrix_7_7(my_ivn2_io_Stationary_matrix_7_7),
    .io_o_vn_0(my_ivn2_io_o_vn_0),
    .io_o_vn_1(my_ivn2_io_o_vn_1),
    .io_o_vn_2(my_ivn2_io_o_vn_2),
    .io_o_vn_3(my_ivn2_io_o_vn_3),
    .io_o_vn2_0(my_ivn2_io_o_vn2_0),
    .io_o_vn2_1(my_ivn2_io_o_vn2_1),
    .io_o_vn2_2(my_ivn2_io_o_vn2_2),
    .io_o_vn2_3(my_ivn2_io_o_vn2_3)
  );
  ivncontrol4_2 my_ivn3 ( // @[ivntop.scala 47:25]
    .clock(my_ivn3_clock),
    .reset(my_ivn3_reset),
    .io_Stationary_matrix_0_0(my_ivn3_io_Stationary_matrix_0_0),
    .io_Stationary_matrix_0_1(my_ivn3_io_Stationary_matrix_0_1),
    .io_Stationary_matrix_0_2(my_ivn3_io_Stationary_matrix_0_2),
    .io_Stationary_matrix_0_3(my_ivn3_io_Stationary_matrix_0_3),
    .io_Stationary_matrix_0_4(my_ivn3_io_Stationary_matrix_0_4),
    .io_Stationary_matrix_0_5(my_ivn3_io_Stationary_matrix_0_5),
    .io_Stationary_matrix_0_6(my_ivn3_io_Stationary_matrix_0_6),
    .io_Stationary_matrix_0_7(my_ivn3_io_Stationary_matrix_0_7),
    .io_Stationary_matrix_1_0(my_ivn3_io_Stationary_matrix_1_0),
    .io_Stationary_matrix_1_1(my_ivn3_io_Stationary_matrix_1_1),
    .io_Stationary_matrix_1_2(my_ivn3_io_Stationary_matrix_1_2),
    .io_Stationary_matrix_1_3(my_ivn3_io_Stationary_matrix_1_3),
    .io_Stationary_matrix_1_4(my_ivn3_io_Stationary_matrix_1_4),
    .io_Stationary_matrix_1_5(my_ivn3_io_Stationary_matrix_1_5),
    .io_Stationary_matrix_1_6(my_ivn3_io_Stationary_matrix_1_6),
    .io_Stationary_matrix_1_7(my_ivn3_io_Stationary_matrix_1_7),
    .io_Stationary_matrix_2_0(my_ivn3_io_Stationary_matrix_2_0),
    .io_Stationary_matrix_2_1(my_ivn3_io_Stationary_matrix_2_1),
    .io_Stationary_matrix_2_2(my_ivn3_io_Stationary_matrix_2_2),
    .io_Stationary_matrix_2_3(my_ivn3_io_Stationary_matrix_2_3),
    .io_Stationary_matrix_2_4(my_ivn3_io_Stationary_matrix_2_4),
    .io_Stationary_matrix_2_5(my_ivn3_io_Stationary_matrix_2_5),
    .io_Stationary_matrix_2_6(my_ivn3_io_Stationary_matrix_2_6),
    .io_Stationary_matrix_2_7(my_ivn3_io_Stationary_matrix_2_7),
    .io_Stationary_matrix_3_0(my_ivn3_io_Stationary_matrix_3_0),
    .io_Stationary_matrix_3_1(my_ivn3_io_Stationary_matrix_3_1),
    .io_Stationary_matrix_3_2(my_ivn3_io_Stationary_matrix_3_2),
    .io_Stationary_matrix_3_3(my_ivn3_io_Stationary_matrix_3_3),
    .io_Stationary_matrix_3_4(my_ivn3_io_Stationary_matrix_3_4),
    .io_Stationary_matrix_3_5(my_ivn3_io_Stationary_matrix_3_5),
    .io_Stationary_matrix_3_6(my_ivn3_io_Stationary_matrix_3_6),
    .io_Stationary_matrix_3_7(my_ivn3_io_Stationary_matrix_3_7),
    .io_Stationary_matrix_4_0(my_ivn3_io_Stationary_matrix_4_0),
    .io_Stationary_matrix_4_1(my_ivn3_io_Stationary_matrix_4_1),
    .io_Stationary_matrix_4_2(my_ivn3_io_Stationary_matrix_4_2),
    .io_Stationary_matrix_4_3(my_ivn3_io_Stationary_matrix_4_3),
    .io_Stationary_matrix_4_4(my_ivn3_io_Stationary_matrix_4_4),
    .io_Stationary_matrix_4_5(my_ivn3_io_Stationary_matrix_4_5),
    .io_Stationary_matrix_4_6(my_ivn3_io_Stationary_matrix_4_6),
    .io_Stationary_matrix_4_7(my_ivn3_io_Stationary_matrix_4_7),
    .io_Stationary_matrix_5_0(my_ivn3_io_Stationary_matrix_5_0),
    .io_Stationary_matrix_5_1(my_ivn3_io_Stationary_matrix_5_1),
    .io_Stationary_matrix_5_2(my_ivn3_io_Stationary_matrix_5_2),
    .io_Stationary_matrix_5_3(my_ivn3_io_Stationary_matrix_5_3),
    .io_Stationary_matrix_5_4(my_ivn3_io_Stationary_matrix_5_4),
    .io_Stationary_matrix_5_5(my_ivn3_io_Stationary_matrix_5_5),
    .io_Stationary_matrix_5_6(my_ivn3_io_Stationary_matrix_5_6),
    .io_Stationary_matrix_5_7(my_ivn3_io_Stationary_matrix_5_7),
    .io_Stationary_matrix_6_0(my_ivn3_io_Stationary_matrix_6_0),
    .io_Stationary_matrix_6_1(my_ivn3_io_Stationary_matrix_6_1),
    .io_Stationary_matrix_6_2(my_ivn3_io_Stationary_matrix_6_2),
    .io_Stationary_matrix_6_3(my_ivn3_io_Stationary_matrix_6_3),
    .io_Stationary_matrix_6_4(my_ivn3_io_Stationary_matrix_6_4),
    .io_Stationary_matrix_6_5(my_ivn3_io_Stationary_matrix_6_5),
    .io_Stationary_matrix_6_6(my_ivn3_io_Stationary_matrix_6_6),
    .io_Stationary_matrix_6_7(my_ivn3_io_Stationary_matrix_6_7),
    .io_Stationary_matrix_7_0(my_ivn3_io_Stationary_matrix_7_0),
    .io_Stationary_matrix_7_1(my_ivn3_io_Stationary_matrix_7_1),
    .io_Stationary_matrix_7_2(my_ivn3_io_Stationary_matrix_7_2),
    .io_Stationary_matrix_7_3(my_ivn3_io_Stationary_matrix_7_3),
    .io_Stationary_matrix_7_4(my_ivn3_io_Stationary_matrix_7_4),
    .io_Stationary_matrix_7_5(my_ivn3_io_Stationary_matrix_7_5),
    .io_Stationary_matrix_7_6(my_ivn3_io_Stationary_matrix_7_6),
    .io_Stationary_matrix_7_7(my_ivn3_io_Stationary_matrix_7_7),
    .io_o_vn_0(my_ivn3_io_o_vn_0),
    .io_o_vn_1(my_ivn3_io_o_vn_1),
    .io_o_vn_2(my_ivn3_io_o_vn_2),
    .io_o_vn_3(my_ivn3_io_o_vn_3),
    .io_o_vn2_0(my_ivn3_io_o_vn2_0),
    .io_o_vn2_1(my_ivn3_io_o_vn2_1),
    .io_o_vn2_2(my_ivn3_io_o_vn2_2),
    .io_o_vn2_3(my_ivn3_io_o_vn2_3)
  );
  ivncontrol4_3 my_ivn4 ( // @[ivntop.scala 54:25]
    .clock(my_ivn4_clock),
    .reset(my_ivn4_reset),
    .io_Stationary_matrix_0_0(my_ivn4_io_Stationary_matrix_0_0),
    .io_Stationary_matrix_0_1(my_ivn4_io_Stationary_matrix_0_1),
    .io_Stationary_matrix_0_2(my_ivn4_io_Stationary_matrix_0_2),
    .io_Stationary_matrix_0_3(my_ivn4_io_Stationary_matrix_0_3),
    .io_Stationary_matrix_0_4(my_ivn4_io_Stationary_matrix_0_4),
    .io_Stationary_matrix_0_5(my_ivn4_io_Stationary_matrix_0_5),
    .io_Stationary_matrix_0_6(my_ivn4_io_Stationary_matrix_0_6),
    .io_Stationary_matrix_0_7(my_ivn4_io_Stationary_matrix_0_7),
    .io_Stationary_matrix_1_0(my_ivn4_io_Stationary_matrix_1_0),
    .io_Stationary_matrix_1_1(my_ivn4_io_Stationary_matrix_1_1),
    .io_Stationary_matrix_1_2(my_ivn4_io_Stationary_matrix_1_2),
    .io_Stationary_matrix_1_3(my_ivn4_io_Stationary_matrix_1_3),
    .io_Stationary_matrix_1_4(my_ivn4_io_Stationary_matrix_1_4),
    .io_Stationary_matrix_1_5(my_ivn4_io_Stationary_matrix_1_5),
    .io_Stationary_matrix_1_6(my_ivn4_io_Stationary_matrix_1_6),
    .io_Stationary_matrix_1_7(my_ivn4_io_Stationary_matrix_1_7),
    .io_Stationary_matrix_2_0(my_ivn4_io_Stationary_matrix_2_0),
    .io_Stationary_matrix_2_1(my_ivn4_io_Stationary_matrix_2_1),
    .io_Stationary_matrix_2_2(my_ivn4_io_Stationary_matrix_2_2),
    .io_Stationary_matrix_2_3(my_ivn4_io_Stationary_matrix_2_3),
    .io_Stationary_matrix_2_4(my_ivn4_io_Stationary_matrix_2_4),
    .io_Stationary_matrix_2_5(my_ivn4_io_Stationary_matrix_2_5),
    .io_Stationary_matrix_2_6(my_ivn4_io_Stationary_matrix_2_6),
    .io_Stationary_matrix_2_7(my_ivn4_io_Stationary_matrix_2_7),
    .io_Stationary_matrix_3_0(my_ivn4_io_Stationary_matrix_3_0),
    .io_Stationary_matrix_3_1(my_ivn4_io_Stationary_matrix_3_1),
    .io_Stationary_matrix_3_2(my_ivn4_io_Stationary_matrix_3_2),
    .io_Stationary_matrix_3_3(my_ivn4_io_Stationary_matrix_3_3),
    .io_Stationary_matrix_3_4(my_ivn4_io_Stationary_matrix_3_4),
    .io_Stationary_matrix_3_5(my_ivn4_io_Stationary_matrix_3_5),
    .io_Stationary_matrix_3_6(my_ivn4_io_Stationary_matrix_3_6),
    .io_Stationary_matrix_3_7(my_ivn4_io_Stationary_matrix_3_7),
    .io_Stationary_matrix_4_0(my_ivn4_io_Stationary_matrix_4_0),
    .io_Stationary_matrix_4_1(my_ivn4_io_Stationary_matrix_4_1),
    .io_Stationary_matrix_4_2(my_ivn4_io_Stationary_matrix_4_2),
    .io_Stationary_matrix_4_3(my_ivn4_io_Stationary_matrix_4_3),
    .io_Stationary_matrix_4_4(my_ivn4_io_Stationary_matrix_4_4),
    .io_Stationary_matrix_4_5(my_ivn4_io_Stationary_matrix_4_5),
    .io_Stationary_matrix_4_6(my_ivn4_io_Stationary_matrix_4_6),
    .io_Stationary_matrix_4_7(my_ivn4_io_Stationary_matrix_4_7),
    .io_Stationary_matrix_5_0(my_ivn4_io_Stationary_matrix_5_0),
    .io_Stationary_matrix_5_1(my_ivn4_io_Stationary_matrix_5_1),
    .io_Stationary_matrix_5_2(my_ivn4_io_Stationary_matrix_5_2),
    .io_Stationary_matrix_5_3(my_ivn4_io_Stationary_matrix_5_3),
    .io_Stationary_matrix_5_4(my_ivn4_io_Stationary_matrix_5_4),
    .io_Stationary_matrix_5_5(my_ivn4_io_Stationary_matrix_5_5),
    .io_Stationary_matrix_5_6(my_ivn4_io_Stationary_matrix_5_6),
    .io_Stationary_matrix_5_7(my_ivn4_io_Stationary_matrix_5_7),
    .io_Stationary_matrix_6_0(my_ivn4_io_Stationary_matrix_6_0),
    .io_Stationary_matrix_6_1(my_ivn4_io_Stationary_matrix_6_1),
    .io_Stationary_matrix_6_2(my_ivn4_io_Stationary_matrix_6_2),
    .io_Stationary_matrix_6_3(my_ivn4_io_Stationary_matrix_6_3),
    .io_Stationary_matrix_6_4(my_ivn4_io_Stationary_matrix_6_4),
    .io_Stationary_matrix_6_5(my_ivn4_io_Stationary_matrix_6_5),
    .io_Stationary_matrix_6_6(my_ivn4_io_Stationary_matrix_6_6),
    .io_Stationary_matrix_6_7(my_ivn4_io_Stationary_matrix_6_7),
    .io_Stationary_matrix_7_0(my_ivn4_io_Stationary_matrix_7_0),
    .io_Stationary_matrix_7_1(my_ivn4_io_Stationary_matrix_7_1),
    .io_Stationary_matrix_7_2(my_ivn4_io_Stationary_matrix_7_2),
    .io_Stationary_matrix_7_3(my_ivn4_io_Stationary_matrix_7_3),
    .io_Stationary_matrix_7_4(my_ivn4_io_Stationary_matrix_7_4),
    .io_Stationary_matrix_7_5(my_ivn4_io_Stationary_matrix_7_5),
    .io_Stationary_matrix_7_6(my_ivn4_io_Stationary_matrix_7_6),
    .io_Stationary_matrix_7_7(my_ivn4_io_Stationary_matrix_7_7),
    .io_o_vn_0(my_ivn4_io_o_vn_0),
    .io_o_vn_1(my_ivn4_io_o_vn_1),
    .io_o_vn_2(my_ivn4_io_o_vn_2),
    .io_o_vn_3(my_ivn4_io_o_vn_3),
    .io_o_vn2_0(my_ivn4_io_o_vn2_0),
    .io_o_vn2_1(my_ivn4_io_o_vn2_1),
    .io_o_vn2_2(my_ivn4_io_o_vn2_2),
    .io_o_vn2_3(my_ivn4_io_o_vn2_3)
  );
  ivncontrol4_4 my_ivn5 ( // @[ivntop.scala 61:25]
    .clock(my_ivn5_clock),
    .reset(my_ivn5_reset),
    .io_Stationary_matrix_0_0(my_ivn5_io_Stationary_matrix_0_0),
    .io_Stationary_matrix_0_1(my_ivn5_io_Stationary_matrix_0_1),
    .io_Stationary_matrix_0_2(my_ivn5_io_Stationary_matrix_0_2),
    .io_Stationary_matrix_0_3(my_ivn5_io_Stationary_matrix_0_3),
    .io_Stationary_matrix_0_4(my_ivn5_io_Stationary_matrix_0_4),
    .io_Stationary_matrix_0_5(my_ivn5_io_Stationary_matrix_0_5),
    .io_Stationary_matrix_0_6(my_ivn5_io_Stationary_matrix_0_6),
    .io_Stationary_matrix_0_7(my_ivn5_io_Stationary_matrix_0_7),
    .io_Stationary_matrix_1_0(my_ivn5_io_Stationary_matrix_1_0),
    .io_Stationary_matrix_1_1(my_ivn5_io_Stationary_matrix_1_1),
    .io_Stationary_matrix_1_2(my_ivn5_io_Stationary_matrix_1_2),
    .io_Stationary_matrix_1_3(my_ivn5_io_Stationary_matrix_1_3),
    .io_Stationary_matrix_1_4(my_ivn5_io_Stationary_matrix_1_4),
    .io_Stationary_matrix_1_5(my_ivn5_io_Stationary_matrix_1_5),
    .io_Stationary_matrix_1_6(my_ivn5_io_Stationary_matrix_1_6),
    .io_Stationary_matrix_1_7(my_ivn5_io_Stationary_matrix_1_7),
    .io_Stationary_matrix_2_0(my_ivn5_io_Stationary_matrix_2_0),
    .io_Stationary_matrix_2_1(my_ivn5_io_Stationary_matrix_2_1),
    .io_Stationary_matrix_2_2(my_ivn5_io_Stationary_matrix_2_2),
    .io_Stationary_matrix_2_3(my_ivn5_io_Stationary_matrix_2_3),
    .io_Stationary_matrix_2_4(my_ivn5_io_Stationary_matrix_2_4),
    .io_Stationary_matrix_2_5(my_ivn5_io_Stationary_matrix_2_5),
    .io_Stationary_matrix_2_6(my_ivn5_io_Stationary_matrix_2_6),
    .io_Stationary_matrix_2_7(my_ivn5_io_Stationary_matrix_2_7),
    .io_Stationary_matrix_3_0(my_ivn5_io_Stationary_matrix_3_0),
    .io_Stationary_matrix_3_1(my_ivn5_io_Stationary_matrix_3_1),
    .io_Stationary_matrix_3_2(my_ivn5_io_Stationary_matrix_3_2),
    .io_Stationary_matrix_3_3(my_ivn5_io_Stationary_matrix_3_3),
    .io_Stationary_matrix_3_4(my_ivn5_io_Stationary_matrix_3_4),
    .io_Stationary_matrix_3_5(my_ivn5_io_Stationary_matrix_3_5),
    .io_Stationary_matrix_3_6(my_ivn5_io_Stationary_matrix_3_6),
    .io_Stationary_matrix_3_7(my_ivn5_io_Stationary_matrix_3_7),
    .io_Stationary_matrix_4_0(my_ivn5_io_Stationary_matrix_4_0),
    .io_Stationary_matrix_4_1(my_ivn5_io_Stationary_matrix_4_1),
    .io_Stationary_matrix_4_2(my_ivn5_io_Stationary_matrix_4_2),
    .io_Stationary_matrix_4_3(my_ivn5_io_Stationary_matrix_4_3),
    .io_Stationary_matrix_4_4(my_ivn5_io_Stationary_matrix_4_4),
    .io_Stationary_matrix_4_5(my_ivn5_io_Stationary_matrix_4_5),
    .io_Stationary_matrix_4_6(my_ivn5_io_Stationary_matrix_4_6),
    .io_Stationary_matrix_4_7(my_ivn5_io_Stationary_matrix_4_7),
    .io_Stationary_matrix_5_0(my_ivn5_io_Stationary_matrix_5_0),
    .io_Stationary_matrix_5_1(my_ivn5_io_Stationary_matrix_5_1),
    .io_Stationary_matrix_5_2(my_ivn5_io_Stationary_matrix_5_2),
    .io_Stationary_matrix_5_3(my_ivn5_io_Stationary_matrix_5_3),
    .io_Stationary_matrix_5_4(my_ivn5_io_Stationary_matrix_5_4),
    .io_Stationary_matrix_5_5(my_ivn5_io_Stationary_matrix_5_5),
    .io_Stationary_matrix_5_6(my_ivn5_io_Stationary_matrix_5_6),
    .io_Stationary_matrix_5_7(my_ivn5_io_Stationary_matrix_5_7),
    .io_Stationary_matrix_6_0(my_ivn5_io_Stationary_matrix_6_0),
    .io_Stationary_matrix_6_1(my_ivn5_io_Stationary_matrix_6_1),
    .io_Stationary_matrix_6_2(my_ivn5_io_Stationary_matrix_6_2),
    .io_Stationary_matrix_6_3(my_ivn5_io_Stationary_matrix_6_3),
    .io_Stationary_matrix_6_4(my_ivn5_io_Stationary_matrix_6_4),
    .io_Stationary_matrix_6_5(my_ivn5_io_Stationary_matrix_6_5),
    .io_Stationary_matrix_6_6(my_ivn5_io_Stationary_matrix_6_6),
    .io_Stationary_matrix_6_7(my_ivn5_io_Stationary_matrix_6_7),
    .io_Stationary_matrix_7_0(my_ivn5_io_Stationary_matrix_7_0),
    .io_Stationary_matrix_7_1(my_ivn5_io_Stationary_matrix_7_1),
    .io_Stationary_matrix_7_2(my_ivn5_io_Stationary_matrix_7_2),
    .io_Stationary_matrix_7_3(my_ivn5_io_Stationary_matrix_7_3),
    .io_Stationary_matrix_7_4(my_ivn5_io_Stationary_matrix_7_4),
    .io_Stationary_matrix_7_5(my_ivn5_io_Stationary_matrix_7_5),
    .io_Stationary_matrix_7_6(my_ivn5_io_Stationary_matrix_7_6),
    .io_Stationary_matrix_7_7(my_ivn5_io_Stationary_matrix_7_7),
    .io_o_vn_0(my_ivn5_io_o_vn_0),
    .io_o_vn_1(my_ivn5_io_o_vn_1),
    .io_o_vn_2(my_ivn5_io_o_vn_2),
    .io_o_vn_3(my_ivn5_io_o_vn_3),
    .io_o_vn2_0(my_ivn5_io_o_vn2_0),
    .io_o_vn2_1(my_ivn5_io_o_vn2_1),
    .io_o_vn2_2(my_ivn5_io_o_vn2_2),
    .io_o_vn2_3(my_ivn5_io_o_vn2_3)
  );
  ivncontrol4_5 my_ivn6 ( // @[ivntop.scala 68:25]
    .clock(my_ivn6_clock),
    .reset(my_ivn6_reset),
    .io_Stationary_matrix_0_0(my_ivn6_io_Stationary_matrix_0_0),
    .io_Stationary_matrix_0_1(my_ivn6_io_Stationary_matrix_0_1),
    .io_Stationary_matrix_0_2(my_ivn6_io_Stationary_matrix_0_2),
    .io_Stationary_matrix_0_3(my_ivn6_io_Stationary_matrix_0_3),
    .io_Stationary_matrix_0_4(my_ivn6_io_Stationary_matrix_0_4),
    .io_Stationary_matrix_0_5(my_ivn6_io_Stationary_matrix_0_5),
    .io_Stationary_matrix_0_6(my_ivn6_io_Stationary_matrix_0_6),
    .io_Stationary_matrix_0_7(my_ivn6_io_Stationary_matrix_0_7),
    .io_Stationary_matrix_1_0(my_ivn6_io_Stationary_matrix_1_0),
    .io_Stationary_matrix_1_1(my_ivn6_io_Stationary_matrix_1_1),
    .io_Stationary_matrix_1_2(my_ivn6_io_Stationary_matrix_1_2),
    .io_Stationary_matrix_1_3(my_ivn6_io_Stationary_matrix_1_3),
    .io_Stationary_matrix_1_4(my_ivn6_io_Stationary_matrix_1_4),
    .io_Stationary_matrix_1_5(my_ivn6_io_Stationary_matrix_1_5),
    .io_Stationary_matrix_1_6(my_ivn6_io_Stationary_matrix_1_6),
    .io_Stationary_matrix_1_7(my_ivn6_io_Stationary_matrix_1_7),
    .io_Stationary_matrix_2_0(my_ivn6_io_Stationary_matrix_2_0),
    .io_Stationary_matrix_2_1(my_ivn6_io_Stationary_matrix_2_1),
    .io_Stationary_matrix_2_2(my_ivn6_io_Stationary_matrix_2_2),
    .io_Stationary_matrix_2_3(my_ivn6_io_Stationary_matrix_2_3),
    .io_Stationary_matrix_2_4(my_ivn6_io_Stationary_matrix_2_4),
    .io_Stationary_matrix_2_5(my_ivn6_io_Stationary_matrix_2_5),
    .io_Stationary_matrix_2_6(my_ivn6_io_Stationary_matrix_2_6),
    .io_Stationary_matrix_2_7(my_ivn6_io_Stationary_matrix_2_7),
    .io_Stationary_matrix_3_0(my_ivn6_io_Stationary_matrix_3_0),
    .io_Stationary_matrix_3_1(my_ivn6_io_Stationary_matrix_3_1),
    .io_Stationary_matrix_3_2(my_ivn6_io_Stationary_matrix_3_2),
    .io_Stationary_matrix_3_3(my_ivn6_io_Stationary_matrix_3_3),
    .io_Stationary_matrix_3_4(my_ivn6_io_Stationary_matrix_3_4),
    .io_Stationary_matrix_3_5(my_ivn6_io_Stationary_matrix_3_5),
    .io_Stationary_matrix_3_6(my_ivn6_io_Stationary_matrix_3_6),
    .io_Stationary_matrix_3_7(my_ivn6_io_Stationary_matrix_3_7),
    .io_Stationary_matrix_4_0(my_ivn6_io_Stationary_matrix_4_0),
    .io_Stationary_matrix_4_1(my_ivn6_io_Stationary_matrix_4_1),
    .io_Stationary_matrix_4_2(my_ivn6_io_Stationary_matrix_4_2),
    .io_Stationary_matrix_4_3(my_ivn6_io_Stationary_matrix_4_3),
    .io_Stationary_matrix_4_4(my_ivn6_io_Stationary_matrix_4_4),
    .io_Stationary_matrix_4_5(my_ivn6_io_Stationary_matrix_4_5),
    .io_Stationary_matrix_4_6(my_ivn6_io_Stationary_matrix_4_6),
    .io_Stationary_matrix_4_7(my_ivn6_io_Stationary_matrix_4_7),
    .io_Stationary_matrix_5_0(my_ivn6_io_Stationary_matrix_5_0),
    .io_Stationary_matrix_5_1(my_ivn6_io_Stationary_matrix_5_1),
    .io_Stationary_matrix_5_2(my_ivn6_io_Stationary_matrix_5_2),
    .io_Stationary_matrix_5_3(my_ivn6_io_Stationary_matrix_5_3),
    .io_Stationary_matrix_5_4(my_ivn6_io_Stationary_matrix_5_4),
    .io_Stationary_matrix_5_5(my_ivn6_io_Stationary_matrix_5_5),
    .io_Stationary_matrix_5_6(my_ivn6_io_Stationary_matrix_5_6),
    .io_Stationary_matrix_5_7(my_ivn6_io_Stationary_matrix_5_7),
    .io_Stationary_matrix_6_0(my_ivn6_io_Stationary_matrix_6_0),
    .io_Stationary_matrix_6_1(my_ivn6_io_Stationary_matrix_6_1),
    .io_Stationary_matrix_6_2(my_ivn6_io_Stationary_matrix_6_2),
    .io_Stationary_matrix_6_3(my_ivn6_io_Stationary_matrix_6_3),
    .io_Stationary_matrix_6_4(my_ivn6_io_Stationary_matrix_6_4),
    .io_Stationary_matrix_6_5(my_ivn6_io_Stationary_matrix_6_5),
    .io_Stationary_matrix_6_6(my_ivn6_io_Stationary_matrix_6_6),
    .io_Stationary_matrix_6_7(my_ivn6_io_Stationary_matrix_6_7),
    .io_Stationary_matrix_7_0(my_ivn6_io_Stationary_matrix_7_0),
    .io_Stationary_matrix_7_1(my_ivn6_io_Stationary_matrix_7_1),
    .io_Stationary_matrix_7_2(my_ivn6_io_Stationary_matrix_7_2),
    .io_Stationary_matrix_7_3(my_ivn6_io_Stationary_matrix_7_3),
    .io_Stationary_matrix_7_4(my_ivn6_io_Stationary_matrix_7_4),
    .io_Stationary_matrix_7_5(my_ivn6_io_Stationary_matrix_7_5),
    .io_Stationary_matrix_7_6(my_ivn6_io_Stationary_matrix_7_6),
    .io_Stationary_matrix_7_7(my_ivn6_io_Stationary_matrix_7_7),
    .io_o_vn_0(my_ivn6_io_o_vn_0),
    .io_o_vn_1(my_ivn6_io_o_vn_1),
    .io_o_vn_2(my_ivn6_io_o_vn_2),
    .io_o_vn_3(my_ivn6_io_o_vn_3),
    .io_o_vn2_0(my_ivn6_io_o_vn2_0),
    .io_o_vn2_1(my_ivn6_io_o_vn2_1),
    .io_o_vn2_2(my_ivn6_io_o_vn2_2),
    .io_o_vn2_3(my_ivn6_io_o_vn2_3)
  );
  ivncontrol4_6 my_ivn7 ( // @[ivntop.scala 75:25]
    .clock(my_ivn7_clock),
    .reset(my_ivn7_reset),
    .io_Stationary_matrix_0_0(my_ivn7_io_Stationary_matrix_0_0),
    .io_Stationary_matrix_0_1(my_ivn7_io_Stationary_matrix_0_1),
    .io_Stationary_matrix_0_2(my_ivn7_io_Stationary_matrix_0_2),
    .io_Stationary_matrix_0_3(my_ivn7_io_Stationary_matrix_0_3),
    .io_Stationary_matrix_0_4(my_ivn7_io_Stationary_matrix_0_4),
    .io_Stationary_matrix_0_5(my_ivn7_io_Stationary_matrix_0_5),
    .io_Stationary_matrix_0_6(my_ivn7_io_Stationary_matrix_0_6),
    .io_Stationary_matrix_0_7(my_ivn7_io_Stationary_matrix_0_7),
    .io_Stationary_matrix_1_0(my_ivn7_io_Stationary_matrix_1_0),
    .io_Stationary_matrix_1_1(my_ivn7_io_Stationary_matrix_1_1),
    .io_Stationary_matrix_1_2(my_ivn7_io_Stationary_matrix_1_2),
    .io_Stationary_matrix_1_3(my_ivn7_io_Stationary_matrix_1_3),
    .io_Stationary_matrix_1_4(my_ivn7_io_Stationary_matrix_1_4),
    .io_Stationary_matrix_1_5(my_ivn7_io_Stationary_matrix_1_5),
    .io_Stationary_matrix_1_6(my_ivn7_io_Stationary_matrix_1_6),
    .io_Stationary_matrix_1_7(my_ivn7_io_Stationary_matrix_1_7),
    .io_Stationary_matrix_2_0(my_ivn7_io_Stationary_matrix_2_0),
    .io_Stationary_matrix_2_1(my_ivn7_io_Stationary_matrix_2_1),
    .io_Stationary_matrix_2_2(my_ivn7_io_Stationary_matrix_2_2),
    .io_Stationary_matrix_2_3(my_ivn7_io_Stationary_matrix_2_3),
    .io_Stationary_matrix_2_4(my_ivn7_io_Stationary_matrix_2_4),
    .io_Stationary_matrix_2_5(my_ivn7_io_Stationary_matrix_2_5),
    .io_Stationary_matrix_2_6(my_ivn7_io_Stationary_matrix_2_6),
    .io_Stationary_matrix_2_7(my_ivn7_io_Stationary_matrix_2_7),
    .io_Stationary_matrix_3_0(my_ivn7_io_Stationary_matrix_3_0),
    .io_Stationary_matrix_3_1(my_ivn7_io_Stationary_matrix_3_1),
    .io_Stationary_matrix_3_2(my_ivn7_io_Stationary_matrix_3_2),
    .io_Stationary_matrix_3_3(my_ivn7_io_Stationary_matrix_3_3),
    .io_Stationary_matrix_3_4(my_ivn7_io_Stationary_matrix_3_4),
    .io_Stationary_matrix_3_5(my_ivn7_io_Stationary_matrix_3_5),
    .io_Stationary_matrix_3_6(my_ivn7_io_Stationary_matrix_3_6),
    .io_Stationary_matrix_3_7(my_ivn7_io_Stationary_matrix_3_7),
    .io_Stationary_matrix_4_0(my_ivn7_io_Stationary_matrix_4_0),
    .io_Stationary_matrix_4_1(my_ivn7_io_Stationary_matrix_4_1),
    .io_Stationary_matrix_4_2(my_ivn7_io_Stationary_matrix_4_2),
    .io_Stationary_matrix_4_3(my_ivn7_io_Stationary_matrix_4_3),
    .io_Stationary_matrix_4_4(my_ivn7_io_Stationary_matrix_4_4),
    .io_Stationary_matrix_4_5(my_ivn7_io_Stationary_matrix_4_5),
    .io_Stationary_matrix_4_6(my_ivn7_io_Stationary_matrix_4_6),
    .io_Stationary_matrix_4_7(my_ivn7_io_Stationary_matrix_4_7),
    .io_Stationary_matrix_5_0(my_ivn7_io_Stationary_matrix_5_0),
    .io_Stationary_matrix_5_1(my_ivn7_io_Stationary_matrix_5_1),
    .io_Stationary_matrix_5_2(my_ivn7_io_Stationary_matrix_5_2),
    .io_Stationary_matrix_5_3(my_ivn7_io_Stationary_matrix_5_3),
    .io_Stationary_matrix_5_4(my_ivn7_io_Stationary_matrix_5_4),
    .io_Stationary_matrix_5_5(my_ivn7_io_Stationary_matrix_5_5),
    .io_Stationary_matrix_5_6(my_ivn7_io_Stationary_matrix_5_6),
    .io_Stationary_matrix_5_7(my_ivn7_io_Stationary_matrix_5_7),
    .io_Stationary_matrix_6_0(my_ivn7_io_Stationary_matrix_6_0),
    .io_Stationary_matrix_6_1(my_ivn7_io_Stationary_matrix_6_1),
    .io_Stationary_matrix_6_2(my_ivn7_io_Stationary_matrix_6_2),
    .io_Stationary_matrix_6_3(my_ivn7_io_Stationary_matrix_6_3),
    .io_Stationary_matrix_6_4(my_ivn7_io_Stationary_matrix_6_4),
    .io_Stationary_matrix_6_5(my_ivn7_io_Stationary_matrix_6_5),
    .io_Stationary_matrix_6_6(my_ivn7_io_Stationary_matrix_6_6),
    .io_Stationary_matrix_6_7(my_ivn7_io_Stationary_matrix_6_7),
    .io_Stationary_matrix_7_0(my_ivn7_io_Stationary_matrix_7_0),
    .io_Stationary_matrix_7_1(my_ivn7_io_Stationary_matrix_7_1),
    .io_Stationary_matrix_7_2(my_ivn7_io_Stationary_matrix_7_2),
    .io_Stationary_matrix_7_3(my_ivn7_io_Stationary_matrix_7_3),
    .io_Stationary_matrix_7_4(my_ivn7_io_Stationary_matrix_7_4),
    .io_Stationary_matrix_7_5(my_ivn7_io_Stationary_matrix_7_5),
    .io_Stationary_matrix_7_6(my_ivn7_io_Stationary_matrix_7_6),
    .io_Stationary_matrix_7_7(my_ivn7_io_Stationary_matrix_7_7),
    .io_o_vn_0(my_ivn7_io_o_vn_0),
    .io_o_vn_1(my_ivn7_io_o_vn_1),
    .io_o_vn_2(my_ivn7_io_o_vn_2),
    .io_o_vn_3(my_ivn7_io_o_vn_3),
    .io_o_vn2_0(my_ivn7_io_o_vn2_0),
    .io_o_vn2_1(my_ivn7_io_o_vn2_1),
    .io_o_vn2_2(my_ivn7_io_o_vn2_2),
    .io_o_vn2_3(my_ivn7_io_o_vn2_3)
  );
  ivncontrol4_7 my_ivn8 ( // @[ivntop.scala 82:25]
    .clock(my_ivn8_clock),
    .reset(my_ivn8_reset),
    .io_Stationary_matrix_0_0(my_ivn8_io_Stationary_matrix_0_0),
    .io_Stationary_matrix_0_1(my_ivn8_io_Stationary_matrix_0_1),
    .io_Stationary_matrix_0_2(my_ivn8_io_Stationary_matrix_0_2),
    .io_Stationary_matrix_0_3(my_ivn8_io_Stationary_matrix_0_3),
    .io_Stationary_matrix_0_4(my_ivn8_io_Stationary_matrix_0_4),
    .io_Stationary_matrix_0_5(my_ivn8_io_Stationary_matrix_0_5),
    .io_Stationary_matrix_0_6(my_ivn8_io_Stationary_matrix_0_6),
    .io_Stationary_matrix_0_7(my_ivn8_io_Stationary_matrix_0_7),
    .io_Stationary_matrix_1_0(my_ivn8_io_Stationary_matrix_1_0),
    .io_Stationary_matrix_1_1(my_ivn8_io_Stationary_matrix_1_1),
    .io_Stationary_matrix_1_2(my_ivn8_io_Stationary_matrix_1_2),
    .io_Stationary_matrix_1_3(my_ivn8_io_Stationary_matrix_1_3),
    .io_Stationary_matrix_1_4(my_ivn8_io_Stationary_matrix_1_4),
    .io_Stationary_matrix_1_5(my_ivn8_io_Stationary_matrix_1_5),
    .io_Stationary_matrix_1_6(my_ivn8_io_Stationary_matrix_1_6),
    .io_Stationary_matrix_1_7(my_ivn8_io_Stationary_matrix_1_7),
    .io_Stationary_matrix_2_0(my_ivn8_io_Stationary_matrix_2_0),
    .io_Stationary_matrix_2_1(my_ivn8_io_Stationary_matrix_2_1),
    .io_Stationary_matrix_2_2(my_ivn8_io_Stationary_matrix_2_2),
    .io_Stationary_matrix_2_3(my_ivn8_io_Stationary_matrix_2_3),
    .io_Stationary_matrix_2_4(my_ivn8_io_Stationary_matrix_2_4),
    .io_Stationary_matrix_2_5(my_ivn8_io_Stationary_matrix_2_5),
    .io_Stationary_matrix_2_6(my_ivn8_io_Stationary_matrix_2_6),
    .io_Stationary_matrix_2_7(my_ivn8_io_Stationary_matrix_2_7),
    .io_Stationary_matrix_3_0(my_ivn8_io_Stationary_matrix_3_0),
    .io_Stationary_matrix_3_1(my_ivn8_io_Stationary_matrix_3_1),
    .io_Stationary_matrix_3_2(my_ivn8_io_Stationary_matrix_3_2),
    .io_Stationary_matrix_3_3(my_ivn8_io_Stationary_matrix_3_3),
    .io_Stationary_matrix_3_4(my_ivn8_io_Stationary_matrix_3_4),
    .io_Stationary_matrix_3_5(my_ivn8_io_Stationary_matrix_3_5),
    .io_Stationary_matrix_3_6(my_ivn8_io_Stationary_matrix_3_6),
    .io_Stationary_matrix_3_7(my_ivn8_io_Stationary_matrix_3_7),
    .io_Stationary_matrix_4_0(my_ivn8_io_Stationary_matrix_4_0),
    .io_Stationary_matrix_4_1(my_ivn8_io_Stationary_matrix_4_1),
    .io_Stationary_matrix_4_2(my_ivn8_io_Stationary_matrix_4_2),
    .io_Stationary_matrix_4_3(my_ivn8_io_Stationary_matrix_4_3),
    .io_Stationary_matrix_4_4(my_ivn8_io_Stationary_matrix_4_4),
    .io_Stationary_matrix_4_5(my_ivn8_io_Stationary_matrix_4_5),
    .io_Stationary_matrix_4_6(my_ivn8_io_Stationary_matrix_4_6),
    .io_Stationary_matrix_4_7(my_ivn8_io_Stationary_matrix_4_7),
    .io_Stationary_matrix_5_0(my_ivn8_io_Stationary_matrix_5_0),
    .io_Stationary_matrix_5_1(my_ivn8_io_Stationary_matrix_5_1),
    .io_Stationary_matrix_5_2(my_ivn8_io_Stationary_matrix_5_2),
    .io_Stationary_matrix_5_3(my_ivn8_io_Stationary_matrix_5_3),
    .io_Stationary_matrix_5_4(my_ivn8_io_Stationary_matrix_5_4),
    .io_Stationary_matrix_5_5(my_ivn8_io_Stationary_matrix_5_5),
    .io_Stationary_matrix_5_6(my_ivn8_io_Stationary_matrix_5_6),
    .io_Stationary_matrix_5_7(my_ivn8_io_Stationary_matrix_5_7),
    .io_Stationary_matrix_6_0(my_ivn8_io_Stationary_matrix_6_0),
    .io_Stationary_matrix_6_1(my_ivn8_io_Stationary_matrix_6_1),
    .io_Stationary_matrix_6_2(my_ivn8_io_Stationary_matrix_6_2),
    .io_Stationary_matrix_6_3(my_ivn8_io_Stationary_matrix_6_3),
    .io_Stationary_matrix_6_4(my_ivn8_io_Stationary_matrix_6_4),
    .io_Stationary_matrix_6_5(my_ivn8_io_Stationary_matrix_6_5),
    .io_Stationary_matrix_6_6(my_ivn8_io_Stationary_matrix_6_6),
    .io_Stationary_matrix_6_7(my_ivn8_io_Stationary_matrix_6_7),
    .io_Stationary_matrix_7_0(my_ivn8_io_Stationary_matrix_7_0),
    .io_Stationary_matrix_7_1(my_ivn8_io_Stationary_matrix_7_1),
    .io_Stationary_matrix_7_2(my_ivn8_io_Stationary_matrix_7_2),
    .io_Stationary_matrix_7_3(my_ivn8_io_Stationary_matrix_7_3),
    .io_Stationary_matrix_7_4(my_ivn8_io_Stationary_matrix_7_4),
    .io_Stationary_matrix_7_5(my_ivn8_io_Stationary_matrix_7_5),
    .io_Stationary_matrix_7_6(my_ivn8_io_Stationary_matrix_7_6),
    .io_Stationary_matrix_7_7(my_ivn8_io_Stationary_matrix_7_7),
    .io_o_vn_0(my_ivn8_io_o_vn_0),
    .io_o_vn_1(my_ivn8_io_o_vn_1),
    .io_o_vn_2(my_ivn8_io_o_vn_2),
    .io_o_vn_3(my_ivn8_io_o_vn_3),
    .io_o_vn2_0(my_ivn8_io_o_vn2_0),
    .io_o_vn2_1(my_ivn8_io_o_vn2_1),
    .io_o_vn2_2(my_ivn8_io_o_vn2_2),
    .io_o_vn2_3(my_ivn8_io_o_vn2_3)
  );
  assign io_ProcessValid = my_ivn1_io_ProcessValid; // @[ivntop.scala 37:21]
  assign io_o_vn_0_0 = my_ivn1_io_o_vn_0; // @[ivntop.scala 95:16]
  assign io_o_vn_0_1 = my_ivn1_io_o_vn_1; // @[ivntop.scala 95:16]
  assign io_o_vn_0_2 = my_ivn1_io_o_vn_2; // @[ivntop.scala 95:16]
  assign io_o_vn_0_3 = my_ivn1_io_o_vn_3; // @[ivntop.scala 95:16]
  assign io_o_vn_1_0 = my_ivn1_io_o_vn2_0; // @[ivntop.scala 96:16]
  assign io_o_vn_1_1 = my_ivn1_io_o_vn2_1; // @[ivntop.scala 96:16]
  assign io_o_vn_1_2 = my_ivn1_io_o_vn2_2; // @[ivntop.scala 96:16]
  assign io_o_vn_1_3 = my_ivn1_io_o_vn2_3; // @[ivntop.scala 96:16]
  assign io_o_vn_2_0 = my_ivn2_io_o_vn_0; // @[ivntop.scala 97:16]
  assign io_o_vn_2_1 = my_ivn2_io_o_vn_1; // @[ivntop.scala 97:16]
  assign io_o_vn_2_2 = my_ivn2_io_o_vn_2; // @[ivntop.scala 97:16]
  assign io_o_vn_2_3 = my_ivn2_io_o_vn_3; // @[ivntop.scala 97:16]
  assign io_o_vn_3_0 = my_ivn2_io_o_vn2_0; // @[ivntop.scala 98:16]
  assign io_o_vn_3_1 = my_ivn2_io_o_vn2_1; // @[ivntop.scala 98:16]
  assign io_o_vn_3_2 = my_ivn2_io_o_vn2_2; // @[ivntop.scala 98:16]
  assign io_o_vn_3_3 = my_ivn2_io_o_vn2_3; // @[ivntop.scala 98:16]
  assign io_o_vn_4_0 = my_ivn3_io_o_vn_0; // @[ivntop.scala 99:16]
  assign io_o_vn_4_1 = my_ivn3_io_o_vn_1; // @[ivntop.scala 99:16]
  assign io_o_vn_4_2 = my_ivn3_io_o_vn_2; // @[ivntop.scala 99:16]
  assign io_o_vn_4_3 = my_ivn3_io_o_vn_3; // @[ivntop.scala 99:16]
  assign io_o_vn_5_0 = my_ivn3_io_o_vn2_0; // @[ivntop.scala 100:16]
  assign io_o_vn_5_1 = my_ivn3_io_o_vn2_1; // @[ivntop.scala 100:16]
  assign io_o_vn_5_2 = my_ivn3_io_o_vn2_2; // @[ivntop.scala 100:16]
  assign io_o_vn_5_3 = my_ivn3_io_o_vn2_3; // @[ivntop.scala 100:16]
  assign io_o_vn_6_0 = my_ivn4_io_o_vn_0; // @[ivntop.scala 101:16]
  assign io_o_vn_6_1 = my_ivn4_io_o_vn_1; // @[ivntop.scala 101:16]
  assign io_o_vn_6_2 = my_ivn4_io_o_vn_2; // @[ivntop.scala 101:16]
  assign io_o_vn_6_3 = my_ivn4_io_o_vn_3; // @[ivntop.scala 101:16]
  assign io_o_vn_7_0 = my_ivn4_io_o_vn2_0; // @[ivntop.scala 102:16]
  assign io_o_vn_7_1 = my_ivn4_io_o_vn2_1; // @[ivntop.scala 102:16]
  assign io_o_vn_7_2 = my_ivn4_io_o_vn2_2; // @[ivntop.scala 102:16]
  assign io_o_vn_7_3 = my_ivn4_io_o_vn2_3; // @[ivntop.scala 102:16]
  assign io_o_vn_8_0 = my_ivn5_io_o_vn_0; // @[ivntop.scala 103:16]
  assign io_o_vn_8_1 = my_ivn5_io_o_vn_1; // @[ivntop.scala 103:16]
  assign io_o_vn_8_2 = my_ivn5_io_o_vn_2; // @[ivntop.scala 103:16]
  assign io_o_vn_8_3 = my_ivn5_io_o_vn_3; // @[ivntop.scala 103:16]
  assign io_o_vn_9_0 = my_ivn5_io_o_vn2_0; // @[ivntop.scala 104:16]
  assign io_o_vn_9_1 = my_ivn5_io_o_vn2_1; // @[ivntop.scala 104:16]
  assign io_o_vn_9_2 = my_ivn5_io_o_vn2_2; // @[ivntop.scala 104:16]
  assign io_o_vn_9_3 = my_ivn5_io_o_vn2_3; // @[ivntop.scala 104:16]
  assign io_o_vn_10_0 = my_ivn6_io_o_vn_0; // @[ivntop.scala 105:17]
  assign io_o_vn_10_1 = my_ivn6_io_o_vn_1; // @[ivntop.scala 105:17]
  assign io_o_vn_10_2 = my_ivn6_io_o_vn_2; // @[ivntop.scala 105:17]
  assign io_o_vn_10_3 = my_ivn6_io_o_vn_3; // @[ivntop.scala 105:17]
  assign io_o_vn_11_0 = my_ivn6_io_o_vn2_0; // @[ivntop.scala 106:17]
  assign io_o_vn_11_1 = my_ivn6_io_o_vn2_1; // @[ivntop.scala 106:17]
  assign io_o_vn_11_2 = my_ivn6_io_o_vn2_2; // @[ivntop.scala 106:17]
  assign io_o_vn_11_3 = my_ivn6_io_o_vn2_3; // @[ivntop.scala 106:17]
  assign io_o_vn_12_0 = my_ivn7_io_o_vn_0; // @[ivntop.scala 107:17]
  assign io_o_vn_12_1 = my_ivn7_io_o_vn_1; // @[ivntop.scala 107:17]
  assign io_o_vn_12_2 = my_ivn7_io_o_vn_2; // @[ivntop.scala 107:17]
  assign io_o_vn_12_3 = my_ivn7_io_o_vn_3; // @[ivntop.scala 107:17]
  assign io_o_vn_13_0 = my_ivn7_io_o_vn2_0; // @[ivntop.scala 108:17]
  assign io_o_vn_13_1 = my_ivn7_io_o_vn2_1; // @[ivntop.scala 108:17]
  assign io_o_vn_13_2 = my_ivn7_io_o_vn2_2; // @[ivntop.scala 108:17]
  assign io_o_vn_13_3 = my_ivn7_io_o_vn2_3; // @[ivntop.scala 108:17]
  assign io_o_vn_14_0 = my_ivn8_io_o_vn_0; // @[ivntop.scala 109:17]
  assign io_o_vn_14_1 = my_ivn8_io_o_vn_1; // @[ivntop.scala 109:17]
  assign io_o_vn_14_2 = my_ivn8_io_o_vn_2; // @[ivntop.scala 109:17]
  assign io_o_vn_14_3 = my_ivn8_io_o_vn_3; // @[ivntop.scala 109:17]
  assign io_o_vn_15_0 = my_ivn8_io_o_vn2_0; // @[ivntop.scala 110:17]
  assign io_o_vn_15_1 = my_ivn8_io_o_vn2_1; // @[ivntop.scala 110:17]
  assign io_o_vn_15_2 = my_ivn8_io_o_vn2_2; // @[ivntop.scala 110:17]
  assign io_o_vn_15_3 = my_ivn8_io_o_vn2_3; // @[ivntop.scala 110:17]
  assign my_stationary_clock = clock;
  assign my_stationary_reset = reset;
  assign my_stationary_io_Stationary_matrix_0_0 = io_Stationary_matrix_0_0; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_0_1 = io_Stationary_matrix_0_1; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_0_2 = io_Stationary_matrix_0_2; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_0_3 = io_Stationary_matrix_0_3; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_0_4 = io_Stationary_matrix_0_4; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_0_5 = io_Stationary_matrix_0_5; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_0_6 = io_Stationary_matrix_0_6; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_0_7 = io_Stationary_matrix_0_7; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_1_0 = io_Stationary_matrix_1_0; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_1_1 = io_Stationary_matrix_1_1; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_1_2 = io_Stationary_matrix_1_2; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_1_3 = io_Stationary_matrix_1_3; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_1_4 = io_Stationary_matrix_1_4; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_1_5 = io_Stationary_matrix_1_5; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_1_6 = io_Stationary_matrix_1_6; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_1_7 = io_Stationary_matrix_1_7; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_2_0 = io_Stationary_matrix_2_0; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_2_1 = io_Stationary_matrix_2_1; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_2_2 = io_Stationary_matrix_2_2; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_2_3 = io_Stationary_matrix_2_3; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_2_4 = io_Stationary_matrix_2_4; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_2_5 = io_Stationary_matrix_2_5; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_2_6 = io_Stationary_matrix_2_6; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_2_7 = io_Stationary_matrix_2_7; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_3_0 = io_Stationary_matrix_3_0; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_3_1 = io_Stationary_matrix_3_1; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_3_2 = io_Stationary_matrix_3_2; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_3_3 = io_Stationary_matrix_3_3; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_3_4 = io_Stationary_matrix_3_4; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_3_5 = io_Stationary_matrix_3_5; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_3_6 = io_Stationary_matrix_3_6; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_3_7 = io_Stationary_matrix_3_7; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_4_0 = io_Stationary_matrix_4_0; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_4_1 = io_Stationary_matrix_4_1; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_4_2 = io_Stationary_matrix_4_2; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_4_3 = io_Stationary_matrix_4_3; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_4_4 = io_Stationary_matrix_4_4; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_4_5 = io_Stationary_matrix_4_5; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_4_6 = io_Stationary_matrix_4_6; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_4_7 = io_Stationary_matrix_4_7; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_5_0 = io_Stationary_matrix_5_0; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_5_1 = io_Stationary_matrix_5_1; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_5_2 = io_Stationary_matrix_5_2; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_5_3 = io_Stationary_matrix_5_3; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_5_4 = io_Stationary_matrix_5_4; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_5_5 = io_Stationary_matrix_5_5; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_5_6 = io_Stationary_matrix_5_6; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_5_7 = io_Stationary_matrix_5_7; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_6_0 = io_Stationary_matrix_6_0; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_6_1 = io_Stationary_matrix_6_1; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_6_2 = io_Stationary_matrix_6_2; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_6_3 = io_Stationary_matrix_6_3; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_6_4 = io_Stationary_matrix_6_4; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_6_5 = io_Stationary_matrix_6_5; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_6_6 = io_Stationary_matrix_6_6; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_6_7 = io_Stationary_matrix_6_7; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_7_0 = io_Stationary_matrix_7_0; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_7_1 = io_Stationary_matrix_7_1; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_7_2 = io_Stationary_matrix_7_2; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_7_3 = io_Stationary_matrix_7_3; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_7_4 = io_Stationary_matrix_7_4; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_7_5 = io_Stationary_matrix_7_5; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_7_6 = io_Stationary_matrix_7_6; // @[ivntop.scala 20:40]
  assign my_stationary_io_Stationary_matrix_7_7 = io_Stationary_matrix_7_7; // @[ivntop.scala 20:40]
  assign my_ivn1_clock = clock;
  assign my_ivn1_reset = reset;
  assign my_ivn1_io_Stationary_matrix_0_0 = my_stationary_io_o_Stationary_matrix1_0_0; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_0_1 = my_stationary_io_o_Stationary_matrix1_0_1; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_0_2 = my_stationary_io_o_Stationary_matrix1_0_2; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_0_3 = my_stationary_io_o_Stationary_matrix1_0_3; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_0_4 = my_stationary_io_o_Stationary_matrix1_0_4; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_0_5 = my_stationary_io_o_Stationary_matrix1_0_5; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_0_6 = my_stationary_io_o_Stationary_matrix1_0_6; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_0_7 = my_stationary_io_o_Stationary_matrix1_0_7; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_1_0 = my_stationary_io_o_Stationary_matrix1_1_0; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_1_1 = my_stationary_io_o_Stationary_matrix1_1_1; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_1_2 = my_stationary_io_o_Stationary_matrix1_1_2; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_1_3 = my_stationary_io_o_Stationary_matrix1_1_3; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_1_4 = my_stationary_io_o_Stationary_matrix1_1_4; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_1_5 = my_stationary_io_o_Stationary_matrix1_1_5; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_1_6 = my_stationary_io_o_Stationary_matrix1_1_6; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_1_7 = my_stationary_io_o_Stationary_matrix1_1_7; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_2_0 = my_stationary_io_o_Stationary_matrix1_2_0; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_2_1 = my_stationary_io_o_Stationary_matrix1_2_1; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_2_2 = my_stationary_io_o_Stationary_matrix1_2_2; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_2_3 = my_stationary_io_o_Stationary_matrix1_2_3; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_2_4 = my_stationary_io_o_Stationary_matrix1_2_4; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_2_5 = my_stationary_io_o_Stationary_matrix1_2_5; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_2_6 = my_stationary_io_o_Stationary_matrix1_2_6; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_2_7 = my_stationary_io_o_Stationary_matrix1_2_7; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_3_0 = my_stationary_io_o_Stationary_matrix1_3_0; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_3_1 = my_stationary_io_o_Stationary_matrix1_3_1; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_3_2 = my_stationary_io_o_Stationary_matrix1_3_2; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_3_3 = my_stationary_io_o_Stationary_matrix1_3_3; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_3_4 = my_stationary_io_o_Stationary_matrix1_3_4; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_3_5 = my_stationary_io_o_Stationary_matrix1_3_5; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_3_6 = my_stationary_io_o_Stationary_matrix1_3_6; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_3_7 = my_stationary_io_o_Stationary_matrix1_3_7; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_4_0 = my_stationary_io_o_Stationary_matrix1_4_0; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_4_1 = my_stationary_io_o_Stationary_matrix1_4_1; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_4_2 = my_stationary_io_o_Stationary_matrix1_4_2; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_4_3 = my_stationary_io_o_Stationary_matrix1_4_3; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_4_4 = my_stationary_io_o_Stationary_matrix1_4_4; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_4_5 = my_stationary_io_o_Stationary_matrix1_4_5; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_4_6 = my_stationary_io_o_Stationary_matrix1_4_6; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_4_7 = my_stationary_io_o_Stationary_matrix1_4_7; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_5_0 = my_stationary_io_o_Stationary_matrix1_5_0; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_5_1 = my_stationary_io_o_Stationary_matrix1_5_1; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_5_2 = my_stationary_io_o_Stationary_matrix1_5_2; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_5_3 = my_stationary_io_o_Stationary_matrix1_5_3; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_5_4 = my_stationary_io_o_Stationary_matrix1_5_4; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_5_5 = my_stationary_io_o_Stationary_matrix1_5_5; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_5_6 = my_stationary_io_o_Stationary_matrix1_5_6; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_5_7 = my_stationary_io_o_Stationary_matrix1_5_7; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_6_0 = my_stationary_io_o_Stationary_matrix1_6_0; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_6_1 = my_stationary_io_o_Stationary_matrix1_6_1; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_6_2 = my_stationary_io_o_Stationary_matrix1_6_2; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_6_3 = my_stationary_io_o_Stationary_matrix1_6_3; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_6_4 = my_stationary_io_o_Stationary_matrix1_6_4; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_6_5 = my_stationary_io_o_Stationary_matrix1_6_5; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_6_6 = my_stationary_io_o_Stationary_matrix1_6_6; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_6_7 = my_stationary_io_o_Stationary_matrix1_6_7; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_7_0 = my_stationary_io_o_Stationary_matrix1_7_0; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_7_1 = my_stationary_io_o_Stationary_matrix1_7_1; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_7_2 = my_stationary_io_o_Stationary_matrix1_7_2; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_7_3 = my_stationary_io_o_Stationary_matrix1_7_3; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_7_4 = my_stationary_io_o_Stationary_matrix1_7_4; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_7_5 = my_stationary_io_o_Stationary_matrix1_7_5; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_7_6 = my_stationary_io_o_Stationary_matrix1_7_6; // @[ivntop.scala 33:34]
  assign my_ivn1_io_Stationary_matrix_7_7 = my_stationary_io_o_Stationary_matrix1_7_7; // @[ivntop.scala 33:34]
  assign my_ivn2_clock = clock;
  assign my_ivn2_reset = reset;
  assign my_ivn2_io_Stationary_matrix_0_0 = my_stationary_io_o_Stationary_matrix2_0_0; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_0_1 = my_stationary_io_o_Stationary_matrix2_0_1; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_0_2 = my_stationary_io_o_Stationary_matrix2_0_2; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_0_3 = my_stationary_io_o_Stationary_matrix2_0_3; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_0_4 = my_stationary_io_o_Stationary_matrix2_0_4; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_0_5 = my_stationary_io_o_Stationary_matrix2_0_5; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_0_6 = my_stationary_io_o_Stationary_matrix2_0_6; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_0_7 = my_stationary_io_o_Stationary_matrix2_0_7; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_1_0 = my_stationary_io_o_Stationary_matrix2_1_0; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_1_1 = my_stationary_io_o_Stationary_matrix2_1_1; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_1_2 = my_stationary_io_o_Stationary_matrix2_1_2; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_1_3 = my_stationary_io_o_Stationary_matrix2_1_3; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_1_4 = my_stationary_io_o_Stationary_matrix2_1_4; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_1_5 = my_stationary_io_o_Stationary_matrix2_1_5; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_1_6 = my_stationary_io_o_Stationary_matrix2_1_6; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_1_7 = my_stationary_io_o_Stationary_matrix2_1_7; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_2_0 = my_stationary_io_o_Stationary_matrix2_2_0; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_2_1 = my_stationary_io_o_Stationary_matrix2_2_1; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_2_2 = my_stationary_io_o_Stationary_matrix2_2_2; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_2_3 = my_stationary_io_o_Stationary_matrix2_2_3; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_2_4 = my_stationary_io_o_Stationary_matrix2_2_4; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_2_5 = my_stationary_io_o_Stationary_matrix2_2_5; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_2_6 = my_stationary_io_o_Stationary_matrix2_2_6; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_2_7 = my_stationary_io_o_Stationary_matrix2_2_7; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_3_0 = my_stationary_io_o_Stationary_matrix2_3_0; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_3_1 = my_stationary_io_o_Stationary_matrix2_3_1; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_3_2 = my_stationary_io_o_Stationary_matrix2_3_2; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_3_3 = my_stationary_io_o_Stationary_matrix2_3_3; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_3_4 = my_stationary_io_o_Stationary_matrix2_3_4; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_3_5 = my_stationary_io_o_Stationary_matrix2_3_5; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_3_6 = my_stationary_io_o_Stationary_matrix2_3_6; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_3_7 = my_stationary_io_o_Stationary_matrix2_3_7; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_4_0 = my_stationary_io_o_Stationary_matrix2_4_0; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_4_1 = my_stationary_io_o_Stationary_matrix2_4_1; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_4_2 = my_stationary_io_o_Stationary_matrix2_4_2; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_4_3 = my_stationary_io_o_Stationary_matrix2_4_3; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_4_4 = my_stationary_io_o_Stationary_matrix2_4_4; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_4_5 = my_stationary_io_o_Stationary_matrix2_4_5; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_4_6 = my_stationary_io_o_Stationary_matrix2_4_6; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_4_7 = my_stationary_io_o_Stationary_matrix2_4_7; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_5_0 = my_stationary_io_o_Stationary_matrix2_5_0; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_5_1 = my_stationary_io_o_Stationary_matrix2_5_1; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_5_2 = my_stationary_io_o_Stationary_matrix2_5_2; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_5_3 = my_stationary_io_o_Stationary_matrix2_5_3; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_5_4 = my_stationary_io_o_Stationary_matrix2_5_4; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_5_5 = my_stationary_io_o_Stationary_matrix2_5_5; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_5_6 = my_stationary_io_o_Stationary_matrix2_5_6; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_5_7 = my_stationary_io_o_Stationary_matrix2_5_7; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_6_0 = my_stationary_io_o_Stationary_matrix2_6_0; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_6_1 = my_stationary_io_o_Stationary_matrix2_6_1; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_6_2 = my_stationary_io_o_Stationary_matrix2_6_2; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_6_3 = my_stationary_io_o_Stationary_matrix2_6_3; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_6_4 = my_stationary_io_o_Stationary_matrix2_6_4; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_6_5 = my_stationary_io_o_Stationary_matrix2_6_5; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_6_6 = my_stationary_io_o_Stationary_matrix2_6_6; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_6_7 = my_stationary_io_o_Stationary_matrix2_6_7; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_7_0 = my_stationary_io_o_Stationary_matrix2_7_0; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_7_1 = my_stationary_io_o_Stationary_matrix2_7_1; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_7_2 = my_stationary_io_o_Stationary_matrix2_7_2; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_7_3 = my_stationary_io_o_Stationary_matrix2_7_3; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_7_4 = my_stationary_io_o_Stationary_matrix2_7_4; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_7_5 = my_stationary_io_o_Stationary_matrix2_7_5; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_7_6 = my_stationary_io_o_Stationary_matrix2_7_6; // @[ivntop.scala 41:34]
  assign my_ivn2_io_Stationary_matrix_7_7 = my_stationary_io_o_Stationary_matrix2_7_7; // @[ivntop.scala 41:34]
  assign my_ivn3_clock = clock;
  assign my_ivn3_reset = reset;
  assign my_ivn3_io_Stationary_matrix_0_0 = my_stationary_io_o_Stationary_matrix3_0_0; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_0_1 = my_stationary_io_o_Stationary_matrix3_0_1; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_0_2 = my_stationary_io_o_Stationary_matrix3_0_2; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_0_3 = my_stationary_io_o_Stationary_matrix3_0_3; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_0_4 = my_stationary_io_o_Stationary_matrix3_0_4; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_0_5 = my_stationary_io_o_Stationary_matrix3_0_5; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_0_6 = my_stationary_io_o_Stationary_matrix3_0_6; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_0_7 = my_stationary_io_o_Stationary_matrix3_0_7; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_1_0 = my_stationary_io_o_Stationary_matrix3_1_0; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_1_1 = my_stationary_io_o_Stationary_matrix3_1_1; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_1_2 = my_stationary_io_o_Stationary_matrix3_1_2; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_1_3 = my_stationary_io_o_Stationary_matrix3_1_3; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_1_4 = my_stationary_io_o_Stationary_matrix3_1_4; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_1_5 = my_stationary_io_o_Stationary_matrix3_1_5; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_1_6 = my_stationary_io_o_Stationary_matrix3_1_6; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_1_7 = my_stationary_io_o_Stationary_matrix3_1_7; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_2_0 = my_stationary_io_o_Stationary_matrix3_2_0; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_2_1 = my_stationary_io_o_Stationary_matrix3_2_1; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_2_2 = my_stationary_io_o_Stationary_matrix3_2_2; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_2_3 = my_stationary_io_o_Stationary_matrix3_2_3; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_2_4 = my_stationary_io_o_Stationary_matrix3_2_4; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_2_5 = my_stationary_io_o_Stationary_matrix3_2_5; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_2_6 = my_stationary_io_o_Stationary_matrix3_2_6; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_2_7 = my_stationary_io_o_Stationary_matrix3_2_7; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_3_0 = my_stationary_io_o_Stationary_matrix3_3_0; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_3_1 = my_stationary_io_o_Stationary_matrix3_3_1; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_3_2 = my_stationary_io_o_Stationary_matrix3_3_2; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_3_3 = my_stationary_io_o_Stationary_matrix3_3_3; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_3_4 = my_stationary_io_o_Stationary_matrix3_3_4; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_3_5 = my_stationary_io_o_Stationary_matrix3_3_5; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_3_6 = my_stationary_io_o_Stationary_matrix3_3_6; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_3_7 = my_stationary_io_o_Stationary_matrix3_3_7; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_4_0 = my_stationary_io_o_Stationary_matrix3_4_0; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_4_1 = my_stationary_io_o_Stationary_matrix3_4_1; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_4_2 = my_stationary_io_o_Stationary_matrix3_4_2; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_4_3 = my_stationary_io_o_Stationary_matrix3_4_3; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_4_4 = my_stationary_io_o_Stationary_matrix3_4_4; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_4_5 = my_stationary_io_o_Stationary_matrix3_4_5; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_4_6 = my_stationary_io_o_Stationary_matrix3_4_6; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_4_7 = my_stationary_io_o_Stationary_matrix3_4_7; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_5_0 = my_stationary_io_o_Stationary_matrix3_5_0; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_5_1 = my_stationary_io_o_Stationary_matrix3_5_1; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_5_2 = my_stationary_io_o_Stationary_matrix3_5_2; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_5_3 = my_stationary_io_o_Stationary_matrix3_5_3; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_5_4 = my_stationary_io_o_Stationary_matrix3_5_4; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_5_5 = my_stationary_io_o_Stationary_matrix3_5_5; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_5_6 = my_stationary_io_o_Stationary_matrix3_5_6; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_5_7 = my_stationary_io_o_Stationary_matrix3_5_7; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_6_0 = my_stationary_io_o_Stationary_matrix3_6_0; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_6_1 = my_stationary_io_o_Stationary_matrix3_6_1; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_6_2 = my_stationary_io_o_Stationary_matrix3_6_2; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_6_3 = my_stationary_io_o_Stationary_matrix3_6_3; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_6_4 = my_stationary_io_o_Stationary_matrix3_6_4; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_6_5 = my_stationary_io_o_Stationary_matrix3_6_5; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_6_6 = my_stationary_io_o_Stationary_matrix3_6_6; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_6_7 = my_stationary_io_o_Stationary_matrix3_6_7; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_7_0 = my_stationary_io_o_Stationary_matrix3_7_0; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_7_1 = my_stationary_io_o_Stationary_matrix3_7_1; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_7_2 = my_stationary_io_o_Stationary_matrix3_7_2; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_7_3 = my_stationary_io_o_Stationary_matrix3_7_3; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_7_4 = my_stationary_io_o_Stationary_matrix3_7_4; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_7_5 = my_stationary_io_o_Stationary_matrix3_7_5; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_7_6 = my_stationary_io_o_Stationary_matrix3_7_6; // @[ivntop.scala 48:34]
  assign my_ivn3_io_Stationary_matrix_7_7 = my_stationary_io_o_Stationary_matrix3_7_7; // @[ivntop.scala 48:34]
  assign my_ivn4_clock = clock;
  assign my_ivn4_reset = reset;
  assign my_ivn4_io_Stationary_matrix_0_0 = my_stationary_io_o_Stationary_matrix4_0_0; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_0_1 = my_stationary_io_o_Stationary_matrix4_0_1; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_0_2 = my_stationary_io_o_Stationary_matrix4_0_2; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_0_3 = my_stationary_io_o_Stationary_matrix4_0_3; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_0_4 = my_stationary_io_o_Stationary_matrix4_0_4; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_0_5 = my_stationary_io_o_Stationary_matrix4_0_5; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_0_6 = my_stationary_io_o_Stationary_matrix4_0_6; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_0_7 = my_stationary_io_o_Stationary_matrix4_0_7; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_1_0 = my_stationary_io_o_Stationary_matrix4_1_0; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_1_1 = my_stationary_io_o_Stationary_matrix4_1_1; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_1_2 = my_stationary_io_o_Stationary_matrix4_1_2; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_1_3 = my_stationary_io_o_Stationary_matrix4_1_3; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_1_4 = my_stationary_io_o_Stationary_matrix4_1_4; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_1_5 = my_stationary_io_o_Stationary_matrix4_1_5; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_1_6 = my_stationary_io_o_Stationary_matrix4_1_6; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_1_7 = my_stationary_io_o_Stationary_matrix4_1_7; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_2_0 = my_stationary_io_o_Stationary_matrix4_2_0; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_2_1 = my_stationary_io_o_Stationary_matrix4_2_1; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_2_2 = my_stationary_io_o_Stationary_matrix4_2_2; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_2_3 = my_stationary_io_o_Stationary_matrix4_2_3; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_2_4 = my_stationary_io_o_Stationary_matrix4_2_4; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_2_5 = my_stationary_io_o_Stationary_matrix4_2_5; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_2_6 = my_stationary_io_o_Stationary_matrix4_2_6; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_2_7 = my_stationary_io_o_Stationary_matrix4_2_7; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_3_0 = my_stationary_io_o_Stationary_matrix4_3_0; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_3_1 = my_stationary_io_o_Stationary_matrix4_3_1; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_3_2 = my_stationary_io_o_Stationary_matrix4_3_2; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_3_3 = my_stationary_io_o_Stationary_matrix4_3_3; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_3_4 = my_stationary_io_o_Stationary_matrix4_3_4; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_3_5 = my_stationary_io_o_Stationary_matrix4_3_5; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_3_6 = my_stationary_io_o_Stationary_matrix4_3_6; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_3_7 = my_stationary_io_o_Stationary_matrix4_3_7; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_4_0 = my_stationary_io_o_Stationary_matrix4_4_0; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_4_1 = my_stationary_io_o_Stationary_matrix4_4_1; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_4_2 = my_stationary_io_o_Stationary_matrix4_4_2; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_4_3 = my_stationary_io_o_Stationary_matrix4_4_3; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_4_4 = my_stationary_io_o_Stationary_matrix4_4_4; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_4_5 = my_stationary_io_o_Stationary_matrix4_4_5; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_4_6 = my_stationary_io_o_Stationary_matrix4_4_6; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_4_7 = my_stationary_io_o_Stationary_matrix4_4_7; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_5_0 = my_stationary_io_o_Stationary_matrix4_5_0; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_5_1 = my_stationary_io_o_Stationary_matrix4_5_1; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_5_2 = my_stationary_io_o_Stationary_matrix4_5_2; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_5_3 = my_stationary_io_o_Stationary_matrix4_5_3; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_5_4 = my_stationary_io_o_Stationary_matrix4_5_4; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_5_5 = my_stationary_io_o_Stationary_matrix4_5_5; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_5_6 = my_stationary_io_o_Stationary_matrix4_5_6; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_5_7 = my_stationary_io_o_Stationary_matrix4_5_7; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_6_0 = my_stationary_io_o_Stationary_matrix4_6_0; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_6_1 = my_stationary_io_o_Stationary_matrix4_6_1; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_6_2 = my_stationary_io_o_Stationary_matrix4_6_2; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_6_3 = my_stationary_io_o_Stationary_matrix4_6_3; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_6_4 = my_stationary_io_o_Stationary_matrix4_6_4; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_6_5 = my_stationary_io_o_Stationary_matrix4_6_5; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_6_6 = my_stationary_io_o_Stationary_matrix4_6_6; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_6_7 = my_stationary_io_o_Stationary_matrix4_6_7; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_7_0 = my_stationary_io_o_Stationary_matrix4_7_0; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_7_1 = my_stationary_io_o_Stationary_matrix4_7_1; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_7_2 = my_stationary_io_o_Stationary_matrix4_7_2; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_7_3 = my_stationary_io_o_Stationary_matrix4_7_3; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_7_4 = my_stationary_io_o_Stationary_matrix4_7_4; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_7_5 = my_stationary_io_o_Stationary_matrix4_7_5; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_7_6 = my_stationary_io_o_Stationary_matrix4_7_6; // @[ivntop.scala 55:34]
  assign my_ivn4_io_Stationary_matrix_7_7 = my_stationary_io_o_Stationary_matrix4_7_7; // @[ivntop.scala 55:34]
  assign my_ivn5_clock = clock;
  assign my_ivn5_reset = reset;
  assign my_ivn5_io_Stationary_matrix_0_0 = my_stationary_io_o_Stationary_matrix5_0_0; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_0_1 = my_stationary_io_o_Stationary_matrix5_0_1; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_0_2 = my_stationary_io_o_Stationary_matrix5_0_2; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_0_3 = my_stationary_io_o_Stationary_matrix5_0_3; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_0_4 = my_stationary_io_o_Stationary_matrix5_0_4; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_0_5 = my_stationary_io_o_Stationary_matrix5_0_5; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_0_6 = my_stationary_io_o_Stationary_matrix5_0_6; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_0_7 = my_stationary_io_o_Stationary_matrix5_0_7; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_1_0 = my_stationary_io_o_Stationary_matrix5_1_0; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_1_1 = my_stationary_io_o_Stationary_matrix5_1_1; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_1_2 = my_stationary_io_o_Stationary_matrix5_1_2; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_1_3 = my_stationary_io_o_Stationary_matrix5_1_3; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_1_4 = my_stationary_io_o_Stationary_matrix5_1_4; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_1_5 = my_stationary_io_o_Stationary_matrix5_1_5; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_1_6 = my_stationary_io_o_Stationary_matrix5_1_6; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_1_7 = my_stationary_io_o_Stationary_matrix5_1_7; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_2_0 = my_stationary_io_o_Stationary_matrix5_2_0; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_2_1 = my_stationary_io_o_Stationary_matrix5_2_1; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_2_2 = my_stationary_io_o_Stationary_matrix5_2_2; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_2_3 = my_stationary_io_o_Stationary_matrix5_2_3; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_2_4 = my_stationary_io_o_Stationary_matrix5_2_4; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_2_5 = my_stationary_io_o_Stationary_matrix5_2_5; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_2_6 = my_stationary_io_o_Stationary_matrix5_2_6; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_2_7 = my_stationary_io_o_Stationary_matrix5_2_7; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_3_0 = my_stationary_io_o_Stationary_matrix5_3_0; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_3_1 = my_stationary_io_o_Stationary_matrix5_3_1; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_3_2 = my_stationary_io_o_Stationary_matrix5_3_2; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_3_3 = my_stationary_io_o_Stationary_matrix5_3_3; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_3_4 = my_stationary_io_o_Stationary_matrix5_3_4; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_3_5 = my_stationary_io_o_Stationary_matrix5_3_5; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_3_6 = my_stationary_io_o_Stationary_matrix5_3_6; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_3_7 = my_stationary_io_o_Stationary_matrix5_3_7; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_4_0 = my_stationary_io_o_Stationary_matrix5_4_0; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_4_1 = my_stationary_io_o_Stationary_matrix5_4_1; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_4_2 = my_stationary_io_o_Stationary_matrix5_4_2; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_4_3 = my_stationary_io_o_Stationary_matrix5_4_3; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_4_4 = my_stationary_io_o_Stationary_matrix5_4_4; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_4_5 = my_stationary_io_o_Stationary_matrix5_4_5; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_4_6 = my_stationary_io_o_Stationary_matrix5_4_6; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_4_7 = my_stationary_io_o_Stationary_matrix5_4_7; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_5_0 = my_stationary_io_o_Stationary_matrix5_5_0; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_5_1 = my_stationary_io_o_Stationary_matrix5_5_1; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_5_2 = my_stationary_io_o_Stationary_matrix5_5_2; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_5_3 = my_stationary_io_o_Stationary_matrix5_5_3; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_5_4 = my_stationary_io_o_Stationary_matrix5_5_4; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_5_5 = my_stationary_io_o_Stationary_matrix5_5_5; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_5_6 = my_stationary_io_o_Stationary_matrix5_5_6; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_5_7 = my_stationary_io_o_Stationary_matrix5_5_7; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_6_0 = my_stationary_io_o_Stationary_matrix5_6_0; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_6_1 = my_stationary_io_o_Stationary_matrix5_6_1; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_6_2 = my_stationary_io_o_Stationary_matrix5_6_2; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_6_3 = my_stationary_io_o_Stationary_matrix5_6_3; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_6_4 = my_stationary_io_o_Stationary_matrix5_6_4; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_6_5 = my_stationary_io_o_Stationary_matrix5_6_5; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_6_6 = my_stationary_io_o_Stationary_matrix5_6_6; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_6_7 = my_stationary_io_o_Stationary_matrix5_6_7; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_7_0 = my_stationary_io_o_Stationary_matrix5_7_0; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_7_1 = my_stationary_io_o_Stationary_matrix5_7_1; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_7_2 = my_stationary_io_o_Stationary_matrix5_7_2; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_7_3 = my_stationary_io_o_Stationary_matrix5_7_3; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_7_4 = my_stationary_io_o_Stationary_matrix5_7_4; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_7_5 = my_stationary_io_o_Stationary_matrix5_7_5; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_7_6 = my_stationary_io_o_Stationary_matrix5_7_6; // @[ivntop.scala 62:34]
  assign my_ivn5_io_Stationary_matrix_7_7 = my_stationary_io_o_Stationary_matrix5_7_7; // @[ivntop.scala 62:34]
  assign my_ivn6_clock = clock;
  assign my_ivn6_reset = reset;
  assign my_ivn6_io_Stationary_matrix_0_0 = my_stationary_io_o_Stationary_matrix6_0_0; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_0_1 = my_stationary_io_o_Stationary_matrix6_0_1; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_0_2 = my_stationary_io_o_Stationary_matrix6_0_2; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_0_3 = my_stationary_io_o_Stationary_matrix6_0_3; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_0_4 = my_stationary_io_o_Stationary_matrix6_0_4; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_0_5 = my_stationary_io_o_Stationary_matrix6_0_5; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_0_6 = my_stationary_io_o_Stationary_matrix6_0_6; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_0_7 = my_stationary_io_o_Stationary_matrix6_0_7; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_1_0 = my_stationary_io_o_Stationary_matrix6_1_0; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_1_1 = my_stationary_io_o_Stationary_matrix6_1_1; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_1_2 = my_stationary_io_o_Stationary_matrix6_1_2; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_1_3 = my_stationary_io_o_Stationary_matrix6_1_3; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_1_4 = my_stationary_io_o_Stationary_matrix6_1_4; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_1_5 = my_stationary_io_o_Stationary_matrix6_1_5; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_1_6 = my_stationary_io_o_Stationary_matrix6_1_6; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_1_7 = my_stationary_io_o_Stationary_matrix6_1_7; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_2_0 = my_stationary_io_o_Stationary_matrix6_2_0; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_2_1 = my_stationary_io_o_Stationary_matrix6_2_1; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_2_2 = my_stationary_io_o_Stationary_matrix6_2_2; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_2_3 = my_stationary_io_o_Stationary_matrix6_2_3; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_2_4 = my_stationary_io_o_Stationary_matrix6_2_4; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_2_5 = my_stationary_io_o_Stationary_matrix6_2_5; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_2_6 = my_stationary_io_o_Stationary_matrix6_2_6; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_2_7 = my_stationary_io_o_Stationary_matrix6_2_7; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_3_0 = my_stationary_io_o_Stationary_matrix6_3_0; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_3_1 = my_stationary_io_o_Stationary_matrix6_3_1; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_3_2 = my_stationary_io_o_Stationary_matrix6_3_2; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_3_3 = my_stationary_io_o_Stationary_matrix6_3_3; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_3_4 = my_stationary_io_o_Stationary_matrix6_3_4; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_3_5 = my_stationary_io_o_Stationary_matrix6_3_5; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_3_6 = my_stationary_io_o_Stationary_matrix6_3_6; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_3_7 = my_stationary_io_o_Stationary_matrix6_3_7; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_4_0 = my_stationary_io_o_Stationary_matrix6_4_0; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_4_1 = my_stationary_io_o_Stationary_matrix6_4_1; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_4_2 = my_stationary_io_o_Stationary_matrix6_4_2; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_4_3 = my_stationary_io_o_Stationary_matrix6_4_3; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_4_4 = my_stationary_io_o_Stationary_matrix6_4_4; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_4_5 = my_stationary_io_o_Stationary_matrix6_4_5; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_4_6 = my_stationary_io_o_Stationary_matrix6_4_6; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_4_7 = my_stationary_io_o_Stationary_matrix6_4_7; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_5_0 = my_stationary_io_o_Stationary_matrix6_5_0; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_5_1 = my_stationary_io_o_Stationary_matrix6_5_1; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_5_2 = my_stationary_io_o_Stationary_matrix6_5_2; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_5_3 = my_stationary_io_o_Stationary_matrix6_5_3; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_5_4 = my_stationary_io_o_Stationary_matrix6_5_4; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_5_5 = my_stationary_io_o_Stationary_matrix6_5_5; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_5_6 = my_stationary_io_o_Stationary_matrix6_5_6; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_5_7 = my_stationary_io_o_Stationary_matrix6_5_7; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_6_0 = my_stationary_io_o_Stationary_matrix6_6_0; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_6_1 = my_stationary_io_o_Stationary_matrix6_6_1; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_6_2 = my_stationary_io_o_Stationary_matrix6_6_2; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_6_3 = my_stationary_io_o_Stationary_matrix6_6_3; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_6_4 = my_stationary_io_o_Stationary_matrix6_6_4; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_6_5 = my_stationary_io_o_Stationary_matrix6_6_5; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_6_6 = my_stationary_io_o_Stationary_matrix6_6_6; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_6_7 = my_stationary_io_o_Stationary_matrix6_6_7; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_7_0 = my_stationary_io_o_Stationary_matrix6_7_0; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_7_1 = my_stationary_io_o_Stationary_matrix6_7_1; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_7_2 = my_stationary_io_o_Stationary_matrix6_7_2; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_7_3 = my_stationary_io_o_Stationary_matrix6_7_3; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_7_4 = my_stationary_io_o_Stationary_matrix6_7_4; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_7_5 = my_stationary_io_o_Stationary_matrix6_7_5; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_7_6 = my_stationary_io_o_Stationary_matrix6_7_6; // @[ivntop.scala 69:34]
  assign my_ivn6_io_Stationary_matrix_7_7 = my_stationary_io_o_Stationary_matrix6_7_7; // @[ivntop.scala 69:34]
  assign my_ivn7_clock = clock;
  assign my_ivn7_reset = reset;
  assign my_ivn7_io_Stationary_matrix_0_0 = my_stationary_io_o_Stationary_matrix7_0_0; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_0_1 = my_stationary_io_o_Stationary_matrix7_0_1; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_0_2 = my_stationary_io_o_Stationary_matrix7_0_2; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_0_3 = my_stationary_io_o_Stationary_matrix7_0_3; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_0_4 = my_stationary_io_o_Stationary_matrix7_0_4; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_0_5 = my_stationary_io_o_Stationary_matrix7_0_5; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_0_6 = my_stationary_io_o_Stationary_matrix7_0_6; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_0_7 = my_stationary_io_o_Stationary_matrix7_0_7; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_1_0 = my_stationary_io_o_Stationary_matrix7_1_0; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_1_1 = my_stationary_io_o_Stationary_matrix7_1_1; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_1_2 = my_stationary_io_o_Stationary_matrix7_1_2; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_1_3 = my_stationary_io_o_Stationary_matrix7_1_3; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_1_4 = my_stationary_io_o_Stationary_matrix7_1_4; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_1_5 = my_stationary_io_o_Stationary_matrix7_1_5; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_1_6 = my_stationary_io_o_Stationary_matrix7_1_6; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_1_7 = my_stationary_io_o_Stationary_matrix7_1_7; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_2_0 = my_stationary_io_o_Stationary_matrix7_2_0; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_2_1 = my_stationary_io_o_Stationary_matrix7_2_1; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_2_2 = my_stationary_io_o_Stationary_matrix7_2_2; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_2_3 = my_stationary_io_o_Stationary_matrix7_2_3; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_2_4 = my_stationary_io_o_Stationary_matrix7_2_4; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_2_5 = my_stationary_io_o_Stationary_matrix7_2_5; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_2_6 = my_stationary_io_o_Stationary_matrix7_2_6; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_2_7 = my_stationary_io_o_Stationary_matrix7_2_7; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_3_0 = my_stationary_io_o_Stationary_matrix7_3_0; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_3_1 = my_stationary_io_o_Stationary_matrix7_3_1; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_3_2 = my_stationary_io_o_Stationary_matrix7_3_2; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_3_3 = my_stationary_io_o_Stationary_matrix7_3_3; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_3_4 = my_stationary_io_o_Stationary_matrix7_3_4; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_3_5 = my_stationary_io_o_Stationary_matrix7_3_5; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_3_6 = my_stationary_io_o_Stationary_matrix7_3_6; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_3_7 = my_stationary_io_o_Stationary_matrix7_3_7; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_4_0 = my_stationary_io_o_Stationary_matrix7_4_0; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_4_1 = my_stationary_io_o_Stationary_matrix7_4_1; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_4_2 = my_stationary_io_o_Stationary_matrix7_4_2; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_4_3 = my_stationary_io_o_Stationary_matrix7_4_3; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_4_4 = my_stationary_io_o_Stationary_matrix7_4_4; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_4_5 = my_stationary_io_o_Stationary_matrix7_4_5; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_4_6 = my_stationary_io_o_Stationary_matrix7_4_6; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_4_7 = my_stationary_io_o_Stationary_matrix7_4_7; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_5_0 = my_stationary_io_o_Stationary_matrix7_5_0; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_5_1 = my_stationary_io_o_Stationary_matrix7_5_1; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_5_2 = my_stationary_io_o_Stationary_matrix7_5_2; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_5_3 = my_stationary_io_o_Stationary_matrix7_5_3; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_5_4 = my_stationary_io_o_Stationary_matrix7_5_4; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_5_5 = my_stationary_io_o_Stationary_matrix7_5_5; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_5_6 = my_stationary_io_o_Stationary_matrix7_5_6; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_5_7 = my_stationary_io_o_Stationary_matrix7_5_7; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_6_0 = my_stationary_io_o_Stationary_matrix7_6_0; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_6_1 = my_stationary_io_o_Stationary_matrix7_6_1; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_6_2 = my_stationary_io_o_Stationary_matrix7_6_2; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_6_3 = my_stationary_io_o_Stationary_matrix7_6_3; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_6_4 = my_stationary_io_o_Stationary_matrix7_6_4; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_6_5 = my_stationary_io_o_Stationary_matrix7_6_5; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_6_6 = my_stationary_io_o_Stationary_matrix7_6_6; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_6_7 = my_stationary_io_o_Stationary_matrix7_6_7; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_7_0 = my_stationary_io_o_Stationary_matrix7_7_0; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_7_1 = my_stationary_io_o_Stationary_matrix7_7_1; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_7_2 = my_stationary_io_o_Stationary_matrix7_7_2; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_7_3 = my_stationary_io_o_Stationary_matrix7_7_3; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_7_4 = my_stationary_io_o_Stationary_matrix7_7_4; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_7_5 = my_stationary_io_o_Stationary_matrix7_7_5; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_7_6 = my_stationary_io_o_Stationary_matrix7_7_6; // @[ivntop.scala 76:34]
  assign my_ivn7_io_Stationary_matrix_7_7 = my_stationary_io_o_Stationary_matrix7_7_7; // @[ivntop.scala 76:34]
  assign my_ivn8_clock = clock;
  assign my_ivn8_reset = reset;
  assign my_ivn8_io_Stationary_matrix_0_0 = my_stationary_io_o_Stationary_matrix8_0_0; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_0_1 = my_stationary_io_o_Stationary_matrix8_0_1; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_0_2 = my_stationary_io_o_Stationary_matrix8_0_2; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_0_3 = my_stationary_io_o_Stationary_matrix8_0_3; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_0_4 = my_stationary_io_o_Stationary_matrix8_0_4; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_0_5 = my_stationary_io_o_Stationary_matrix8_0_5; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_0_6 = my_stationary_io_o_Stationary_matrix8_0_6; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_0_7 = my_stationary_io_o_Stationary_matrix8_0_7; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_1_0 = my_stationary_io_o_Stationary_matrix8_1_0; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_1_1 = my_stationary_io_o_Stationary_matrix8_1_1; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_1_2 = my_stationary_io_o_Stationary_matrix8_1_2; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_1_3 = my_stationary_io_o_Stationary_matrix8_1_3; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_1_4 = my_stationary_io_o_Stationary_matrix8_1_4; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_1_5 = my_stationary_io_o_Stationary_matrix8_1_5; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_1_6 = my_stationary_io_o_Stationary_matrix8_1_6; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_1_7 = my_stationary_io_o_Stationary_matrix8_1_7; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_2_0 = my_stationary_io_o_Stationary_matrix8_2_0; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_2_1 = my_stationary_io_o_Stationary_matrix8_2_1; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_2_2 = my_stationary_io_o_Stationary_matrix8_2_2; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_2_3 = my_stationary_io_o_Stationary_matrix8_2_3; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_2_4 = my_stationary_io_o_Stationary_matrix8_2_4; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_2_5 = my_stationary_io_o_Stationary_matrix8_2_5; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_2_6 = my_stationary_io_o_Stationary_matrix8_2_6; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_2_7 = my_stationary_io_o_Stationary_matrix8_2_7; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_3_0 = my_stationary_io_o_Stationary_matrix8_3_0; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_3_1 = my_stationary_io_o_Stationary_matrix8_3_1; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_3_2 = my_stationary_io_o_Stationary_matrix8_3_2; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_3_3 = my_stationary_io_o_Stationary_matrix8_3_3; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_3_4 = my_stationary_io_o_Stationary_matrix8_3_4; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_3_5 = my_stationary_io_o_Stationary_matrix8_3_5; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_3_6 = my_stationary_io_o_Stationary_matrix8_3_6; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_3_7 = my_stationary_io_o_Stationary_matrix8_3_7; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_4_0 = my_stationary_io_o_Stationary_matrix8_4_0; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_4_1 = my_stationary_io_o_Stationary_matrix8_4_1; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_4_2 = my_stationary_io_o_Stationary_matrix8_4_2; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_4_3 = my_stationary_io_o_Stationary_matrix8_4_3; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_4_4 = my_stationary_io_o_Stationary_matrix8_4_4; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_4_5 = my_stationary_io_o_Stationary_matrix8_4_5; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_4_6 = my_stationary_io_o_Stationary_matrix8_4_6; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_4_7 = my_stationary_io_o_Stationary_matrix8_4_7; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_5_0 = my_stationary_io_o_Stationary_matrix8_5_0; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_5_1 = my_stationary_io_o_Stationary_matrix8_5_1; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_5_2 = my_stationary_io_o_Stationary_matrix8_5_2; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_5_3 = my_stationary_io_o_Stationary_matrix8_5_3; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_5_4 = my_stationary_io_o_Stationary_matrix8_5_4; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_5_5 = my_stationary_io_o_Stationary_matrix8_5_5; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_5_6 = my_stationary_io_o_Stationary_matrix8_5_6; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_5_7 = my_stationary_io_o_Stationary_matrix8_5_7; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_6_0 = my_stationary_io_o_Stationary_matrix8_6_0; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_6_1 = my_stationary_io_o_Stationary_matrix8_6_1; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_6_2 = my_stationary_io_o_Stationary_matrix8_6_2; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_6_3 = my_stationary_io_o_Stationary_matrix8_6_3; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_6_4 = my_stationary_io_o_Stationary_matrix8_6_4; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_6_5 = my_stationary_io_o_Stationary_matrix8_6_5; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_6_6 = my_stationary_io_o_Stationary_matrix8_6_6; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_6_7 = my_stationary_io_o_Stationary_matrix8_6_7; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_7_0 = my_stationary_io_o_Stationary_matrix8_7_0; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_7_1 = my_stationary_io_o_Stationary_matrix8_7_1; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_7_2 = my_stationary_io_o_Stationary_matrix8_7_2; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_7_3 = my_stationary_io_o_Stationary_matrix8_7_3; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_7_4 = my_stationary_io_o_Stationary_matrix8_7_4; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_7_5 = my_stationary_io_o_Stationary_matrix8_7_5; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_7_6 = my_stationary_io_o_Stationary_matrix8_7_6; // @[ivntop.scala 83:34]
  assign my_ivn8_io_Stationary_matrix_7_7 = my_stationary_io_o_Stationary_matrix8_7_7; // @[ivntop.scala 83:34]
endmodule
