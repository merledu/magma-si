module ReductionMux(
  input  [31:0] io_i_data_0,
  input  [31:0] io_i_data_1,
  output [31:0] io_o_data_0,
  output [31:0] io_o_data_1
);
  assign io_o_data_0 = io_i_data_0; // @[ReductionMux.scala 33:39 35:18 37:18]
  assign io_o_data_1 = io_i_data_1; // @[ReductionMux.scala 39:22]
endmodule
module SimpleAdder(
  input  [31:0] io_A,
  input  [31:0] io_B,
  output [31:0] io_O
);
  assign io_O = io_A + io_B; // @[SimpleAdder.scala 14:18]
endmodule
module EdgeAdderSwitch(
  input         clock,
  input         reset,
  input         io_i_valid,
  input  [63:0] io_i_data_bus_0,
  input  [63:0] io_i_data_bus_1,
  input  [2:0]  io_i_add_en,
  input  [4:0]  io_i_cmd,
  output [63:0] io_o_vn,
  output [1:0]  io_o_vn_valid,
  output [31:0] io_o_adder
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] reductionMux_io_i_data_0; // @[EdgeAdderSwitch.scala 23:28]
  wire [31:0] reductionMux_io_i_data_1; // @[EdgeAdderSwitch.scala 23:28]
  wire [31:0] reductionMux_io_o_data_0; // @[EdgeAdderSwitch.scala 23:28]
  wire [31:0] reductionMux_io_o_data_1; // @[EdgeAdderSwitch.scala 23:28]
  wire [31:0] adder32_io_A; // @[EdgeAdderSwitch.scala 27:23]
  wire [31:0] adder32_io_B; // @[EdgeAdderSwitch.scala 27:23]
  wire [31:0] adder32_io_O; // @[EdgeAdderSwitch.scala 27:23]
  reg  r_valid; // @[EdgeAdderSwitch.scala 31:24]
  reg [31:0] r_adder; // @[EdgeAdderSwitch.scala 32:24]
  reg [63:0] r_vn; // @[EdgeAdderSwitch.scala 33:21]
  reg [1:0] r_vn_valid; // @[EdgeAdderSwitch.scala 34:27]
  reg [2:0] r_add_en; // @[EdgeAdderSwitch.scala 35:25]
  wire [95:0] _r_vn_T = {io_i_data_bus_0,32'h0}; // @[Cat.scala 33:92]
  wire [95:0] _r_vn_T_1 = {32'h0,io_i_data_bus_1}; // @[Cat.scala 33:92]
  wire [63:0] _r_vn_T_2 = {reductionMux_io_o_data_0,reductionMux_io_o_data_1}; // @[Cat.scala 33:92]
  wire [1:0] _GEN_0 = 5'h0 == io_i_cmd ? 2'h0 : r_vn_valid; // @[EdgeAdderSwitch.scala 42:23 58:20 34:27]
  wire [63:0] _GEN_1 = 5'h5 == io_i_cmd ? _r_vn_T_2 : r_vn; // @[EdgeAdderSwitch.scala 42:23 54:14 33:21]
  wire [1:0] _GEN_2 = 5'h5 == io_i_cmd ? 2'h3 : _GEN_0; // @[EdgeAdderSwitch.scala 42:23 55:20]
  wire [31:0] _GEN_3 = 5'h4 == io_i_cmd ? reductionMux_io_o_data_0 : r_adder; // @[EdgeAdderSwitch.scala 42:23 49:17 32:24]
  wire [95:0] _GEN_4 = 5'h4 == io_i_cmd ? _r_vn_T_1 : {{32'd0}, _GEN_1}; // @[EdgeAdderSwitch.scala 42:23 50:14]
  wire [1:0] _GEN_5 = 5'h4 == io_i_cmd ? 2'h2 : _GEN_2; // @[EdgeAdderSwitch.scala 42:23 51:20]
  wire [95:0] _GEN_7 = 5'h3 == io_i_cmd ? _r_vn_T : _GEN_4; // @[EdgeAdderSwitch.scala 42:23 45:14]
  wire [95:0] _GEN_10 = r_valid ? _GEN_7 : {{32'd0}, r_vn}; // @[EdgeAdderSwitch.scala 33:21 41:25]
  wire [95:0] _GEN_13 = reset ? 96'h0 : _GEN_10; // @[EdgeAdderSwitch.scala 37:14 39:10]
  wire [31:0] _GEN_15 = r_add_en == 3'h0 ? r_adder : adder32_io_O; // @[EdgeAdderSwitch.scala 68:22 69:18 71:18]
  wire [95:0] _GEN_19 = reset ? 96'h0 : _GEN_13; // @[EdgeAdderSwitch.scala 33:{21,21}]
  ReductionMux reductionMux ( // @[EdgeAdderSwitch.scala 23:28]
    .io_i_data_0(reductionMux_io_i_data_0),
    .io_i_data_1(reductionMux_io_i_data_1),
    .io_o_data_0(reductionMux_io_o_data_0),
    .io_o_data_1(reductionMux_io_o_data_1)
  );
  SimpleAdder adder32 ( // @[EdgeAdderSwitch.scala 27:23]
    .io_A(adder32_io_A),
    .io_B(adder32_io_B),
    .io_O(adder32_io_O)
  );
  assign io_o_vn = reset ? 64'h0 : r_vn; // @[EdgeAdderSwitch.scala 63:14 65:13 73:13]
  assign io_o_vn_valid = reset ? 2'h0 : r_vn_valid; // @[EdgeAdderSwitch.scala 63:14 66:19 74:19]
  assign io_o_adder = reset ? 32'h0 : _GEN_15; // @[EdgeAdderSwitch.scala 63:14 64:16]
  assign reductionMux_io_i_data_0 = io_i_data_bus_0[31:0]; // @[EdgeAdderSwitch.scala 24:26]
  assign reductionMux_io_i_data_1 = io_i_data_bus_1[31:0]; // @[EdgeAdderSwitch.scala 24:26]
  assign adder32_io_A = reductionMux_io_o_data_1; // @[EdgeAdderSwitch.scala 28:16]
  assign adder32_io_B = reductionMux_io_o_data_0; // @[EdgeAdderSwitch.scala 29:16]
  always @(posedge clock) begin
    if (reset) begin // @[EdgeAdderSwitch.scala 31:24]
      r_valid <= 1'h0; // @[EdgeAdderSwitch.scala 31:24]
    end else begin
      r_valid <= io_i_valid; // @[EdgeAdderSwitch.scala 31:24]
    end
    if (reset) begin // @[EdgeAdderSwitch.scala 32:24]
      r_adder <= 32'h0; // @[EdgeAdderSwitch.scala 32:24]
    end else if (reset) begin // @[EdgeAdderSwitch.scala 37:14]
      r_adder <= 32'h0; // @[EdgeAdderSwitch.scala 38:13]
    end else if (r_valid) begin // @[EdgeAdderSwitch.scala 41:25]
      if (5'h3 == io_i_cmd) begin // @[EdgeAdderSwitch.scala 42:23]
        r_adder <= reductionMux_io_o_data_1; // @[EdgeAdderSwitch.scala 44:17]
      end else begin
        r_adder <= _GEN_3;
      end
    end
    r_vn <= _GEN_19[63:0]; // @[EdgeAdderSwitch.scala 33:{21,21}]
    if (reset) begin // @[EdgeAdderSwitch.scala 34:27]
      r_vn_valid <= 2'h0; // @[EdgeAdderSwitch.scala 34:27]
    end else if (reset) begin // @[EdgeAdderSwitch.scala 37:14]
      r_vn_valid <= 2'h0; // @[EdgeAdderSwitch.scala 40:16]
    end else if (r_valid) begin // @[EdgeAdderSwitch.scala 41:25]
      if (5'h3 == io_i_cmd) begin // @[EdgeAdderSwitch.scala 42:23]
        r_vn_valid <= 2'h1; // @[EdgeAdderSwitch.scala 46:20]
      end else begin
        r_vn_valid <= _GEN_5;
      end
    end
    if (reset) begin // @[EdgeAdderSwitch.scala 35:25]
      r_add_en <= 3'h0; // @[EdgeAdderSwitch.scala 35:25]
    end else begin
      r_add_en <= io_i_add_en; // @[EdgeAdderSwitch.scala 35:25]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  r_adder = _RAND_1[31:0];
  _RAND_2 = {2{`RANDOM}};
  r_vn = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  r_vn_valid = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  r_add_en = _RAND_4[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AdderSwitch(
  input         clock,
  input         reset,
  input         io_i_valid,
  input  [31:0] io_i_data_bus_0,
  input  [31:0] io_i_data_bus_1,
  input  [2:0]  io_i_add_en,
  input  [2:0]  io_i_cmd,
  output [1:0]  io_o_vn_valid,
  output [63:0] io_o_vn,
  output [31:0] io_o_adder_0,
  output [31:0] io_o_adder_1
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] reductionMux_io_i_data_0; // @[AdderSwitch.scala 25:28]
  wire [31:0] reductionMux_io_i_data_1; // @[AdderSwitch.scala 25:28]
  wire [31:0] reductionMux_io_o_data_0; // @[AdderSwitch.scala 25:28]
  wire [31:0] reductionMux_io_o_data_1; // @[AdderSwitch.scala 25:28]
  wire [31:0] adder32_io_A; // @[AdderSwitch.scala 29:23]
  wire [31:0] adder32_io_B; // @[AdderSwitch.scala 29:23]
  wire [31:0] adder32_io_O; // @[AdderSwitch.scala 29:23]
  reg [63:0] r_adder; // @[AdderSwitch.scala 33:24]
  reg [63:0] r_vn; // @[AdderSwitch.scala 34:21]
  reg [1:0] r_vn_valid; // @[AdderSwitch.scala 35:27]
  reg [2:0] r_add_en; // @[AdderSwitch.scala 36:25]
  wire [63:0] _r_adder_T = {reductionMux_io_o_data_0,reductionMux_io_o_data_1}; // @[Cat.scala 33:92]
  wire [62:0] _r_adder_T_1 = {31'h0,reductionMux_io_o_data_1}; // @[Cat.scala 33:92]
  wire [62:0] _r_adder_T_2 = {reductionMux_io_o_data_0,31'h0}; // @[Cat.scala 33:92]
  wire [1:0] _GEN_0 = 3'h0 == io_i_cmd ? 2'h0 : r_vn_valid; // @[AdderSwitch.scala 43:23 63:20 35:27]
  wire [63:0] _GEN_1 = 3'h5 == io_i_cmd ? _r_adder_T : r_vn; // @[AdderSwitch.scala 43:23 59:14 34:21]
  wire [1:0] _GEN_2 = 3'h5 == io_i_cmd ? 2'h3 : _GEN_0; // @[AdderSwitch.scala 43:23 60:20]
  wire [63:0] _GEN_3 = 3'h4 == io_i_cmd ? {{1'd0}, _r_adder_T_2} : r_adder; // @[AdderSwitch.scala 43:23 54:17 33:24]
  wire [63:0] _GEN_4 = 3'h4 == io_i_cmd ? {{32'd0}, io_i_data_bus_1} : _GEN_1; // @[AdderSwitch.scala 43:23 55:14]
  wire [1:0] _GEN_5 = 3'h4 == io_i_cmd ? 2'h2 : _GEN_2; // @[AdderSwitch.scala 43:23 56:20]
  wire [63:0] _GEN_6 = 3'h3 == io_i_cmd ? {{1'd0}, _r_adder_T_1} : _GEN_3; // @[AdderSwitch.scala 43:23 49:17]
  wire [63:0] _GEN_7 = 3'h3 == io_i_cmd ? {{32'd0}, io_i_data_bus_0} : _GEN_4; // @[AdderSwitch.scala 43:23 50:14]
  wire [1:0] _GEN_8 = 3'h3 == io_i_cmd ? 2'h1 : _GEN_5; // @[AdderSwitch.scala 43:23 51:20]
  wire [31:0] _WIRE_2_0 = adder32_io_O; // @[AdderSwitch.scala 76:{28,28}]
  wire [31:0] _GEN_18 = r_add_en == 3'h0 ? r_adder[31:0] : _WIRE_2_0; // @[AdderSwitch.scala 73:22 74:18 76:18]
  wire [31:0] _GEN_19 = r_add_en == 3'h0 ? r_adder[63:32] : _WIRE_2_0; // @[AdderSwitch.scala 73:22 74:18 76:18]
  ReductionMux reductionMux ( // @[AdderSwitch.scala 25:28]
    .io_i_data_0(reductionMux_io_i_data_0),
    .io_i_data_1(reductionMux_io_i_data_1),
    .io_o_data_0(reductionMux_io_o_data_0),
    .io_o_data_1(reductionMux_io_o_data_1)
  );
  SimpleAdder adder32 ( // @[AdderSwitch.scala 29:23]
    .io_A(adder32_io_A),
    .io_B(adder32_io_B),
    .io_O(adder32_io_O)
  );
  assign io_o_vn_valid = reset ? 2'h0 : r_vn_valid; // @[AdderSwitch.scala 68:14 71:19 79:19]
  assign io_o_vn = reset ? 64'h0 : r_vn; // @[AdderSwitch.scala 68:14 70:13 78:13]
  assign io_o_adder_0 = reset ? 32'h0 : _GEN_18; // @[AdderSwitch.scala 68:14 69:16]
  assign io_o_adder_1 = reset ? 32'h0 : _GEN_19; // @[AdderSwitch.scala 68:14 69:16]
  assign reductionMux_io_i_data_0 = io_i_data_bus_0; // @[AdderSwitch.scala 26:26]
  assign reductionMux_io_i_data_1 = io_i_data_bus_1; // @[AdderSwitch.scala 26:26]
  assign adder32_io_A = reductionMux_io_o_data_1; // @[AdderSwitch.scala 30:16]
  assign adder32_io_B = reductionMux_io_o_data_0; // @[AdderSwitch.scala 31:16]
  always @(posedge clock) begin
    if (reset) begin // @[AdderSwitch.scala 33:24]
      r_adder <= 64'h0; // @[AdderSwitch.scala 33:24]
    end else if (reset) begin // @[AdderSwitch.scala 38:14]
      r_adder <= 64'h0; // @[AdderSwitch.scala 39:13]
    end else if (io_i_valid) begin // @[AdderSwitch.scala 42:28]
      if (3'h1 == io_i_cmd) begin // @[AdderSwitch.scala 43:23]
        r_adder <= _r_adder_T; // @[AdderSwitch.scala 45:17]
      end else begin
        r_adder <= _GEN_6;
      end
    end
    if (reset) begin // @[AdderSwitch.scala 34:21]
      r_vn <= 64'h0; // @[AdderSwitch.scala 34:21]
    end else if (reset) begin // @[AdderSwitch.scala 38:14]
      r_vn <= 64'h0; // @[AdderSwitch.scala 40:10]
    end else if (io_i_valid) begin // @[AdderSwitch.scala 42:28]
      if (!(3'h1 == io_i_cmd)) begin // @[AdderSwitch.scala 43:23]
        r_vn <= _GEN_7;
      end
    end
    if (reset) begin // @[AdderSwitch.scala 35:27]
      r_vn_valid <= 2'h0; // @[AdderSwitch.scala 35:27]
    end else if (reset) begin // @[AdderSwitch.scala 38:14]
      r_vn_valid <= 2'h0; // @[AdderSwitch.scala 41:16]
    end else if (io_i_valid) begin // @[AdderSwitch.scala 42:28]
      if (3'h1 == io_i_cmd) begin // @[AdderSwitch.scala 43:23]
        r_vn_valid <= 2'h0; // @[AdderSwitch.scala 46:20]
      end else begin
        r_vn_valid <= _GEN_8;
      end
    end
    if (reset) begin // @[AdderSwitch.scala 36:25]
      r_add_en <= 3'h0; // @[AdderSwitch.scala 36:25]
    end else begin
      r_add_en <= io_i_add_en; // @[AdderSwitch.scala 36:25]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  r_adder = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  r_vn = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  r_vn_valid = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  r_add_en = _RAND_3[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ReductionMux_3(
  input  [31:0] io_i_data_0,
  input  [31:0] io_i_data_1,
  input  [31:0] io_i_data_2,
  input  [31:0] io_i_data_3,
  input  [1:0]  io_i_sel,
  output [31:0] io_o_data_0,
  output [31:0] io_o_data_1
);
  wire  w_sel_in_left = io_i_sel[0]; // @[ReductionMux.scala 29:32]
  wire  w_sel_in_right = io_i_sel[1]; // @[ReductionMux.scala 30:33]
  assign io_o_data_0 = w_sel_in_left ? io_i_data_1 : io_i_data_0; // @[ReductionMux.scala 35:{18,18}]
  assign io_o_data_1 = w_sel_in_right ? io_i_data_3 : io_i_data_2; // @[ReductionMux.scala 39:{22,22}]
endmodule
module EdgeAdderSwitch_2(
  input         clock,
  input         reset,
  input         io_i_valid,
  input  [63:0] io_i_data_bus_0,
  input  [63:0] io_i_data_bus_1,
  input  [63:0] io_i_data_bus_2,
  input  [63:0] io_i_data_bus_3,
  input  [2:0]  io_i_add_en,
  input  [4:0]  io_i_cmd,
  input  [1:0]  io_i_sel,
  output [63:0] io_o_vn,
  output [1:0]  io_o_vn_valid,
  output [31:0] io_o_adder
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] reductionMux_io_i_data_0; // @[EdgeAdderSwitch.scala 23:28]
  wire [31:0] reductionMux_io_i_data_1; // @[EdgeAdderSwitch.scala 23:28]
  wire [31:0] reductionMux_io_i_data_2; // @[EdgeAdderSwitch.scala 23:28]
  wire [31:0] reductionMux_io_i_data_3; // @[EdgeAdderSwitch.scala 23:28]
  wire [1:0] reductionMux_io_i_sel; // @[EdgeAdderSwitch.scala 23:28]
  wire [31:0] reductionMux_io_o_data_0; // @[EdgeAdderSwitch.scala 23:28]
  wire [31:0] reductionMux_io_o_data_1; // @[EdgeAdderSwitch.scala 23:28]
  wire [31:0] adder32_io_A; // @[EdgeAdderSwitch.scala 27:23]
  wire [31:0] adder32_io_B; // @[EdgeAdderSwitch.scala 27:23]
  wire [31:0] adder32_io_O; // @[EdgeAdderSwitch.scala 27:23]
  reg  r_valid; // @[EdgeAdderSwitch.scala 31:24]
  reg [31:0] r_adder; // @[EdgeAdderSwitch.scala 32:24]
  reg [63:0] r_vn; // @[EdgeAdderSwitch.scala 33:21]
  reg [1:0] r_vn_valid; // @[EdgeAdderSwitch.scala 34:27]
  reg [2:0] r_add_en; // @[EdgeAdderSwitch.scala 35:25]
  wire [95:0] _r_vn_T = {io_i_data_bus_0,32'h0}; // @[Cat.scala 33:92]
  wire [95:0] _r_vn_T_1 = {32'h0,io_i_data_bus_3}; // @[Cat.scala 33:92]
  wire [63:0] _r_vn_T_2 = {reductionMux_io_o_data_0,reductionMux_io_o_data_1}; // @[Cat.scala 33:92]
  wire [1:0] _GEN_0 = 5'h0 == io_i_cmd ? 2'h0 : r_vn_valid; // @[EdgeAdderSwitch.scala 42:23 58:20 34:27]
  wire [63:0] _GEN_1 = 5'h5 == io_i_cmd ? _r_vn_T_2 : r_vn; // @[EdgeAdderSwitch.scala 42:23 54:14 33:21]
  wire [1:0] _GEN_2 = 5'h5 == io_i_cmd ? 2'h3 : _GEN_0; // @[EdgeAdderSwitch.scala 42:23 55:20]
  wire [31:0] _GEN_3 = 5'h4 == io_i_cmd ? reductionMux_io_o_data_0 : r_adder; // @[EdgeAdderSwitch.scala 42:23 49:17 32:24]
  wire [95:0] _GEN_4 = 5'h4 == io_i_cmd ? _r_vn_T_1 : {{32'd0}, _GEN_1}; // @[EdgeAdderSwitch.scala 42:23 50:14]
  wire [1:0] _GEN_5 = 5'h4 == io_i_cmd ? 2'h2 : _GEN_2; // @[EdgeAdderSwitch.scala 42:23 51:20]
  wire [95:0] _GEN_7 = 5'h3 == io_i_cmd ? _r_vn_T : _GEN_4; // @[EdgeAdderSwitch.scala 42:23 45:14]
  wire [95:0] _GEN_10 = r_valid ? _GEN_7 : {{32'd0}, r_vn}; // @[EdgeAdderSwitch.scala 33:21 41:25]
  wire [95:0] _GEN_13 = reset ? 96'h0 : _GEN_10; // @[EdgeAdderSwitch.scala 37:14 39:10]
  wire [31:0] _GEN_15 = r_add_en == 3'h0 ? r_adder : adder32_io_O; // @[EdgeAdderSwitch.scala 68:22 69:18 71:18]
  wire [95:0] _GEN_19 = reset ? 96'h0 : _GEN_13; // @[EdgeAdderSwitch.scala 33:{21,21}]
  ReductionMux_3 reductionMux ( // @[EdgeAdderSwitch.scala 23:28]
    .io_i_data_0(reductionMux_io_i_data_0),
    .io_i_data_1(reductionMux_io_i_data_1),
    .io_i_data_2(reductionMux_io_i_data_2),
    .io_i_data_3(reductionMux_io_i_data_3),
    .io_i_sel(reductionMux_io_i_sel),
    .io_o_data_0(reductionMux_io_o_data_0),
    .io_o_data_1(reductionMux_io_o_data_1)
  );
  SimpleAdder adder32 ( // @[EdgeAdderSwitch.scala 27:23]
    .io_A(adder32_io_A),
    .io_B(adder32_io_B),
    .io_O(adder32_io_O)
  );
  assign io_o_vn = reset ? 64'h0 : r_vn; // @[EdgeAdderSwitch.scala 63:14 65:13 73:13]
  assign io_o_vn_valid = reset ? 2'h0 : r_vn_valid; // @[EdgeAdderSwitch.scala 63:14 66:19 74:19]
  assign io_o_adder = reset ? 32'h0 : _GEN_15; // @[EdgeAdderSwitch.scala 63:14 64:16]
  assign reductionMux_io_i_data_0 = io_i_data_bus_0[31:0]; // @[EdgeAdderSwitch.scala 24:26]
  assign reductionMux_io_i_data_1 = io_i_data_bus_1[31:0]; // @[EdgeAdderSwitch.scala 24:26]
  assign reductionMux_io_i_data_2 = io_i_data_bus_2[31:0]; // @[EdgeAdderSwitch.scala 24:26]
  assign reductionMux_io_i_data_3 = io_i_data_bus_3[31:0]; // @[EdgeAdderSwitch.scala 24:26]
  assign reductionMux_io_i_sel = io_i_sel; // @[EdgeAdderSwitch.scala 25:25]
  assign adder32_io_A = reductionMux_io_o_data_1; // @[EdgeAdderSwitch.scala 28:16]
  assign adder32_io_B = reductionMux_io_o_data_0; // @[EdgeAdderSwitch.scala 29:16]
  always @(posedge clock) begin
    if (reset) begin // @[EdgeAdderSwitch.scala 31:24]
      r_valid <= 1'h0; // @[EdgeAdderSwitch.scala 31:24]
    end else begin
      r_valid <= io_i_valid; // @[EdgeAdderSwitch.scala 31:24]
    end
    if (reset) begin // @[EdgeAdderSwitch.scala 32:24]
      r_adder <= 32'h0; // @[EdgeAdderSwitch.scala 32:24]
    end else if (reset) begin // @[EdgeAdderSwitch.scala 37:14]
      r_adder <= 32'h0; // @[EdgeAdderSwitch.scala 38:13]
    end else if (r_valid) begin // @[EdgeAdderSwitch.scala 41:25]
      if (5'h3 == io_i_cmd) begin // @[EdgeAdderSwitch.scala 42:23]
        r_adder <= reductionMux_io_o_data_1; // @[EdgeAdderSwitch.scala 44:17]
      end else begin
        r_adder <= _GEN_3;
      end
    end
    r_vn <= _GEN_19[63:0]; // @[EdgeAdderSwitch.scala 33:{21,21}]
    if (reset) begin // @[EdgeAdderSwitch.scala 34:27]
      r_vn_valid <= 2'h0; // @[EdgeAdderSwitch.scala 34:27]
    end else if (reset) begin // @[EdgeAdderSwitch.scala 37:14]
      r_vn_valid <= 2'h0; // @[EdgeAdderSwitch.scala 40:16]
    end else if (r_valid) begin // @[EdgeAdderSwitch.scala 41:25]
      if (5'h3 == io_i_cmd) begin // @[EdgeAdderSwitch.scala 42:23]
        r_vn_valid <= 2'h1; // @[EdgeAdderSwitch.scala 46:20]
      end else begin
        r_vn_valid <= _GEN_5;
      end
    end
    if (reset) begin // @[EdgeAdderSwitch.scala 35:25]
      r_add_en <= 3'h0; // @[EdgeAdderSwitch.scala 35:25]
    end else begin
      r_add_en <= io_i_add_en; // @[EdgeAdderSwitch.scala 35:25]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  r_adder = _RAND_1[31:0];
  _RAND_2 = {2{`RANDOM}};
  r_vn = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  r_vn_valid = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  r_add_en = _RAND_4[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ReductionMux_7(
  input  [31:0] io_i_data_0,
  input  [31:0] io_i_data_1,
  input  [31:0] io_i_data_2,
  input  [31:0] io_i_data_3,
  input  [31:0] io_i_data_4,
  input  [31:0] io_i_data_5,
  input  [3:0]  io_i_sel,
  output [31:0] io_o_data_0,
  output [31:0] io_o_data_1
);
  wire [1:0] w_sel_in_left = io_i_sel[1:0]; // @[ReductionMux.scala 29:32]
  wire [1:0] w_sel_in_right = io_i_sel[3:2]; // @[ReductionMux.scala 30:33]
  wire [31:0] _GEN_1 = 2'h1 == w_sel_in_left ? io_i_data_1 : io_i_data_0; // @[ReductionMux.scala 35:{18,18}]
  wire [31:0] _GEN_2 = 2'h2 == w_sel_in_left ? io_i_data_2 : _GEN_1; // @[ReductionMux.scala 35:{18,18}]
  wire [31:0] _GEN_5 = 2'h1 == w_sel_in_right ? io_i_data_4 : io_i_data_3; // @[ReductionMux.scala 39:{22,22}]
  wire [31:0] _GEN_6 = 2'h2 == w_sel_in_right ? io_i_data_5 : _GEN_5; // @[ReductionMux.scala 39:{22,22}]
  assign io_o_data_0 = w_sel_in_left < 2'h2 ? _GEN_2 : 32'h0; // @[ReductionMux.scala 33:39 35:18 37:18]
  assign io_o_data_1 = w_sel_in_right < 2'h3 ? _GEN_6 : 32'h0; // @[ReductionMux.scala 39:22]
endmodule
module EdgeAdderSwitch_3(
  input         clock,
  input         reset,
  input         io_i_valid,
  input  [63:0] io_i_data_bus_0,
  input  [63:0] io_i_data_bus_1,
  input  [63:0] io_i_data_bus_2,
  input  [63:0] io_i_data_bus_3,
  input  [63:0] io_i_data_bus_4,
  input  [63:0] io_i_data_bus_5,
  input  [2:0]  io_i_add_en,
  input  [4:0]  io_i_cmd,
  input  [3:0]  io_i_sel,
  output [63:0] io_o_vn,
  output [1:0]  io_o_vn_valid,
  output [31:0] io_o_adder
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] reductionMux_io_i_data_0; // @[EdgeAdderSwitch.scala 23:28]
  wire [31:0] reductionMux_io_i_data_1; // @[EdgeAdderSwitch.scala 23:28]
  wire [31:0] reductionMux_io_i_data_2; // @[EdgeAdderSwitch.scala 23:28]
  wire [31:0] reductionMux_io_i_data_3; // @[EdgeAdderSwitch.scala 23:28]
  wire [31:0] reductionMux_io_i_data_4; // @[EdgeAdderSwitch.scala 23:28]
  wire [31:0] reductionMux_io_i_data_5; // @[EdgeAdderSwitch.scala 23:28]
  wire [3:0] reductionMux_io_i_sel; // @[EdgeAdderSwitch.scala 23:28]
  wire [31:0] reductionMux_io_o_data_0; // @[EdgeAdderSwitch.scala 23:28]
  wire [31:0] reductionMux_io_o_data_1; // @[EdgeAdderSwitch.scala 23:28]
  wire [31:0] adder32_io_A; // @[EdgeAdderSwitch.scala 27:23]
  wire [31:0] adder32_io_B; // @[EdgeAdderSwitch.scala 27:23]
  wire [31:0] adder32_io_O; // @[EdgeAdderSwitch.scala 27:23]
  reg  r_valid; // @[EdgeAdderSwitch.scala 31:24]
  reg [31:0] r_adder; // @[EdgeAdderSwitch.scala 32:24]
  reg [63:0] r_vn; // @[EdgeAdderSwitch.scala 33:21]
  reg [1:0] r_vn_valid; // @[EdgeAdderSwitch.scala 34:27]
  reg [2:0] r_add_en; // @[EdgeAdderSwitch.scala 35:25]
  wire [95:0] _r_vn_T = {io_i_data_bus_0,32'h0}; // @[Cat.scala 33:92]
  wire [95:0] _r_vn_T_1 = {32'h0,io_i_data_bus_5}; // @[Cat.scala 33:92]
  wire [63:0] _r_vn_T_2 = {reductionMux_io_o_data_0,reductionMux_io_o_data_1}; // @[Cat.scala 33:92]
  wire [1:0] _GEN_0 = 5'h0 == io_i_cmd ? 2'h0 : r_vn_valid; // @[EdgeAdderSwitch.scala 42:23 58:20 34:27]
  wire [63:0] _GEN_1 = 5'h5 == io_i_cmd ? _r_vn_T_2 : r_vn; // @[EdgeAdderSwitch.scala 42:23 54:14 33:21]
  wire [1:0] _GEN_2 = 5'h5 == io_i_cmd ? 2'h3 : _GEN_0; // @[EdgeAdderSwitch.scala 42:23 55:20]
  wire [31:0] _GEN_3 = 5'h4 == io_i_cmd ? reductionMux_io_o_data_0 : r_adder; // @[EdgeAdderSwitch.scala 42:23 49:17 32:24]
  wire [95:0] _GEN_4 = 5'h4 == io_i_cmd ? _r_vn_T_1 : {{32'd0}, _GEN_1}; // @[EdgeAdderSwitch.scala 42:23 50:14]
  wire [1:0] _GEN_5 = 5'h4 == io_i_cmd ? 2'h2 : _GEN_2; // @[EdgeAdderSwitch.scala 42:23 51:20]
  wire [95:0] _GEN_7 = 5'h3 == io_i_cmd ? _r_vn_T : _GEN_4; // @[EdgeAdderSwitch.scala 42:23 45:14]
  wire [95:0] _GEN_10 = r_valid ? _GEN_7 : {{32'd0}, r_vn}; // @[EdgeAdderSwitch.scala 33:21 41:25]
  wire [95:0] _GEN_13 = reset ? 96'h0 : _GEN_10; // @[EdgeAdderSwitch.scala 37:14 39:10]
  wire [31:0] _GEN_15 = r_add_en == 3'h0 ? r_adder : adder32_io_O; // @[EdgeAdderSwitch.scala 68:22 69:18 71:18]
  wire [95:0] _GEN_19 = reset ? 96'h0 : _GEN_13; // @[EdgeAdderSwitch.scala 33:{21,21}]
  ReductionMux_7 reductionMux ( // @[EdgeAdderSwitch.scala 23:28]
    .io_i_data_0(reductionMux_io_i_data_0),
    .io_i_data_1(reductionMux_io_i_data_1),
    .io_i_data_2(reductionMux_io_i_data_2),
    .io_i_data_3(reductionMux_io_i_data_3),
    .io_i_data_4(reductionMux_io_i_data_4),
    .io_i_data_5(reductionMux_io_i_data_5),
    .io_i_sel(reductionMux_io_i_sel),
    .io_o_data_0(reductionMux_io_o_data_0),
    .io_o_data_1(reductionMux_io_o_data_1)
  );
  SimpleAdder adder32 ( // @[EdgeAdderSwitch.scala 27:23]
    .io_A(adder32_io_A),
    .io_B(adder32_io_B),
    .io_O(adder32_io_O)
  );
  assign io_o_vn = reset ? 64'h0 : r_vn; // @[EdgeAdderSwitch.scala 63:14 65:13 73:13]
  assign io_o_vn_valid = reset ? 2'h0 : r_vn_valid; // @[EdgeAdderSwitch.scala 63:14 66:19 74:19]
  assign io_o_adder = reset ? 32'h0 : _GEN_15; // @[EdgeAdderSwitch.scala 63:14 64:16]
  assign reductionMux_io_i_data_0 = io_i_data_bus_0[31:0]; // @[EdgeAdderSwitch.scala 24:26]
  assign reductionMux_io_i_data_1 = io_i_data_bus_1[31:0]; // @[EdgeAdderSwitch.scala 24:26]
  assign reductionMux_io_i_data_2 = io_i_data_bus_2[31:0]; // @[EdgeAdderSwitch.scala 24:26]
  assign reductionMux_io_i_data_3 = io_i_data_bus_3[31:0]; // @[EdgeAdderSwitch.scala 24:26]
  assign reductionMux_io_i_data_4 = io_i_data_bus_4[31:0]; // @[EdgeAdderSwitch.scala 24:26]
  assign reductionMux_io_i_data_5 = io_i_data_bus_5[31:0]; // @[EdgeAdderSwitch.scala 24:26]
  assign reductionMux_io_i_sel = io_i_sel; // @[EdgeAdderSwitch.scala 25:25]
  assign adder32_io_A = reductionMux_io_o_data_1; // @[EdgeAdderSwitch.scala 28:16]
  assign adder32_io_B = reductionMux_io_o_data_0; // @[EdgeAdderSwitch.scala 29:16]
  always @(posedge clock) begin
    if (reset) begin // @[EdgeAdderSwitch.scala 31:24]
      r_valid <= 1'h0; // @[EdgeAdderSwitch.scala 31:24]
    end else begin
      r_valid <= io_i_valid; // @[EdgeAdderSwitch.scala 31:24]
    end
    if (reset) begin // @[EdgeAdderSwitch.scala 32:24]
      r_adder <= 32'h0; // @[EdgeAdderSwitch.scala 32:24]
    end else if (reset) begin // @[EdgeAdderSwitch.scala 37:14]
      r_adder <= 32'h0; // @[EdgeAdderSwitch.scala 38:13]
    end else if (r_valid) begin // @[EdgeAdderSwitch.scala 41:25]
      if (5'h3 == io_i_cmd) begin // @[EdgeAdderSwitch.scala 42:23]
        r_adder <= reductionMux_io_o_data_1; // @[EdgeAdderSwitch.scala 44:17]
      end else begin
        r_adder <= _GEN_3;
      end
    end
    r_vn <= _GEN_19[63:0]; // @[EdgeAdderSwitch.scala 33:{21,21}]
    if (reset) begin // @[EdgeAdderSwitch.scala 34:27]
      r_vn_valid <= 2'h0; // @[EdgeAdderSwitch.scala 34:27]
    end else if (reset) begin // @[EdgeAdderSwitch.scala 37:14]
      r_vn_valid <= 2'h0; // @[EdgeAdderSwitch.scala 40:16]
    end else if (r_valid) begin // @[EdgeAdderSwitch.scala 41:25]
      if (5'h3 == io_i_cmd) begin // @[EdgeAdderSwitch.scala 42:23]
        r_vn_valid <= 2'h1; // @[EdgeAdderSwitch.scala 46:20]
      end else begin
        r_vn_valid <= _GEN_5;
      end
    end
    if (reset) begin // @[EdgeAdderSwitch.scala 35:25]
      r_add_en <= 3'h0; // @[EdgeAdderSwitch.scala 35:25]
    end else begin
      r_add_en <= io_i_add_en; // @[EdgeAdderSwitch.scala 35:25]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  r_adder = _RAND_1[31:0];
  _RAND_2 = {2{`RANDOM}};
  r_vn = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  r_vn_valid = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  r_add_en = _RAND_4[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AdderSwitch_7(
  input         clock,
  input         reset,
  input         io_i_valid,
  input  [31:0] io_i_data_bus_0,
  input  [31:0] io_i_data_bus_1,
  input  [31:0] io_i_data_bus_2,
  input  [31:0] io_i_data_bus_3,
  input  [2:0]  io_i_add_en,
  input  [2:0]  io_i_cmd,
  input  [1:0]  io_i_sel,
  output [1:0]  io_o_vn_valid,
  output [63:0] io_o_vn,
  output [31:0] io_o_adder_0,
  output [31:0] io_o_adder_1
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] reductionMux_io_i_data_0; // @[AdderSwitch.scala 25:28]
  wire [31:0] reductionMux_io_i_data_1; // @[AdderSwitch.scala 25:28]
  wire [31:0] reductionMux_io_i_data_2; // @[AdderSwitch.scala 25:28]
  wire [31:0] reductionMux_io_i_data_3; // @[AdderSwitch.scala 25:28]
  wire [1:0] reductionMux_io_i_sel; // @[AdderSwitch.scala 25:28]
  wire [31:0] reductionMux_io_o_data_0; // @[AdderSwitch.scala 25:28]
  wire [31:0] reductionMux_io_o_data_1; // @[AdderSwitch.scala 25:28]
  wire [31:0] adder32_io_A; // @[AdderSwitch.scala 29:23]
  wire [31:0] adder32_io_B; // @[AdderSwitch.scala 29:23]
  wire [31:0] adder32_io_O; // @[AdderSwitch.scala 29:23]
  reg [63:0] r_adder; // @[AdderSwitch.scala 33:24]
  reg [63:0] r_vn; // @[AdderSwitch.scala 34:21]
  reg [1:0] r_vn_valid; // @[AdderSwitch.scala 35:27]
  reg [2:0] r_add_en; // @[AdderSwitch.scala 36:25]
  wire [63:0] _r_adder_T = {reductionMux_io_o_data_0,reductionMux_io_o_data_1}; // @[Cat.scala 33:92]
  wire [62:0] _r_adder_T_1 = {31'h0,reductionMux_io_o_data_1}; // @[Cat.scala 33:92]
  wire [62:0] _r_adder_T_2 = {reductionMux_io_o_data_0,31'h0}; // @[Cat.scala 33:92]
  wire [1:0] _GEN_0 = 3'h0 == io_i_cmd ? 2'h0 : r_vn_valid; // @[AdderSwitch.scala 43:23 63:20 35:27]
  wire [63:0] _GEN_1 = 3'h5 == io_i_cmd ? _r_adder_T : r_vn; // @[AdderSwitch.scala 43:23 59:14 34:21]
  wire [1:0] _GEN_2 = 3'h5 == io_i_cmd ? 2'h3 : _GEN_0; // @[AdderSwitch.scala 43:23 60:20]
  wire [63:0] _GEN_3 = 3'h4 == io_i_cmd ? {{1'd0}, _r_adder_T_2} : r_adder; // @[AdderSwitch.scala 43:23 54:17 33:24]
  wire [63:0] _GEN_4 = 3'h4 == io_i_cmd ? {{32'd0}, io_i_data_bus_1} : _GEN_1; // @[AdderSwitch.scala 43:23 55:14]
  wire [1:0] _GEN_5 = 3'h4 == io_i_cmd ? 2'h2 : _GEN_2; // @[AdderSwitch.scala 43:23 56:20]
  wire [63:0] _GEN_6 = 3'h3 == io_i_cmd ? {{1'd0}, _r_adder_T_1} : _GEN_3; // @[AdderSwitch.scala 43:23 49:17]
  wire [63:0] _GEN_7 = 3'h3 == io_i_cmd ? {{32'd0}, io_i_data_bus_0} : _GEN_4; // @[AdderSwitch.scala 43:23 50:14]
  wire [1:0] _GEN_8 = 3'h3 == io_i_cmd ? 2'h1 : _GEN_5; // @[AdderSwitch.scala 43:23 51:20]
  wire [31:0] _WIRE_2_0 = adder32_io_O; // @[AdderSwitch.scala 76:{28,28}]
  wire [31:0] _GEN_18 = r_add_en == 3'h0 ? r_adder[31:0] : _WIRE_2_0; // @[AdderSwitch.scala 73:22 74:18 76:18]
  wire [31:0] _GEN_19 = r_add_en == 3'h0 ? r_adder[63:32] : _WIRE_2_0; // @[AdderSwitch.scala 73:22 74:18 76:18]
  ReductionMux_3 reductionMux ( // @[AdderSwitch.scala 25:28]
    .io_i_data_0(reductionMux_io_i_data_0),
    .io_i_data_1(reductionMux_io_i_data_1),
    .io_i_data_2(reductionMux_io_i_data_2),
    .io_i_data_3(reductionMux_io_i_data_3),
    .io_i_sel(reductionMux_io_i_sel),
    .io_o_data_0(reductionMux_io_o_data_0),
    .io_o_data_1(reductionMux_io_o_data_1)
  );
  SimpleAdder adder32 ( // @[AdderSwitch.scala 29:23]
    .io_A(adder32_io_A),
    .io_B(adder32_io_B),
    .io_O(adder32_io_O)
  );
  assign io_o_vn_valid = reset ? 2'h0 : r_vn_valid; // @[AdderSwitch.scala 68:14 71:19 79:19]
  assign io_o_vn = reset ? 64'h0 : r_vn; // @[AdderSwitch.scala 68:14 70:13 78:13]
  assign io_o_adder_0 = reset ? 32'h0 : _GEN_18; // @[AdderSwitch.scala 68:14 69:16]
  assign io_o_adder_1 = reset ? 32'h0 : _GEN_19; // @[AdderSwitch.scala 68:14 69:16]
  assign reductionMux_io_i_data_0 = io_i_data_bus_0; // @[AdderSwitch.scala 26:26]
  assign reductionMux_io_i_data_1 = io_i_data_bus_1; // @[AdderSwitch.scala 26:26]
  assign reductionMux_io_i_data_2 = io_i_data_bus_2; // @[AdderSwitch.scala 26:26]
  assign reductionMux_io_i_data_3 = io_i_data_bus_3; // @[AdderSwitch.scala 26:26]
  assign reductionMux_io_i_sel = io_i_sel; // @[AdderSwitch.scala 27:25]
  assign adder32_io_A = reductionMux_io_o_data_1; // @[AdderSwitch.scala 30:16]
  assign adder32_io_B = reductionMux_io_o_data_0; // @[AdderSwitch.scala 31:16]
  always @(posedge clock) begin
    if (reset) begin // @[AdderSwitch.scala 33:24]
      r_adder <= 64'h0; // @[AdderSwitch.scala 33:24]
    end else if (reset) begin // @[AdderSwitch.scala 38:14]
      r_adder <= 64'h0; // @[AdderSwitch.scala 39:13]
    end else if (io_i_valid) begin // @[AdderSwitch.scala 42:28]
      if (3'h1 == io_i_cmd) begin // @[AdderSwitch.scala 43:23]
        r_adder <= _r_adder_T; // @[AdderSwitch.scala 45:17]
      end else begin
        r_adder <= _GEN_6;
      end
    end
    if (reset) begin // @[AdderSwitch.scala 34:21]
      r_vn <= 64'h0; // @[AdderSwitch.scala 34:21]
    end else if (reset) begin // @[AdderSwitch.scala 38:14]
      r_vn <= 64'h0; // @[AdderSwitch.scala 40:10]
    end else if (io_i_valid) begin // @[AdderSwitch.scala 42:28]
      if (!(3'h1 == io_i_cmd)) begin // @[AdderSwitch.scala 43:23]
        r_vn <= _GEN_7;
      end
    end
    if (reset) begin // @[AdderSwitch.scala 35:27]
      r_vn_valid <= 2'h0; // @[AdderSwitch.scala 35:27]
    end else if (reset) begin // @[AdderSwitch.scala 38:14]
      r_vn_valid <= 2'h0; // @[AdderSwitch.scala 41:16]
    end else if (io_i_valid) begin // @[AdderSwitch.scala 42:28]
      if (3'h1 == io_i_cmd) begin // @[AdderSwitch.scala 43:23]
        r_vn_valid <= 2'h0; // @[AdderSwitch.scala 46:20]
      end else begin
        r_vn_valid <= _GEN_8;
      end
    end
    if (reset) begin // @[AdderSwitch.scala 36:25]
      r_add_en <= 3'h0; // @[AdderSwitch.scala 36:25]
    end else begin
      r_add_en <= io_i_add_en; // @[AdderSwitch.scala 36:25]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  r_adder = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  r_vn = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  r_vn_valid = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  r_add_en = _RAND_3[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ReductionMux_15(
  input  [31:0] io_i_data_0,
  input  [31:0] io_i_data_1,
  input  [31:0] io_i_data_2,
  input  [31:0] io_i_data_3,
  input  [31:0] io_i_data_4,
  input  [31:0] io_i_data_5,
  input  [31:0] io_i_data_6,
  input  [31:0] io_i_data_7,
  input  [3:0]  io_i_sel,
  output [31:0] io_o_data_0,
  output [31:0] io_o_data_1
);
  wire [1:0] w_sel_in_left = io_i_sel[1:0]; // @[ReductionMux.scala 29:32]
  wire [1:0] w_sel_in_right = io_i_sel[3:2]; // @[ReductionMux.scala 30:33]
  wire [31:0] _GEN_1 = 2'h1 == w_sel_in_left ? io_i_data_1 : io_i_data_0; // @[ReductionMux.scala 35:{18,18}]
  wire [31:0] _GEN_2 = 2'h2 == w_sel_in_left ? io_i_data_2 : _GEN_1; // @[ReductionMux.scala 35:{18,18}]
  wire [31:0] _GEN_3 = 2'h3 == w_sel_in_left ? io_i_data_3 : _GEN_2; // @[ReductionMux.scala 35:{18,18}]
  wire [31:0] _GEN_6 = 2'h1 == w_sel_in_right ? io_i_data_5 : io_i_data_4; // @[ReductionMux.scala 39:{22,22}]
  wire [31:0] _GEN_7 = 2'h2 == w_sel_in_right ? io_i_data_6 : _GEN_6; // @[ReductionMux.scala 39:{22,22}]
  assign io_o_data_0 = w_sel_in_left < 2'h2 ? _GEN_3 : 32'h0; // @[ReductionMux.scala 33:39 35:18 37:18]
  assign io_o_data_1 = 2'h3 == w_sel_in_right ? io_i_data_7 : _GEN_7; // @[ReductionMux.scala 39:{22,22}]
endmodule
module EdgeAdderSwitch_4(
  input         clock,
  input         reset,
  input         io_i_valid,
  input  [63:0] io_i_data_bus_0,
  input  [63:0] io_i_data_bus_1,
  input  [63:0] io_i_data_bus_2,
  input  [63:0] io_i_data_bus_3,
  input  [63:0] io_i_data_bus_4,
  input  [63:0] io_i_data_bus_5,
  input  [63:0] io_i_data_bus_6,
  input  [63:0] io_i_data_bus_7,
  input  [2:0]  io_i_add_en,
  input  [4:0]  io_i_cmd,
  input  [3:0]  io_i_sel,
  output [63:0] io_o_vn,
  output [1:0]  io_o_vn_valid,
  output [31:0] io_o_adder
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] reductionMux_io_i_data_0; // @[EdgeAdderSwitch.scala 23:28]
  wire [31:0] reductionMux_io_i_data_1; // @[EdgeAdderSwitch.scala 23:28]
  wire [31:0] reductionMux_io_i_data_2; // @[EdgeAdderSwitch.scala 23:28]
  wire [31:0] reductionMux_io_i_data_3; // @[EdgeAdderSwitch.scala 23:28]
  wire [31:0] reductionMux_io_i_data_4; // @[EdgeAdderSwitch.scala 23:28]
  wire [31:0] reductionMux_io_i_data_5; // @[EdgeAdderSwitch.scala 23:28]
  wire [31:0] reductionMux_io_i_data_6; // @[EdgeAdderSwitch.scala 23:28]
  wire [31:0] reductionMux_io_i_data_7; // @[EdgeAdderSwitch.scala 23:28]
  wire [3:0] reductionMux_io_i_sel; // @[EdgeAdderSwitch.scala 23:28]
  wire [31:0] reductionMux_io_o_data_0; // @[EdgeAdderSwitch.scala 23:28]
  wire [31:0] reductionMux_io_o_data_1; // @[EdgeAdderSwitch.scala 23:28]
  wire [31:0] adder32_io_A; // @[EdgeAdderSwitch.scala 27:23]
  wire [31:0] adder32_io_B; // @[EdgeAdderSwitch.scala 27:23]
  wire [31:0] adder32_io_O; // @[EdgeAdderSwitch.scala 27:23]
  reg  r_valid; // @[EdgeAdderSwitch.scala 31:24]
  reg [31:0] r_adder; // @[EdgeAdderSwitch.scala 32:24]
  reg [63:0] r_vn; // @[EdgeAdderSwitch.scala 33:21]
  reg [1:0] r_vn_valid; // @[EdgeAdderSwitch.scala 34:27]
  reg [2:0] r_add_en; // @[EdgeAdderSwitch.scala 35:25]
  wire [95:0] _r_vn_T = {io_i_data_bus_0,32'h0}; // @[Cat.scala 33:92]
  wire [95:0] _r_vn_T_1 = {32'h0,io_i_data_bus_7}; // @[Cat.scala 33:92]
  wire [63:0] _r_vn_T_2 = {reductionMux_io_o_data_0,reductionMux_io_o_data_1}; // @[Cat.scala 33:92]
  wire [1:0] _GEN_0 = 5'h0 == io_i_cmd ? 2'h0 : r_vn_valid; // @[EdgeAdderSwitch.scala 42:23 58:20 34:27]
  wire [63:0] _GEN_1 = 5'h5 == io_i_cmd ? _r_vn_T_2 : r_vn; // @[EdgeAdderSwitch.scala 42:23 54:14 33:21]
  wire [1:0] _GEN_2 = 5'h5 == io_i_cmd ? 2'h3 : _GEN_0; // @[EdgeAdderSwitch.scala 42:23 55:20]
  wire [31:0] _GEN_3 = 5'h4 == io_i_cmd ? reductionMux_io_o_data_0 : r_adder; // @[EdgeAdderSwitch.scala 42:23 49:17 32:24]
  wire [95:0] _GEN_4 = 5'h4 == io_i_cmd ? _r_vn_T_1 : {{32'd0}, _GEN_1}; // @[EdgeAdderSwitch.scala 42:23 50:14]
  wire [1:0] _GEN_5 = 5'h4 == io_i_cmd ? 2'h2 : _GEN_2; // @[EdgeAdderSwitch.scala 42:23 51:20]
  wire [95:0] _GEN_7 = 5'h3 == io_i_cmd ? _r_vn_T : _GEN_4; // @[EdgeAdderSwitch.scala 42:23 45:14]
  wire [95:0] _GEN_10 = r_valid ? _GEN_7 : {{32'd0}, r_vn}; // @[EdgeAdderSwitch.scala 33:21 41:25]
  wire [95:0] _GEN_13 = reset ? 96'h0 : _GEN_10; // @[EdgeAdderSwitch.scala 37:14 39:10]
  wire [31:0] _GEN_15 = r_add_en == 3'h0 ? r_adder : adder32_io_O; // @[EdgeAdderSwitch.scala 68:22 69:18 71:18]
  wire [95:0] _GEN_19 = reset ? 96'h0 : _GEN_13; // @[EdgeAdderSwitch.scala 33:{21,21}]
  ReductionMux_15 reductionMux ( // @[EdgeAdderSwitch.scala 23:28]
    .io_i_data_0(reductionMux_io_i_data_0),
    .io_i_data_1(reductionMux_io_i_data_1),
    .io_i_data_2(reductionMux_io_i_data_2),
    .io_i_data_3(reductionMux_io_i_data_3),
    .io_i_data_4(reductionMux_io_i_data_4),
    .io_i_data_5(reductionMux_io_i_data_5),
    .io_i_data_6(reductionMux_io_i_data_6),
    .io_i_data_7(reductionMux_io_i_data_7),
    .io_i_sel(reductionMux_io_i_sel),
    .io_o_data_0(reductionMux_io_o_data_0),
    .io_o_data_1(reductionMux_io_o_data_1)
  );
  SimpleAdder adder32 ( // @[EdgeAdderSwitch.scala 27:23]
    .io_A(adder32_io_A),
    .io_B(adder32_io_B),
    .io_O(adder32_io_O)
  );
  assign io_o_vn = reset ? 64'h0 : r_vn; // @[EdgeAdderSwitch.scala 63:14 65:13 73:13]
  assign io_o_vn_valid = reset ? 2'h0 : r_vn_valid; // @[EdgeAdderSwitch.scala 63:14 66:19 74:19]
  assign io_o_adder = reset ? 32'h0 : _GEN_15; // @[EdgeAdderSwitch.scala 63:14 64:16]
  assign reductionMux_io_i_data_0 = io_i_data_bus_0[31:0]; // @[EdgeAdderSwitch.scala 24:26]
  assign reductionMux_io_i_data_1 = io_i_data_bus_1[31:0]; // @[EdgeAdderSwitch.scala 24:26]
  assign reductionMux_io_i_data_2 = io_i_data_bus_2[31:0]; // @[EdgeAdderSwitch.scala 24:26]
  assign reductionMux_io_i_data_3 = io_i_data_bus_3[31:0]; // @[EdgeAdderSwitch.scala 24:26]
  assign reductionMux_io_i_data_4 = io_i_data_bus_4[31:0]; // @[EdgeAdderSwitch.scala 24:26]
  assign reductionMux_io_i_data_5 = io_i_data_bus_5[31:0]; // @[EdgeAdderSwitch.scala 24:26]
  assign reductionMux_io_i_data_6 = io_i_data_bus_6[31:0]; // @[EdgeAdderSwitch.scala 24:26]
  assign reductionMux_io_i_data_7 = io_i_data_bus_7[31:0]; // @[EdgeAdderSwitch.scala 24:26]
  assign reductionMux_io_i_sel = io_i_sel; // @[EdgeAdderSwitch.scala 25:25]
  assign adder32_io_A = reductionMux_io_o_data_1; // @[EdgeAdderSwitch.scala 28:16]
  assign adder32_io_B = reductionMux_io_o_data_0; // @[EdgeAdderSwitch.scala 29:16]
  always @(posedge clock) begin
    if (reset) begin // @[EdgeAdderSwitch.scala 31:24]
      r_valid <= 1'h0; // @[EdgeAdderSwitch.scala 31:24]
    end else begin
      r_valid <= io_i_valid; // @[EdgeAdderSwitch.scala 31:24]
    end
    if (reset) begin // @[EdgeAdderSwitch.scala 32:24]
      r_adder <= 32'h0; // @[EdgeAdderSwitch.scala 32:24]
    end else if (reset) begin // @[EdgeAdderSwitch.scala 37:14]
      r_adder <= 32'h0; // @[EdgeAdderSwitch.scala 38:13]
    end else if (r_valid) begin // @[EdgeAdderSwitch.scala 41:25]
      if (5'h3 == io_i_cmd) begin // @[EdgeAdderSwitch.scala 42:23]
        r_adder <= reductionMux_io_o_data_1; // @[EdgeAdderSwitch.scala 44:17]
      end else begin
        r_adder <= _GEN_3;
      end
    end
    r_vn <= _GEN_19[63:0]; // @[EdgeAdderSwitch.scala 33:{21,21}]
    if (reset) begin // @[EdgeAdderSwitch.scala 34:27]
      r_vn_valid <= 2'h0; // @[EdgeAdderSwitch.scala 34:27]
    end else if (reset) begin // @[EdgeAdderSwitch.scala 37:14]
      r_vn_valid <= 2'h0; // @[EdgeAdderSwitch.scala 40:16]
    end else if (r_valid) begin // @[EdgeAdderSwitch.scala 41:25]
      if (5'h3 == io_i_cmd) begin // @[EdgeAdderSwitch.scala 42:23]
        r_vn_valid <= 2'h1; // @[EdgeAdderSwitch.scala 46:20]
      end else begin
        r_vn_valid <= _GEN_5;
      end
    end
    if (reset) begin // @[EdgeAdderSwitch.scala 35:25]
      r_add_en <= 3'h0; // @[EdgeAdderSwitch.scala 35:25]
    end else begin
      r_add_en <= io_i_add_en; // @[EdgeAdderSwitch.scala 35:25]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  r_adder = _RAND_1[31:0];
  _RAND_2 = {2{`RANDOM}};
  r_vn = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  r_vn_valid = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  r_add_en = _RAND_4[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FanNetworkcom(
  input         clock,
  input         reset,
  input         io_i_valid,
  input  [31:0] io_i_data_bus_0,
  input  [31:0] io_i_data_bus_1,
  input  [31:0] io_i_data_bus_2,
  input  [31:0] io_i_data_bus_3,
  input  [31:0] io_i_data_bus_4,
  input  [31:0] io_i_data_bus_5,
  input  [31:0] io_i_data_bus_6,
  input  [31:0] io_i_data_bus_7,
  input  [31:0] io_i_data_bus_8,
  input  [31:0] io_i_data_bus_9,
  input  [31:0] io_i_data_bus_10,
  input  [31:0] io_i_data_bus_11,
  input  [31:0] io_i_data_bus_12,
  input  [31:0] io_i_data_bus_13,
  input  [31:0] io_i_data_bus_14,
  input  [31:0] io_i_data_bus_15,
  input  [31:0] io_i_data_bus_16,
  input  [31:0] io_i_data_bus_17,
  input  [31:0] io_i_data_bus_18,
  input  [31:0] io_i_data_bus_19,
  input  [31:0] io_i_data_bus_20,
  input  [31:0] io_i_data_bus_21,
  input  [31:0] io_i_data_bus_22,
  input  [31:0] io_i_data_bus_23,
  input  [31:0] io_i_data_bus_24,
  input  [31:0] io_i_data_bus_25,
  input  [31:0] io_i_data_bus_26,
  input  [31:0] io_i_data_bus_27,
  input  [31:0] io_i_data_bus_28,
  input  [31:0] io_i_data_bus_29,
  input  [31:0] io_i_data_bus_30,
  input  [31:0] io_i_data_bus_31,
  input         io_i_add_en_bus_0,
  input         io_i_add_en_bus_1,
  input         io_i_add_en_bus_2,
  input         io_i_add_en_bus_3,
  input         io_i_add_en_bus_4,
  input         io_i_add_en_bus_5,
  input         io_i_add_en_bus_6,
  input         io_i_add_en_bus_7,
  input         io_i_add_en_bus_8,
  input         io_i_add_en_bus_9,
  input         io_i_add_en_bus_10,
  input         io_i_add_en_bus_11,
  input         io_i_add_en_bus_12,
  input         io_i_add_en_bus_13,
  input         io_i_add_en_bus_14,
  input         io_i_add_en_bus_15,
  input         io_i_add_en_bus_16,
  input         io_i_add_en_bus_17,
  input         io_i_add_en_bus_18,
  input         io_i_add_en_bus_19,
  input         io_i_add_en_bus_20,
  input         io_i_add_en_bus_21,
  input         io_i_add_en_bus_22,
  input         io_i_add_en_bus_23,
  input         io_i_add_en_bus_24,
  input         io_i_add_en_bus_25,
  input         io_i_add_en_bus_26,
  input         io_i_add_en_bus_27,
  input         io_i_add_en_bus_28,
  input         io_i_add_en_bus_29,
  input         io_i_add_en_bus_30,
  input  [2:0]  io_i_cmd_bus_0,
  input  [2:0]  io_i_cmd_bus_1,
  input  [2:0]  io_i_cmd_bus_2,
  input  [2:0]  io_i_cmd_bus_3,
  input  [2:0]  io_i_cmd_bus_4,
  input  [2:0]  io_i_cmd_bus_5,
  input  [2:0]  io_i_cmd_bus_6,
  input  [2:0]  io_i_cmd_bus_7,
  input  [2:0]  io_i_cmd_bus_8,
  input  [2:0]  io_i_cmd_bus_9,
  input  [2:0]  io_i_cmd_bus_10,
  input  [2:0]  io_i_cmd_bus_11,
  input  [2:0]  io_i_cmd_bus_12,
  input  [2:0]  io_i_cmd_bus_13,
  input  [2:0]  io_i_cmd_bus_14,
  input  [2:0]  io_i_cmd_bus_15,
  input  [2:0]  io_i_cmd_bus_16,
  input  [2:0]  io_i_cmd_bus_17,
  input  [2:0]  io_i_cmd_bus_18,
  input  [2:0]  io_i_cmd_bus_19,
  input  [2:0]  io_i_cmd_bus_20,
  input  [2:0]  io_i_cmd_bus_21,
  input  [2:0]  io_i_cmd_bus_22,
  input  [2:0]  io_i_cmd_bus_23,
  input  [2:0]  io_i_cmd_bus_24,
  input  [2:0]  io_i_cmd_bus_25,
  input  [2:0]  io_i_cmd_bus_26,
  input  [2:0]  io_i_cmd_bus_27,
  input  [2:0]  io_i_cmd_bus_28,
  input  [2:0]  io_i_cmd_bus_29,
  input  [2:0]  io_i_cmd_bus_30,
  input         io_i_sel_bus_0,
  input         io_i_sel_bus_1,
  input         io_i_sel_bus_2,
  input         io_i_sel_bus_3,
  input         io_i_sel_bus_4,
  input         io_i_sel_bus_5,
  input         io_i_sel_bus_6,
  input         io_i_sel_bus_7,
  input         io_i_sel_bus_8,
  input         io_i_sel_bus_9,
  input         io_i_sel_bus_10,
  input         io_i_sel_bus_11,
  input         io_i_sel_bus_12,
  input         io_i_sel_bus_13,
  input         io_i_sel_bus_14,
  input         io_i_sel_bus_15,
  input         io_i_sel_bus_16,
  input         io_i_sel_bus_17,
  input         io_i_sel_bus_18,
  input         io_i_sel_bus_19,
  output        io_o_valid_0,
  output        io_o_valid_1,
  output        io_o_valid_2,
  output        io_o_valid_3,
  output        io_o_valid_4,
  output        io_o_valid_5,
  output        io_o_valid_6,
  output        io_o_valid_7,
  output        io_o_valid_8,
  output        io_o_valid_9,
  output        io_o_valid_10,
  output        io_o_valid_11,
  output        io_o_valid_12,
  output        io_o_valid_13,
  output        io_o_valid_14,
  output        io_o_valid_15,
  output        io_o_valid_16,
  output        io_o_valid_17,
  output        io_o_valid_18,
  output        io_o_valid_19,
  output        io_o_valid_20,
  output        io_o_valid_21,
  output        io_o_valid_22,
  output        io_o_valid_23,
  output        io_o_valid_24,
  output        io_o_valid_25,
  output        io_o_valid_26,
  output        io_o_valid_27,
  output        io_o_valid_28,
  output        io_o_valid_29,
  output        io_o_valid_30,
  output        io_o_valid_31,
  output [31:0] io_o_data_bus_0,
  output [31:0] io_o_data_bus_1,
  output [31:0] io_o_data_bus_2,
  output [31:0] io_o_data_bus_3,
  output [31:0] io_o_data_bus_4,
  output [31:0] io_o_data_bus_5,
  output [31:0] io_o_data_bus_6,
  output [31:0] io_o_data_bus_7,
  output [31:0] io_o_data_bus_8,
  output [31:0] io_o_data_bus_9,
  output [31:0] io_o_data_bus_10,
  output [31:0] io_o_data_bus_11,
  output [31:0] io_o_data_bus_12,
  output [31:0] io_o_data_bus_13,
  output [31:0] io_o_data_bus_14,
  output [31:0] io_o_data_bus_15,
  output [31:0] io_o_data_bus_16,
  output [31:0] io_o_data_bus_17,
  output [31:0] io_o_data_bus_18,
  output [31:0] io_o_data_bus_19,
  output [31:0] io_o_data_bus_20,
  output [31:0] io_o_data_bus_21,
  output [31:0] io_o_data_bus_22,
  output [31:0] io_o_data_bus_23,
  output [31:0] io_o_data_bus_24,
  output [31:0] io_o_data_bus_25,
  output [31:0] io_o_data_bus_26,
  output [31:0] io_o_data_bus_27,
  output [31:0] io_o_data_bus_28,
  output [31:0] io_o_data_bus_29,
  output [31:0] io_o_data_bus_30,
  output [31:0] io_o_data_bus_31
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
`endif // RANDOMIZE_REG_INIT
  wire  my_adder_0_clock; // @[FanNetwork.scala 1018:28]
  wire  my_adder_0_reset; // @[FanNetwork.scala 1018:28]
  wire  my_adder_0_io_i_valid; // @[FanNetwork.scala 1018:28]
  wire [63:0] my_adder_0_io_i_data_bus_0; // @[FanNetwork.scala 1018:28]
  wire [63:0] my_adder_0_io_i_data_bus_1; // @[FanNetwork.scala 1018:28]
  wire [2:0] my_adder_0_io_i_add_en; // @[FanNetwork.scala 1018:28]
  wire [4:0] my_adder_0_io_i_cmd; // @[FanNetwork.scala 1018:28]
  wire [63:0] my_adder_0_io_o_vn; // @[FanNetwork.scala 1018:28]
  wire [1:0] my_adder_0_io_o_vn_valid; // @[FanNetwork.scala 1018:28]
  wire [31:0] my_adder_0_io_o_adder; // @[FanNetwork.scala 1018:28]
  wire  my_adder_1_clock; // @[FanNetwork.scala 1031:28]
  wire  my_adder_1_reset; // @[FanNetwork.scala 1031:28]
  wire  my_adder_1_io_i_valid; // @[FanNetwork.scala 1031:28]
  wire [63:0] my_adder_1_io_i_data_bus_0; // @[FanNetwork.scala 1031:28]
  wire [63:0] my_adder_1_io_i_data_bus_1; // @[FanNetwork.scala 1031:28]
  wire [2:0] my_adder_1_io_i_add_en; // @[FanNetwork.scala 1031:28]
  wire [4:0] my_adder_1_io_i_cmd; // @[FanNetwork.scala 1031:28]
  wire [63:0] my_adder_1_io_o_vn; // @[FanNetwork.scala 1031:28]
  wire [1:0] my_adder_1_io_o_vn_valid; // @[FanNetwork.scala 1031:28]
  wire [31:0] my_adder_1_io_o_adder; // @[FanNetwork.scala 1031:28]
  wire  my_adder_2_clock; // @[FanNetwork.scala 1045:28]
  wire  my_adder_2_reset; // @[FanNetwork.scala 1045:28]
  wire  my_adder_2_io_i_valid; // @[FanNetwork.scala 1045:28]
  wire [31:0] my_adder_2_io_i_data_bus_0; // @[FanNetwork.scala 1045:28]
  wire [31:0] my_adder_2_io_i_data_bus_1; // @[FanNetwork.scala 1045:28]
  wire [2:0] my_adder_2_io_i_add_en; // @[FanNetwork.scala 1045:28]
  wire [2:0] my_adder_2_io_i_cmd; // @[FanNetwork.scala 1045:28]
  wire [1:0] my_adder_2_io_o_vn_valid; // @[FanNetwork.scala 1045:28]
  wire [63:0] my_adder_2_io_o_vn; // @[FanNetwork.scala 1045:28]
  wire [31:0] my_adder_2_io_o_adder_0; // @[FanNetwork.scala 1045:28]
  wire [31:0] my_adder_2_io_o_adder_1; // @[FanNetwork.scala 1045:28]
  wire  my_adder_3_clock; // @[FanNetwork.scala 1064:28]
  wire  my_adder_3_reset; // @[FanNetwork.scala 1064:28]
  wire  my_adder_3_io_i_valid; // @[FanNetwork.scala 1064:28]
  wire [63:0] my_adder_3_io_i_data_bus_0; // @[FanNetwork.scala 1064:28]
  wire [63:0] my_adder_3_io_i_data_bus_1; // @[FanNetwork.scala 1064:28]
  wire [63:0] my_adder_3_io_i_data_bus_2; // @[FanNetwork.scala 1064:28]
  wire [63:0] my_adder_3_io_i_data_bus_3; // @[FanNetwork.scala 1064:28]
  wire [2:0] my_adder_3_io_i_add_en; // @[FanNetwork.scala 1064:28]
  wire [4:0] my_adder_3_io_i_cmd; // @[FanNetwork.scala 1064:28]
  wire [1:0] my_adder_3_io_i_sel; // @[FanNetwork.scala 1064:28]
  wire [63:0] my_adder_3_io_o_vn; // @[FanNetwork.scala 1064:28]
  wire [1:0] my_adder_3_io_o_vn_valid; // @[FanNetwork.scala 1064:28]
  wire [31:0] my_adder_3_io_o_adder; // @[FanNetwork.scala 1064:28]
  wire  my_adder_4_clock; // @[FanNetwork.scala 1081:28]
  wire  my_adder_4_reset; // @[FanNetwork.scala 1081:28]
  wire  my_adder_4_io_i_valid; // @[FanNetwork.scala 1081:28]
  wire [31:0] my_adder_4_io_i_data_bus_0; // @[FanNetwork.scala 1081:28]
  wire [31:0] my_adder_4_io_i_data_bus_1; // @[FanNetwork.scala 1081:28]
  wire [2:0] my_adder_4_io_i_add_en; // @[FanNetwork.scala 1081:28]
  wire [2:0] my_adder_4_io_i_cmd; // @[FanNetwork.scala 1081:28]
  wire [1:0] my_adder_4_io_o_vn_valid; // @[FanNetwork.scala 1081:28]
  wire [63:0] my_adder_4_io_o_vn; // @[FanNetwork.scala 1081:28]
  wire [31:0] my_adder_4_io_o_adder_0; // @[FanNetwork.scala 1081:28]
  wire [31:0] my_adder_4_io_o_adder_1; // @[FanNetwork.scala 1081:28]
  wire  my_adder_5_clock; // @[FanNetwork.scala 1099:28]
  wire  my_adder_5_reset; // @[FanNetwork.scala 1099:28]
  wire  my_adder_5_io_i_valid; // @[FanNetwork.scala 1099:28]
  wire [31:0] my_adder_5_io_i_data_bus_0; // @[FanNetwork.scala 1099:28]
  wire [31:0] my_adder_5_io_i_data_bus_1; // @[FanNetwork.scala 1099:28]
  wire [2:0] my_adder_5_io_i_add_en; // @[FanNetwork.scala 1099:28]
  wire [2:0] my_adder_5_io_i_cmd; // @[FanNetwork.scala 1099:28]
  wire [1:0] my_adder_5_io_o_vn_valid; // @[FanNetwork.scala 1099:28]
  wire [63:0] my_adder_5_io_o_vn; // @[FanNetwork.scala 1099:28]
  wire [31:0] my_adder_5_io_o_adder_0; // @[FanNetwork.scala 1099:28]
  wire [31:0] my_adder_5_io_o_adder_1; // @[FanNetwork.scala 1099:28]
  wire  my_adder_6_clock; // @[FanNetwork.scala 1116:28]
  wire  my_adder_6_reset; // @[FanNetwork.scala 1116:28]
  wire  my_adder_6_io_i_valid; // @[FanNetwork.scala 1116:28]
  wire [31:0] my_adder_6_io_i_data_bus_0; // @[FanNetwork.scala 1116:28]
  wire [31:0] my_adder_6_io_i_data_bus_1; // @[FanNetwork.scala 1116:28]
  wire [2:0] my_adder_6_io_i_add_en; // @[FanNetwork.scala 1116:28]
  wire [2:0] my_adder_6_io_i_cmd; // @[FanNetwork.scala 1116:28]
  wire [1:0] my_adder_6_io_o_vn_valid; // @[FanNetwork.scala 1116:28]
  wire [63:0] my_adder_6_io_o_vn; // @[FanNetwork.scala 1116:28]
  wire [31:0] my_adder_6_io_o_adder_0; // @[FanNetwork.scala 1116:28]
  wire [31:0] my_adder_6_io_o_adder_1; // @[FanNetwork.scala 1116:28]
  wire  my_adder_7_clock; // @[FanNetwork.scala 1133:28]
  wire  my_adder_7_reset; // @[FanNetwork.scala 1133:28]
  wire  my_adder_7_io_i_valid; // @[FanNetwork.scala 1133:28]
  wire [63:0] my_adder_7_io_i_data_bus_0; // @[FanNetwork.scala 1133:28]
  wire [63:0] my_adder_7_io_i_data_bus_1; // @[FanNetwork.scala 1133:28]
  wire [63:0] my_adder_7_io_i_data_bus_2; // @[FanNetwork.scala 1133:28]
  wire [63:0] my_adder_7_io_i_data_bus_3; // @[FanNetwork.scala 1133:28]
  wire [63:0] my_adder_7_io_i_data_bus_4; // @[FanNetwork.scala 1133:28]
  wire [63:0] my_adder_7_io_i_data_bus_5; // @[FanNetwork.scala 1133:28]
  wire [2:0] my_adder_7_io_i_add_en; // @[FanNetwork.scala 1133:28]
  wire [4:0] my_adder_7_io_i_cmd; // @[FanNetwork.scala 1133:28]
  wire [3:0] my_adder_7_io_i_sel; // @[FanNetwork.scala 1133:28]
  wire [63:0] my_adder_7_io_o_vn; // @[FanNetwork.scala 1133:28]
  wire [1:0] my_adder_7_io_o_vn_valid; // @[FanNetwork.scala 1133:28]
  wire [31:0] my_adder_7_io_o_adder; // @[FanNetwork.scala 1133:28]
  wire  my_adder_8_clock; // @[FanNetwork.scala 1152:28]
  wire  my_adder_8_reset; // @[FanNetwork.scala 1152:28]
  wire  my_adder_8_io_i_valid; // @[FanNetwork.scala 1152:28]
  wire [31:0] my_adder_8_io_i_data_bus_0; // @[FanNetwork.scala 1152:28]
  wire [31:0] my_adder_8_io_i_data_bus_1; // @[FanNetwork.scala 1152:28]
  wire [2:0] my_adder_8_io_i_add_en; // @[FanNetwork.scala 1152:28]
  wire [2:0] my_adder_8_io_i_cmd; // @[FanNetwork.scala 1152:28]
  wire [1:0] my_adder_8_io_o_vn_valid; // @[FanNetwork.scala 1152:28]
  wire [63:0] my_adder_8_io_o_vn; // @[FanNetwork.scala 1152:28]
  wire [31:0] my_adder_8_io_o_adder_0; // @[FanNetwork.scala 1152:28]
  wire [31:0] my_adder_8_io_o_adder_1; // @[FanNetwork.scala 1152:28]
  wire  my_adder_9_clock; // @[FanNetwork.scala 1169:28]
  wire  my_adder_9_reset; // @[FanNetwork.scala 1169:28]
  wire  my_adder_9_io_i_valid; // @[FanNetwork.scala 1169:28]
  wire [31:0] my_adder_9_io_i_data_bus_0; // @[FanNetwork.scala 1169:28]
  wire [31:0] my_adder_9_io_i_data_bus_1; // @[FanNetwork.scala 1169:28]
  wire [2:0] my_adder_9_io_i_add_en; // @[FanNetwork.scala 1169:28]
  wire [2:0] my_adder_9_io_i_cmd; // @[FanNetwork.scala 1169:28]
  wire [1:0] my_adder_9_io_o_vn_valid; // @[FanNetwork.scala 1169:28]
  wire [63:0] my_adder_9_io_o_vn; // @[FanNetwork.scala 1169:28]
  wire [31:0] my_adder_9_io_o_adder_0; // @[FanNetwork.scala 1169:28]
  wire [31:0] my_adder_9_io_o_adder_1; // @[FanNetwork.scala 1169:28]
  wire  my_adder_10_clock; // @[FanNetwork.scala 1186:29]
  wire  my_adder_10_reset; // @[FanNetwork.scala 1186:29]
  wire  my_adder_10_io_i_valid; // @[FanNetwork.scala 1186:29]
  wire [31:0] my_adder_10_io_i_data_bus_0; // @[FanNetwork.scala 1186:29]
  wire [31:0] my_adder_10_io_i_data_bus_1; // @[FanNetwork.scala 1186:29]
  wire [2:0] my_adder_10_io_i_add_en; // @[FanNetwork.scala 1186:29]
  wire [2:0] my_adder_10_io_i_cmd; // @[FanNetwork.scala 1186:29]
  wire [1:0] my_adder_10_io_o_vn_valid; // @[FanNetwork.scala 1186:29]
  wire [63:0] my_adder_10_io_o_vn; // @[FanNetwork.scala 1186:29]
  wire [31:0] my_adder_10_io_o_adder_0; // @[FanNetwork.scala 1186:29]
  wire [31:0] my_adder_10_io_o_adder_1; // @[FanNetwork.scala 1186:29]
  wire  my_adder_11_clock; // @[FanNetwork.scala 1204:29]
  wire  my_adder_11_reset; // @[FanNetwork.scala 1204:29]
  wire  my_adder_11_io_i_valid; // @[FanNetwork.scala 1204:29]
  wire [31:0] my_adder_11_io_i_data_bus_0; // @[FanNetwork.scala 1204:29]
  wire [31:0] my_adder_11_io_i_data_bus_1; // @[FanNetwork.scala 1204:29]
  wire [31:0] my_adder_11_io_i_data_bus_2; // @[FanNetwork.scala 1204:29]
  wire [31:0] my_adder_11_io_i_data_bus_3; // @[FanNetwork.scala 1204:29]
  wire [2:0] my_adder_11_io_i_add_en; // @[FanNetwork.scala 1204:29]
  wire [2:0] my_adder_11_io_i_cmd; // @[FanNetwork.scala 1204:29]
  wire [1:0] my_adder_11_io_i_sel; // @[FanNetwork.scala 1204:29]
  wire [1:0] my_adder_11_io_o_vn_valid; // @[FanNetwork.scala 1204:29]
  wire [63:0] my_adder_11_io_o_vn; // @[FanNetwork.scala 1204:29]
  wire [31:0] my_adder_11_io_o_adder_0; // @[FanNetwork.scala 1204:29]
  wire [31:0] my_adder_11_io_o_adder_1; // @[FanNetwork.scala 1204:29]
  wire  my_adder_12_clock; // @[FanNetwork.scala 1225:29]
  wire  my_adder_12_reset; // @[FanNetwork.scala 1225:29]
  wire  my_adder_12_io_i_valid; // @[FanNetwork.scala 1225:29]
  wire [31:0] my_adder_12_io_i_data_bus_0; // @[FanNetwork.scala 1225:29]
  wire [31:0] my_adder_12_io_i_data_bus_1; // @[FanNetwork.scala 1225:29]
  wire [2:0] my_adder_12_io_i_add_en; // @[FanNetwork.scala 1225:29]
  wire [2:0] my_adder_12_io_i_cmd; // @[FanNetwork.scala 1225:29]
  wire [1:0] my_adder_12_io_o_vn_valid; // @[FanNetwork.scala 1225:29]
  wire [63:0] my_adder_12_io_o_vn; // @[FanNetwork.scala 1225:29]
  wire [31:0] my_adder_12_io_o_adder_0; // @[FanNetwork.scala 1225:29]
  wire [31:0] my_adder_12_io_o_adder_1; // @[FanNetwork.scala 1225:29]
  wire  my_adder_13_clock; // @[FanNetwork.scala 1243:29]
  wire  my_adder_13_reset; // @[FanNetwork.scala 1243:29]
  wire  my_adder_13_io_i_valid; // @[FanNetwork.scala 1243:29]
  wire [31:0] my_adder_13_io_i_data_bus_0; // @[FanNetwork.scala 1243:29]
  wire [31:0] my_adder_13_io_i_data_bus_1; // @[FanNetwork.scala 1243:29]
  wire [2:0] my_adder_13_io_i_add_en; // @[FanNetwork.scala 1243:29]
  wire [2:0] my_adder_13_io_i_cmd; // @[FanNetwork.scala 1243:29]
  wire [1:0] my_adder_13_io_o_vn_valid; // @[FanNetwork.scala 1243:29]
  wire [63:0] my_adder_13_io_o_vn; // @[FanNetwork.scala 1243:29]
  wire [31:0] my_adder_13_io_o_adder_0; // @[FanNetwork.scala 1243:29]
  wire [31:0] my_adder_13_io_o_adder_1; // @[FanNetwork.scala 1243:29]
  wire  my_adder_14_clock; // @[FanNetwork.scala 1261:29]
  wire  my_adder_14_reset; // @[FanNetwork.scala 1261:29]
  wire  my_adder_14_io_i_valid; // @[FanNetwork.scala 1261:29]
  wire [31:0] my_adder_14_io_i_data_bus_0; // @[FanNetwork.scala 1261:29]
  wire [31:0] my_adder_14_io_i_data_bus_1; // @[FanNetwork.scala 1261:29]
  wire [2:0] my_adder_14_io_i_add_en; // @[FanNetwork.scala 1261:29]
  wire [2:0] my_adder_14_io_i_cmd; // @[FanNetwork.scala 1261:29]
  wire [1:0] my_adder_14_io_o_vn_valid; // @[FanNetwork.scala 1261:29]
  wire [63:0] my_adder_14_io_o_vn; // @[FanNetwork.scala 1261:29]
  wire [31:0] my_adder_14_io_o_adder_0; // @[FanNetwork.scala 1261:29]
  wire [31:0] my_adder_14_io_o_adder_1; // @[FanNetwork.scala 1261:29]
  wire  my_adder_15_clock; // @[FanNetwork.scala 1279:29]
  wire  my_adder_15_reset; // @[FanNetwork.scala 1279:29]
  wire  my_adder_15_io_i_valid; // @[FanNetwork.scala 1279:29]
  wire [63:0] my_adder_15_io_i_data_bus_0; // @[FanNetwork.scala 1279:29]
  wire [63:0] my_adder_15_io_i_data_bus_1; // @[FanNetwork.scala 1279:29]
  wire [63:0] my_adder_15_io_i_data_bus_2; // @[FanNetwork.scala 1279:29]
  wire [63:0] my_adder_15_io_i_data_bus_3; // @[FanNetwork.scala 1279:29]
  wire [63:0] my_adder_15_io_i_data_bus_4; // @[FanNetwork.scala 1279:29]
  wire [63:0] my_adder_15_io_i_data_bus_5; // @[FanNetwork.scala 1279:29]
  wire [63:0] my_adder_15_io_i_data_bus_6; // @[FanNetwork.scala 1279:29]
  wire [63:0] my_adder_15_io_i_data_bus_7; // @[FanNetwork.scala 1279:29]
  wire [2:0] my_adder_15_io_i_add_en; // @[FanNetwork.scala 1279:29]
  wire [4:0] my_adder_15_io_i_cmd; // @[FanNetwork.scala 1279:29]
  wire [3:0] my_adder_15_io_i_sel; // @[FanNetwork.scala 1279:29]
  wire [63:0] my_adder_15_io_o_vn; // @[FanNetwork.scala 1279:29]
  wire [1:0] my_adder_15_io_o_vn_valid; // @[FanNetwork.scala 1279:29]
  wire [31:0] my_adder_15_io_o_adder; // @[FanNetwork.scala 1279:29]
  wire  my_adder_16_clock; // @[FanNetwork.scala 1299:29]
  wire  my_adder_16_reset; // @[FanNetwork.scala 1299:29]
  wire  my_adder_16_io_i_valid; // @[FanNetwork.scala 1299:29]
  wire [31:0] my_adder_16_io_i_data_bus_0; // @[FanNetwork.scala 1299:29]
  wire [31:0] my_adder_16_io_i_data_bus_1; // @[FanNetwork.scala 1299:29]
  wire [2:0] my_adder_16_io_i_add_en; // @[FanNetwork.scala 1299:29]
  wire [2:0] my_adder_16_io_i_cmd; // @[FanNetwork.scala 1299:29]
  wire [1:0] my_adder_16_io_o_vn_valid; // @[FanNetwork.scala 1299:29]
  wire [63:0] my_adder_16_io_o_vn; // @[FanNetwork.scala 1299:29]
  wire [31:0] my_adder_16_io_o_adder_0; // @[FanNetwork.scala 1299:29]
  wire [31:0] my_adder_16_io_o_adder_1; // @[FanNetwork.scala 1299:29]
  wire  my_adder_17_clock; // @[FanNetwork.scala 1317:29]
  wire  my_adder_17_reset; // @[FanNetwork.scala 1317:29]
  wire  my_adder_17_io_i_valid; // @[FanNetwork.scala 1317:29]
  wire [31:0] my_adder_17_io_i_data_bus_0; // @[FanNetwork.scala 1317:29]
  wire [31:0] my_adder_17_io_i_data_bus_1; // @[FanNetwork.scala 1317:29]
  wire [2:0] my_adder_17_io_i_add_en; // @[FanNetwork.scala 1317:29]
  wire [2:0] my_adder_17_io_i_cmd; // @[FanNetwork.scala 1317:29]
  wire [1:0] my_adder_17_io_o_vn_valid; // @[FanNetwork.scala 1317:29]
  wire [63:0] my_adder_17_io_o_vn; // @[FanNetwork.scala 1317:29]
  wire [31:0] my_adder_17_io_o_adder_0; // @[FanNetwork.scala 1317:29]
  wire [31:0] my_adder_17_io_o_adder_1; // @[FanNetwork.scala 1317:29]
  wire  my_adder_18_clock; // @[FanNetwork.scala 1335:29]
  wire  my_adder_18_reset; // @[FanNetwork.scala 1335:29]
  wire  my_adder_18_io_i_valid; // @[FanNetwork.scala 1335:29]
  wire [31:0] my_adder_18_io_i_data_bus_0; // @[FanNetwork.scala 1335:29]
  wire [31:0] my_adder_18_io_i_data_bus_1; // @[FanNetwork.scala 1335:29]
  wire [2:0] my_adder_18_io_i_add_en; // @[FanNetwork.scala 1335:29]
  wire [2:0] my_adder_18_io_i_cmd; // @[FanNetwork.scala 1335:29]
  wire [1:0] my_adder_18_io_o_vn_valid; // @[FanNetwork.scala 1335:29]
  wire [63:0] my_adder_18_io_o_vn; // @[FanNetwork.scala 1335:29]
  wire [31:0] my_adder_18_io_o_adder_0; // @[FanNetwork.scala 1335:29]
  wire [31:0] my_adder_18_io_o_adder_1; // @[FanNetwork.scala 1335:29]
  wire  my_adder_19_clock; // @[FanNetwork.scala 1353:29]
  wire  my_adder_19_reset; // @[FanNetwork.scala 1353:29]
  wire  my_adder_19_io_i_valid; // @[FanNetwork.scala 1353:29]
  wire [31:0] my_adder_19_io_i_data_bus_0; // @[FanNetwork.scala 1353:29]
  wire [31:0] my_adder_19_io_i_data_bus_1; // @[FanNetwork.scala 1353:29]
  wire [31:0] my_adder_19_io_i_data_bus_2; // @[FanNetwork.scala 1353:29]
  wire [31:0] my_adder_19_io_i_data_bus_3; // @[FanNetwork.scala 1353:29]
  wire [2:0] my_adder_19_io_i_add_en; // @[FanNetwork.scala 1353:29]
  wire [2:0] my_adder_19_io_i_cmd; // @[FanNetwork.scala 1353:29]
  wire [1:0] my_adder_19_io_i_sel; // @[FanNetwork.scala 1353:29]
  wire [1:0] my_adder_19_io_o_vn_valid; // @[FanNetwork.scala 1353:29]
  wire [63:0] my_adder_19_io_o_vn; // @[FanNetwork.scala 1353:29]
  wire [31:0] my_adder_19_io_o_adder_0; // @[FanNetwork.scala 1353:29]
  wire [31:0] my_adder_19_io_o_adder_1; // @[FanNetwork.scala 1353:29]
  wire  my_adder_20_clock; // @[FanNetwork.scala 1373:29]
  wire  my_adder_20_reset; // @[FanNetwork.scala 1373:29]
  wire  my_adder_20_io_i_valid; // @[FanNetwork.scala 1373:29]
  wire [31:0] my_adder_20_io_i_data_bus_0; // @[FanNetwork.scala 1373:29]
  wire [31:0] my_adder_20_io_i_data_bus_1; // @[FanNetwork.scala 1373:29]
  wire [2:0] my_adder_20_io_i_add_en; // @[FanNetwork.scala 1373:29]
  wire [2:0] my_adder_20_io_i_cmd; // @[FanNetwork.scala 1373:29]
  wire [1:0] my_adder_20_io_o_vn_valid; // @[FanNetwork.scala 1373:29]
  wire [63:0] my_adder_20_io_o_vn; // @[FanNetwork.scala 1373:29]
  wire [31:0] my_adder_20_io_o_adder_0; // @[FanNetwork.scala 1373:29]
  wire [31:0] my_adder_20_io_o_adder_1; // @[FanNetwork.scala 1373:29]
  wire  my_adder_21_clock; // @[FanNetwork.scala 1393:29]
  wire  my_adder_21_reset; // @[FanNetwork.scala 1393:29]
  wire  my_adder_21_io_i_valid; // @[FanNetwork.scala 1393:29]
  wire [31:0] my_adder_21_io_i_data_bus_0; // @[FanNetwork.scala 1393:29]
  wire [31:0] my_adder_21_io_i_data_bus_1; // @[FanNetwork.scala 1393:29]
  wire [2:0] my_adder_21_io_i_add_en; // @[FanNetwork.scala 1393:29]
  wire [2:0] my_adder_21_io_i_cmd; // @[FanNetwork.scala 1393:29]
  wire [1:0] my_adder_21_io_o_vn_valid; // @[FanNetwork.scala 1393:29]
  wire [63:0] my_adder_21_io_o_vn; // @[FanNetwork.scala 1393:29]
  wire [31:0] my_adder_21_io_o_adder_0; // @[FanNetwork.scala 1393:29]
  wire [31:0] my_adder_21_io_o_adder_1; // @[FanNetwork.scala 1393:29]
  wire  my_adder_22_clock; // @[FanNetwork.scala 1412:29]
  wire  my_adder_22_reset; // @[FanNetwork.scala 1412:29]
  wire  my_adder_22_io_i_valid; // @[FanNetwork.scala 1412:29]
  wire [31:0] my_adder_22_io_i_data_bus_0; // @[FanNetwork.scala 1412:29]
  wire [31:0] my_adder_22_io_i_data_bus_1; // @[FanNetwork.scala 1412:29]
  wire [2:0] my_adder_22_io_i_add_en; // @[FanNetwork.scala 1412:29]
  wire [2:0] my_adder_22_io_i_cmd; // @[FanNetwork.scala 1412:29]
  wire [1:0] my_adder_22_io_o_vn_valid; // @[FanNetwork.scala 1412:29]
  wire [63:0] my_adder_22_io_o_vn; // @[FanNetwork.scala 1412:29]
  wire [31:0] my_adder_22_io_o_adder_0; // @[FanNetwork.scala 1412:29]
  wire [31:0] my_adder_22_io_o_adder_1; // @[FanNetwork.scala 1412:29]
  wire  my_adder_23_clock; // @[FanNetwork.scala 1430:29]
  wire  my_adder_23_reset; // @[FanNetwork.scala 1430:29]
  wire  my_adder_23_io_i_valid; // @[FanNetwork.scala 1430:29]
  wire [63:0] my_adder_23_io_i_data_bus_0; // @[FanNetwork.scala 1430:29]
  wire [63:0] my_adder_23_io_i_data_bus_1; // @[FanNetwork.scala 1430:29]
  wire [63:0] my_adder_23_io_i_data_bus_2; // @[FanNetwork.scala 1430:29]
  wire [63:0] my_adder_23_io_i_data_bus_3; // @[FanNetwork.scala 1430:29]
  wire [63:0] my_adder_23_io_i_data_bus_4; // @[FanNetwork.scala 1430:29]
  wire [63:0] my_adder_23_io_i_data_bus_5; // @[FanNetwork.scala 1430:29]
  wire [2:0] my_adder_23_io_i_add_en; // @[FanNetwork.scala 1430:29]
  wire [4:0] my_adder_23_io_i_cmd; // @[FanNetwork.scala 1430:29]
  wire [3:0] my_adder_23_io_i_sel; // @[FanNetwork.scala 1430:29]
  wire [63:0] my_adder_23_io_o_vn; // @[FanNetwork.scala 1430:29]
  wire [1:0] my_adder_23_io_o_vn_valid; // @[FanNetwork.scala 1430:29]
  wire [31:0] my_adder_23_io_o_adder; // @[FanNetwork.scala 1430:29]
  wire  my_adder_24_clock; // @[FanNetwork.scala 1447:29]
  wire  my_adder_24_reset; // @[FanNetwork.scala 1447:29]
  wire  my_adder_24_io_i_valid; // @[FanNetwork.scala 1447:29]
  wire [31:0] my_adder_24_io_i_data_bus_0; // @[FanNetwork.scala 1447:29]
  wire [31:0] my_adder_24_io_i_data_bus_1; // @[FanNetwork.scala 1447:29]
  wire [2:0] my_adder_24_io_i_add_en; // @[FanNetwork.scala 1447:29]
  wire [2:0] my_adder_24_io_i_cmd; // @[FanNetwork.scala 1447:29]
  wire [1:0] my_adder_24_io_o_vn_valid; // @[FanNetwork.scala 1447:29]
  wire [63:0] my_adder_24_io_o_vn; // @[FanNetwork.scala 1447:29]
  wire [31:0] my_adder_24_io_o_adder_0; // @[FanNetwork.scala 1447:29]
  wire [31:0] my_adder_24_io_o_adder_1; // @[FanNetwork.scala 1447:29]
  wire  my_adder_25_clock; // @[FanNetwork.scala 1466:29]
  wire  my_adder_25_reset; // @[FanNetwork.scala 1466:29]
  wire  my_adder_25_io_i_valid; // @[FanNetwork.scala 1466:29]
  wire [31:0] my_adder_25_io_i_data_bus_0; // @[FanNetwork.scala 1466:29]
  wire [31:0] my_adder_25_io_i_data_bus_1; // @[FanNetwork.scala 1466:29]
  wire [2:0] my_adder_25_io_i_add_en; // @[FanNetwork.scala 1466:29]
  wire [2:0] my_adder_25_io_i_cmd; // @[FanNetwork.scala 1466:29]
  wire [1:0] my_adder_25_io_o_vn_valid; // @[FanNetwork.scala 1466:29]
  wire [63:0] my_adder_25_io_o_vn; // @[FanNetwork.scala 1466:29]
  wire [31:0] my_adder_25_io_o_adder_0; // @[FanNetwork.scala 1466:29]
  wire [31:0] my_adder_25_io_o_adder_1; // @[FanNetwork.scala 1466:29]
  wire  my_adder_26_clock; // @[FanNetwork.scala 1486:29]
  wire  my_adder_26_reset; // @[FanNetwork.scala 1486:29]
  wire  my_adder_26_io_i_valid; // @[FanNetwork.scala 1486:29]
  wire [31:0] my_adder_26_io_i_data_bus_0; // @[FanNetwork.scala 1486:29]
  wire [31:0] my_adder_26_io_i_data_bus_1; // @[FanNetwork.scala 1486:29]
  wire [2:0] my_adder_26_io_i_add_en; // @[FanNetwork.scala 1486:29]
  wire [2:0] my_adder_26_io_i_cmd; // @[FanNetwork.scala 1486:29]
  wire [1:0] my_adder_26_io_o_vn_valid; // @[FanNetwork.scala 1486:29]
  wire [63:0] my_adder_26_io_o_vn; // @[FanNetwork.scala 1486:29]
  wire [31:0] my_adder_26_io_o_adder_0; // @[FanNetwork.scala 1486:29]
  wire [31:0] my_adder_26_io_o_adder_1; // @[FanNetwork.scala 1486:29]
  wire  my_adder_27_clock; // @[FanNetwork.scala 1504:29]
  wire  my_adder_27_reset; // @[FanNetwork.scala 1504:29]
  wire  my_adder_27_io_i_valid; // @[FanNetwork.scala 1504:29]
  wire [63:0] my_adder_27_io_i_data_bus_0; // @[FanNetwork.scala 1504:29]
  wire [63:0] my_adder_27_io_i_data_bus_1; // @[FanNetwork.scala 1504:29]
  wire [63:0] my_adder_27_io_i_data_bus_2; // @[FanNetwork.scala 1504:29]
  wire [63:0] my_adder_27_io_i_data_bus_3; // @[FanNetwork.scala 1504:29]
  wire [2:0] my_adder_27_io_i_add_en; // @[FanNetwork.scala 1504:29]
  wire [4:0] my_adder_27_io_i_cmd; // @[FanNetwork.scala 1504:29]
  wire [1:0] my_adder_27_io_i_sel; // @[FanNetwork.scala 1504:29]
  wire [63:0] my_adder_27_io_o_vn; // @[FanNetwork.scala 1504:29]
  wire [1:0] my_adder_27_io_o_vn_valid; // @[FanNetwork.scala 1504:29]
  wire [31:0] my_adder_27_io_o_adder; // @[FanNetwork.scala 1504:29]
  wire  my_adder_28_clock; // @[FanNetwork.scala 1525:29]
  wire  my_adder_28_reset; // @[FanNetwork.scala 1525:29]
  wire  my_adder_28_io_i_valid; // @[FanNetwork.scala 1525:29]
  wire [31:0] my_adder_28_io_i_data_bus_0; // @[FanNetwork.scala 1525:29]
  wire [31:0] my_adder_28_io_i_data_bus_1; // @[FanNetwork.scala 1525:29]
  wire [2:0] my_adder_28_io_i_add_en; // @[FanNetwork.scala 1525:29]
  wire [2:0] my_adder_28_io_i_cmd; // @[FanNetwork.scala 1525:29]
  wire [1:0] my_adder_28_io_o_vn_valid; // @[FanNetwork.scala 1525:29]
  wire [63:0] my_adder_28_io_o_vn; // @[FanNetwork.scala 1525:29]
  wire [31:0] my_adder_28_io_o_adder_0; // @[FanNetwork.scala 1525:29]
  wire [31:0] my_adder_28_io_o_adder_1; // @[FanNetwork.scala 1525:29]
  wire  my_adder_29_clock; // @[FanNetwork.scala 1544:29]
  wire  my_adder_29_reset; // @[FanNetwork.scala 1544:29]
  wire  my_adder_29_io_i_valid; // @[FanNetwork.scala 1544:29]
  wire [63:0] my_adder_29_io_i_data_bus_0; // @[FanNetwork.scala 1544:29]
  wire [63:0] my_adder_29_io_i_data_bus_1; // @[FanNetwork.scala 1544:29]
  wire [2:0] my_adder_29_io_i_add_en; // @[FanNetwork.scala 1544:29]
  wire [4:0] my_adder_29_io_i_cmd; // @[FanNetwork.scala 1544:29]
  wire [63:0] my_adder_29_io_o_vn; // @[FanNetwork.scala 1544:29]
  wire [1:0] my_adder_29_io_o_vn_valid; // @[FanNetwork.scala 1544:29]
  wire [31:0] my_adder_29_io_o_adder; // @[FanNetwork.scala 1544:29]
  wire  my_adder_30_clock; // @[FanNetwork.scala 1562:29]
  wire  my_adder_30_reset; // @[FanNetwork.scala 1562:29]
  wire  my_adder_30_io_i_valid; // @[FanNetwork.scala 1562:29]
  wire [63:0] my_adder_30_io_i_data_bus_0; // @[FanNetwork.scala 1562:29]
  wire [63:0] my_adder_30_io_i_data_bus_1; // @[FanNetwork.scala 1562:29]
  wire [2:0] my_adder_30_io_i_add_en; // @[FanNetwork.scala 1562:29]
  wire [4:0] my_adder_30_io_i_cmd; // @[FanNetwork.scala 1562:29]
  wire [63:0] my_adder_30_io_o_vn; // @[FanNetwork.scala 1562:29]
  wire [1:0] my_adder_30_io_o_vn_valid; // @[FanNetwork.scala 1562:29]
  wire [31:0] my_adder_30_io_o_adder; // @[FanNetwork.scala 1562:29]
  reg [31:0] r_fan_ff_lvl_0_to_4_0; // @[FanNetwork.scala 32:38]
  reg [31:0] r_fan_ff_lvl_0_to_4_1; // @[FanNetwork.scala 32:38]
  reg [31:0] r_fan_ff_lvl_0_to_3_0; // @[FanNetwork.scala 33:38]
  reg [31:0] r_fan_ff_lvl_0_to_3_1; // @[FanNetwork.scala 33:38]
  reg [31:0] r_fan_ff_lvl_0_to_3_2; // @[FanNetwork.scala 33:38]
  reg [31:0] r_fan_ff_lvl_0_to_3_3; // @[FanNetwork.scala 33:38]
  reg [31:0] r_fan_ff_lvl_0_to_3_4; // @[FanNetwork.scala 33:38]
  reg [31:0] r_fan_ff_lvl_0_to_3_5; // @[FanNetwork.scala 33:38]
  reg [31:0] r_fan_ff_lvl_0_to_2_0; // @[FanNetwork.scala 34:38]
  reg [31:0] r_fan_ff_lvl_0_to_2_1; // @[FanNetwork.scala 34:38]
  reg [31:0] r_fan_ff_lvl_0_to_2_2; // @[FanNetwork.scala 34:38]
  reg [31:0] r_fan_ff_lvl_0_to_2_3; // @[FanNetwork.scala 34:38]
  reg [31:0] r_fan_ff_lvl_0_to_2_4; // @[FanNetwork.scala 34:38]
  reg [31:0] r_fan_ff_lvl_0_to_2_5; // @[FanNetwork.scala 34:38]
  reg [31:0] r_fan_ff_lvl_0_to_2_6; // @[FanNetwork.scala 34:38]
  reg [31:0] r_fan_ff_lvl_0_to_2_7; // @[FanNetwork.scala 34:38]
  reg [31:0] r_fan_ff_lvl_0_to_2_8; // @[FanNetwork.scala 34:38]
  reg [31:0] r_fan_ff_lvl_0_to_2_9; // @[FanNetwork.scala 34:38]
  reg [31:0] r_fan_ff_lvl_0_to_2_10; // @[FanNetwork.scala 34:38]
  reg [31:0] r_fan_ff_lvl_0_to_2_11; // @[FanNetwork.scala 34:38]
  reg [31:0] r_fan_ff_lvl_0_to_2_12; // @[FanNetwork.scala 34:38]
  reg [31:0] r_fan_ff_lvl_0_to_2_13; // @[FanNetwork.scala 34:38]
  reg [31:0] r_fan_ff_lvl_1_to_4_0; // @[FanNetwork.scala 35:38]
  reg [31:0] r_fan_ff_lvl_1_to_4_1; // @[FanNetwork.scala 35:38]
  reg [31:0] r_fan_ff_lvl_1_to_3_0; // @[FanNetwork.scala 36:38]
  reg [31:0] r_fan_ff_lvl_1_to_3_1; // @[FanNetwork.scala 36:38]
  reg [31:0] r_fan_ff_lvl_1_to_3_2; // @[FanNetwork.scala 36:38]
  reg [31:0] r_fan_ff_lvl_1_to_3_3; // @[FanNetwork.scala 36:38]
  reg [31:0] r_fan_ff_lvl_1_to_3_4; // @[FanNetwork.scala 36:38]
  reg [31:0] r_fan_ff_lvl_1_to_3_5; // @[FanNetwork.scala 36:38]
  reg [31:0] r_fan_ff_lvl_2_to_4_0; // @[FanNetwork.scala 37:38]
  reg [31:0] r_fan_ff_lvl_2_to_4_1; // @[FanNetwork.scala 37:38]
  reg [31:0] r_lvl_output_ff_0; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_1; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_2; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_3; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_6; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_7; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_8; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_9; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_10; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_11; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_12; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_13; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_14; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_15; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_16; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_17; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_18; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_19; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_20; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_21; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_22; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_23; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_24; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_25; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_26; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_27; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_28; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_29; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_30; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_31; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_32; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_33; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_34; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_35; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_37; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_38; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_39; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_40; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_41; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_42; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_43; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_44; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_45; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_46; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_47; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_48; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_49; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_50; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_51; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_52; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_53; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_54; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_55; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_56; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_57; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_58; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_59; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_60; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_61; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_62; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_63; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_64; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_65; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_66; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_67; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_68; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_69; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_70; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_71; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_72; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_73; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_74; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_75; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_76; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_77; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_78; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_79; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_80; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_81; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_82; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_83; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_84; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_85; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_86; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_87; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_88; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_89; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_90; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_91; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_92; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_93; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_94; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_95; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_96; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_97; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_98; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_99; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_100; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_101; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_102; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_103; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_104; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_105; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_106; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_107; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_108; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_109; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_110; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_112; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_113; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_114; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_115; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_116; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_117; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_118; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_119; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_120; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_121; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_122; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_123; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_124; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_125; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_126; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_127; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_128; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_129; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_130; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_131; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_132; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_133; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_134; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_135; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_136; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_137; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_138; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_139; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_140; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_141; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_142; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_143; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_144; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_145; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_146; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_147; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_148; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_149; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_150; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_151; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_152; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_153; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_154; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_155; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_156; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_157; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_158; // @[FanNetwork.scala 50:34]
  reg [31:0] r_lvl_output_ff_159; // @[FanNetwork.scala 50:34]
  reg  r_lvl_output_ff_valid_0; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_1; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_2; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_3; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_4; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_5; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_6; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_7; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_8; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_9; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_10; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_11; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_12; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_13; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_14; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_15; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_16; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_17; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_18; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_19; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_20; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_21; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_22; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_23; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_24; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_25; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_26; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_27; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_28; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_29; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_30; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_31; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_32; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_33; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_34; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_35; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_36; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_37; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_38; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_39; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_40; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_41; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_42; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_43; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_44; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_45; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_46; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_47; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_48; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_49; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_50; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_51; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_52; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_53; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_54; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_55; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_56; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_57; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_58; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_59; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_60; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_61; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_62; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_63; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_64; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_65; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_66; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_67; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_68; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_69; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_70; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_71; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_72; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_73; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_74; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_75; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_76; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_77; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_78; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_79; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_80; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_81; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_82; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_83; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_84; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_85; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_86; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_87; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_88; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_89; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_90; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_91; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_92; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_93; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_94; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_95; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_96; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_97; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_98; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_99; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_100; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_101; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_102; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_103; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_104; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_105; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_106; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_107; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_108; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_109; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_110; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_111; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_112; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_113; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_114; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_115; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_116; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_117; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_118; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_119; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_120; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_121; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_122; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_123; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_124; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_125; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_126; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_127; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_128; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_129; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_130; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_131; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_132; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_133; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_134; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_135; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_136; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_137; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_138; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_139; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_140; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_141; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_142; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_143; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_144; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_145; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_146; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_147; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_148; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_149; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_150; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_151; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_152; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_153; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_154; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_155; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_156; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_157; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_158; // @[FanNetwork.scala 51:40]
  reg  r_lvl_output_ff_valid_159; // @[FanNetwork.scala 51:40]
  reg  r_valid_0; // @[FanNetwork.scala 52:26]
  reg  r_valid_1; // @[FanNetwork.scala 52:26]
  reg  r_valid_2; // @[FanNetwork.scala 52:26]
  reg  r_valid_3; // @[FanNetwork.scala 52:26]
  reg  r_valid_4; // @[FanNetwork.scala 52:26]
  reg [31:0] r_final_sum; // @[FanNetwork.scala 54:30]
  reg  r_final_add; // @[FanNetwork.scala 55:30]
  reg  r_final_add2; // @[FanNetwork.scala 56:31]
  wire  w_vn_lvl_0_valid_1 = my_adder_0_io_o_vn_valid[1]; // @[FanNetwork.scala 1028:52]
  wire  w_vn_lvl_0_valid_0 = my_adder_0_io_o_vn_valid[0]; // @[FanNetwork.scala 1027:52]
  wire  _T_9 = w_vn_lvl_0_valid_1 & ~w_vn_lvl_0_valid_0; // @[FanNetwork.scala 88:48]
  wire  _T_14 = ~w_vn_lvl_0_valid_1 & w_vn_lvl_0_valid_0; // @[FanNetwork.scala 93:48]
  wire [31:0] w_vn_lvl_0_0 = my_adder_0_io_o_vn[31:0]; // @[FanNetwork.scala 1025:40]
  wire [31:0] w_vn_lvl_0_1 = my_adder_0_io_o_vn[63:32]; // @[FanNetwork.scala 1026:40]
  wire  _GEN_6 = w_vn_lvl_0_valid_1 & ~w_vn_lvl_0_valid_0 ? 1'h0 : _T_14; // @[FanNetwork.scala 88:83 92:30]
  wire  _GEN_9 = w_vn_lvl_0_valid_1 & w_vn_lvl_0_valid_0 | _T_9; // @[FanNetwork.scala 83:77 86:30]
  wire  _GEN_10 = w_vn_lvl_0_valid_1 & w_vn_lvl_0_valid_0 | _GEN_6; // @[FanNetwork.scala 83:77 87:30]
  wire  w_vn_lvl_0_valid_3 = my_adder_2_io_o_vn_valid[1]; // @[FanNetwork.scala 1058:52]
  wire  w_vn_lvl_0_valid_2 = my_adder_2_io_o_vn_valid[0]; // @[FanNetwork.scala 1057:52]
  wire  _T_24 = w_vn_lvl_0_valid_3 & ~w_vn_lvl_0_valid_2; // @[FanNetwork.scala 111:48]
  wire  _T_29 = ~w_vn_lvl_0_valid_3 & w_vn_lvl_0_valid_2; // @[FanNetwork.scala 116:48]
  wire [31:0] w_vn_lvl_0_2 = my_adder_4_io_o_vn[31:0]; // @[FanNetwork.scala 1089:40]
  wire [31:0] w_vn_lvl_0_3 = my_adder_4_io_o_vn[63:32]; // @[FanNetwork.scala 1090:40]
  wire  _GEN_17 = w_vn_lvl_0_valid_3 & ~w_vn_lvl_0_valid_2 ? 1'h0 : _T_29; // @[FanNetwork.scala 111:83 115:30]
  wire  _GEN_20 = w_vn_lvl_0_valid_3 & w_vn_lvl_0_valid_2 | _T_24; // @[FanNetwork.scala 106:77 109:30]
  wire  _GEN_21 = w_vn_lvl_0_valid_3 & w_vn_lvl_0_valid_2 | _GEN_17; // @[FanNetwork.scala 106:77 110:30]
  wire  w_vn_lvl_0_valid_5 = my_adder_4_io_o_vn_valid[1]; // @[FanNetwork.scala 1093:52]
  wire  w_vn_lvl_0_valid_4 = my_adder_4_io_o_vn_valid[0]; // @[FanNetwork.scala 1092:52]
  wire  _T_39 = w_vn_lvl_0_valid_5 & ~w_vn_lvl_0_valid_4; // @[FanNetwork.scala 133:48]
  wire  _T_44 = ~w_vn_lvl_0_valid_5 & w_vn_lvl_0_valid_4; // @[FanNetwork.scala 138:48]
  wire  _GEN_28 = w_vn_lvl_0_valid_5 & ~w_vn_lvl_0_valid_4 ? 1'h0 : _T_44; // @[FanNetwork.scala 133:83 137:30]
  wire  _GEN_31 = w_vn_lvl_0_valid_5 & w_vn_lvl_0_valid_4 | _T_39; // @[FanNetwork.scala 128:77 131:30]
  wire  _GEN_32 = w_vn_lvl_0_valid_5 & w_vn_lvl_0_valid_4 | _GEN_28; // @[FanNetwork.scala 128:77 132:30]
  wire  w_vn_lvl_0_valid_7 = my_adder_6_io_o_vn_valid[1]; // @[FanNetwork.scala 1128:52]
  wire  w_vn_lvl_0_valid_6 = my_adder_6_io_o_vn_valid[0]; // @[FanNetwork.scala 1127:52]
  wire  _T_54 = w_vn_lvl_0_valid_7 & ~w_vn_lvl_0_valid_6; // @[FanNetwork.scala 156:48]
  wire  _T_59 = ~w_vn_lvl_0_valid_7 & w_vn_lvl_0_valid_6; // @[FanNetwork.scala 161:48]
  wire [31:0] w_vn_lvl_0_6 = my_adder_6_io_o_vn[31:0]; // @[FanNetwork.scala 1124:40]
  wire [31:0] w_vn_lvl_0_7 = my_adder_6_io_o_vn[63:32]; // @[FanNetwork.scala 1125:40]
  wire  _GEN_39 = w_vn_lvl_0_valid_7 & ~w_vn_lvl_0_valid_6 ? 1'h0 : _T_59; // @[FanNetwork.scala 156:83 160:30]
  wire  _GEN_42 = w_vn_lvl_0_valid_7 & w_vn_lvl_0_valid_6 | _T_54; // @[FanNetwork.scala 151:77 154:30]
  wire  _GEN_43 = w_vn_lvl_0_valid_7 & w_vn_lvl_0_valid_6 | _GEN_39; // @[FanNetwork.scala 151:77 155:30]
  wire  w_vn_lvl_0_valid_9 = my_adder_8_io_o_vn_valid[0]; // @[FanNetwork.scala 1164:52]
  wire  w_vn_lvl_0_valid_8 = my_adder_8_io_o_vn_valid[1]; // @[FanNetwork.scala 1163:52]
  wire  _T_66 = w_vn_lvl_0_valid_9 & ~w_vn_lvl_0_valid_8; // @[FanNetwork.scala 179:40]
  wire  _T_70 = ~w_vn_lvl_0_valid_9 & w_vn_lvl_0_valid_8; // @[FanNetwork.scala 184:41]
  wire [31:0] w_vn_lvl_0_8 = my_adder_8_io_o_vn[31:0]; // @[FanNetwork.scala 1160:40]
  wire [31:0] w_vn_lvl_0_9 = my_adder_8_io_o_vn[63:32]; // @[FanNetwork.scala 1161:40]
  wire  _GEN_50 = w_vn_lvl_0_valid_9 & ~w_vn_lvl_0_valid_8 ? 1'h0 : _T_70; // @[FanNetwork.scala 179:68 183:30]
  wire  _GEN_53 = w_vn_lvl_0_valid_9 & w_vn_lvl_0_valid_8 | _T_66; // @[FanNetwork.scala 174:61 177:30]
  wire  _GEN_54 = w_vn_lvl_0_valid_9 & w_vn_lvl_0_valid_8 | _GEN_50; // @[FanNetwork.scala 174:61 178:30]
  wire  w_vn_lvl_0_valid_11 = my_adder_10_io_o_vn_valid[1]; // @[FanNetwork.scala 1198:58]
  wire  w_vn_lvl_0_valid_10 = my_adder_10_io_o_vn_valid[0]; // @[FanNetwork.scala 1197:54]
  wire  _T_77 = w_vn_lvl_0_valid_11 & ~w_vn_lvl_0_valid_10; // @[FanNetwork.scala 202:41]
  wire  _T_81 = ~w_vn_lvl_0_valid_11 & w_vn_lvl_0_valid_10; // @[FanNetwork.scala 207:42]
  wire [31:0] w_vn_lvl_0_10 = my_adder_10_io_o_vn[31:0]; // @[FanNetwork.scala 1194:42]
  wire  _GEN_61 = w_vn_lvl_0_valid_11 & ~w_vn_lvl_0_valid_10 ? 1'h0 : _T_81; // @[FanNetwork.scala 202:70 206:31]
  wire  _GEN_64 = w_vn_lvl_0_valid_11 & w_vn_lvl_0_valid_10 | _T_77; // @[FanNetwork.scala 197:63 200:31]
  wire  _GEN_65 = w_vn_lvl_0_valid_11 & w_vn_lvl_0_valid_10 | _GEN_61; // @[FanNetwork.scala 197:63 201:31]
  wire  w_vn_lvl_0_valid_13 = my_adder_12_io_o_vn_valid[1]; // @[FanNetwork.scala 1237:58]
  wire  w_vn_lvl_0_valid_12 = my_adder_12_io_o_vn_valid[0]; // @[FanNetwork.scala 1236:54]
  wire  _T_88 = w_vn_lvl_0_valid_13 & ~w_vn_lvl_0_valid_12; // @[FanNetwork.scala 225:41]
  wire  _T_92 = ~w_vn_lvl_0_valid_13 & w_vn_lvl_0_valid_12; // @[FanNetwork.scala 230:42]
  wire [31:0] w_vn_lvl_0_12 = my_adder_12_io_o_vn[31:0]; // @[FanNetwork.scala 1233:42]
  wire [31:0] w_vn_lvl_0_13 = my_adder_12_io_o_vn[63:32]; // @[FanNetwork.scala 1234:46]
  wire  _GEN_72 = w_vn_lvl_0_valid_13 & ~w_vn_lvl_0_valid_12 ? 1'h0 : _T_92; // @[FanNetwork.scala 225:70 229:31]
  wire  _GEN_75 = w_vn_lvl_0_valid_13 & w_vn_lvl_0_valid_12 | _T_88; // @[FanNetwork.scala 220:63 223:31]
  wire  _GEN_76 = w_vn_lvl_0_valid_13 & w_vn_lvl_0_valid_12 | _GEN_72; // @[FanNetwork.scala 220:63 224:31]
  wire  w_vn_lvl_0_valid_15 = my_adder_14_io_o_vn_valid[1]; // @[FanNetwork.scala 1273:54]
  wire  w_vn_lvl_0_valid_14 = my_adder_14_io_o_vn_valid[0]; // @[FanNetwork.scala 1272:54]
  wire  _T_99 = w_vn_lvl_0_valid_15 & ~w_vn_lvl_0_valid_14; // @[FanNetwork.scala 248:41]
  wire  _T_103 = ~w_vn_lvl_0_valid_15 & w_vn_lvl_0_valid_14; // @[FanNetwork.scala 253:42]
  wire [31:0] w_vn_lvl_0_14 = my_adder_14_io_o_vn[31:0]; // @[FanNetwork.scala 1269:42]
  wire [31:0] w_vn_lvl_0_15 = my_adder_14_io_o_vn[63:32]; // @[FanNetwork.scala 1270:42]
  wire  _GEN_83 = w_vn_lvl_0_valid_15 & ~w_vn_lvl_0_valid_14 ? 1'h0 : _T_103; // @[FanNetwork.scala 248:70 252:31]
  wire  _GEN_86 = w_vn_lvl_0_valid_15 & w_vn_lvl_0_valid_14 | _T_99; // @[FanNetwork.scala 243:63 246:31]
  wire  _GEN_87 = w_vn_lvl_0_valid_15 & w_vn_lvl_0_valid_14 | _GEN_83; // @[FanNetwork.scala 243:63 247:31]
  wire  w_vn_lvl_0_valid_17 = my_adder_16_io_o_vn_valid[1]; // @[FanNetwork.scala 1311:54]
  wire  w_vn_lvl_0_valid_16 = my_adder_16_io_o_vn_valid[0]; // @[FanNetwork.scala 1310:54]
  wire  _T_110 = w_vn_lvl_0_valid_17 & ~w_vn_lvl_0_valid_16; // @[FanNetwork.scala 271:41]
  wire  _T_114 = ~w_vn_lvl_0_valid_17 & w_vn_lvl_0_valid_16; // @[FanNetwork.scala 276:42]
  wire [31:0] w_vn_lvl_0_16 = my_adder_16_io_o_vn[31:0]; // @[FanNetwork.scala 1307:42]
  wire [31:0] w_vn_lvl_0_17 = my_adder_16_io_o_vn[63:32]; // @[FanNetwork.scala 1308:42]
  wire  _GEN_94 = w_vn_lvl_0_valid_17 & ~w_vn_lvl_0_valid_16 ? 1'h0 : _T_114; // @[FanNetwork.scala 271:70 275:31]
  wire  _GEN_97 = w_vn_lvl_0_valid_17 & w_vn_lvl_0_valid_16 | _T_110; // @[FanNetwork.scala 266:63 269:31]
  wire  _GEN_98 = w_vn_lvl_0_valid_17 & w_vn_lvl_0_valid_16 | _GEN_94; // @[FanNetwork.scala 266:63 270:31]
  wire  w_vn_lvl_0_valid_19 = my_adder_18_io_o_vn_valid[1]; // @[FanNetwork.scala 1347:54]
  wire  w_vn_lvl_0_valid_18 = my_adder_18_io_o_vn_valid[0]; // @[FanNetwork.scala 1346:54]
  wire  _T_121 = w_vn_lvl_0_valid_19 & ~w_vn_lvl_0_valid_18; // @[FanNetwork.scala 294:41]
  wire  _T_125 = ~w_vn_lvl_0_valid_19 & w_vn_lvl_0_valid_18; // @[FanNetwork.scala 299:42]
  wire [31:0] w_vn_lvl_0_18 = my_adder_18_io_o_vn[31:0]; // @[FanNetwork.scala 1343:42]
  wire [31:0] w_vn_lvl_0_19 = my_adder_18_io_o_vn[63:32]; // @[FanNetwork.scala 1344:42]
  wire  _GEN_105 = w_vn_lvl_0_valid_19 & ~w_vn_lvl_0_valid_18 ? 1'h0 : _T_125; // @[FanNetwork.scala 294:70 298:31]
  wire  _GEN_108 = w_vn_lvl_0_valid_19 & w_vn_lvl_0_valid_18 | _T_121; // @[FanNetwork.scala 289:63 292:31]
  wire  _GEN_109 = w_vn_lvl_0_valid_19 & w_vn_lvl_0_valid_18 | _GEN_105; // @[FanNetwork.scala 289:63 293:31]
  wire  w_vn_lvl_0_valid_21 = my_adder_20_io_o_vn_valid[1]; // @[FanNetwork.scala 1385:54]
  wire  w_vn_lvl_0_valid_20 = my_adder_20_io_o_vn_valid[0]; // @[FanNetwork.scala 1384:54]
  wire  _T_132 = w_vn_lvl_0_valid_21 & ~w_vn_lvl_0_valid_20; // @[FanNetwork.scala 317:41]
  wire  _T_136 = ~w_vn_lvl_0_valid_21 & w_vn_lvl_0_valid_20; // @[FanNetwork.scala 322:42]
  wire [31:0] w_vn_lvl_0_20 = my_adder_20_io_o_vn[31:0]; // @[FanNetwork.scala 1381:42]
  wire [31:0] w_vn_lvl_0_21 = my_adder_20_io_o_vn[63:32]; // @[FanNetwork.scala 1382:42]
  wire  _GEN_116 = w_vn_lvl_0_valid_21 & ~w_vn_lvl_0_valid_20 ? 1'h0 : _T_136; // @[FanNetwork.scala 317:70 321:31]
  wire  _GEN_119 = w_vn_lvl_0_valid_21 & w_vn_lvl_0_valid_20 | _T_132; // @[FanNetwork.scala 312:63 315:31]
  wire  _GEN_120 = w_vn_lvl_0_valid_21 & w_vn_lvl_0_valid_20 | _GEN_116; // @[FanNetwork.scala 312:63 316:31]
  wire  w_vn_lvl_0_valid_23 = my_adder_22_io_o_vn_valid[1]; // @[FanNetwork.scala 1424:54]
  wire  w_vn_lvl_0_valid_22 = my_adder_22_io_o_vn_valid[0]; // @[FanNetwork.scala 1423:54]
  wire  _T_143 = w_vn_lvl_0_valid_23 & ~w_vn_lvl_0_valid_22; // @[FanNetwork.scala 340:41]
  wire  _T_147 = ~w_vn_lvl_0_valid_23 & w_vn_lvl_0_valid_22; // @[FanNetwork.scala 345:42]
  wire [31:0] w_vn_lvl_0_22 = my_adder_22_io_o_vn[31:0]; // @[FanNetwork.scala 1420:42]
  wire [31:0] w_vn_lvl_0_23 = my_adder_22_io_o_vn[63:32]; // @[FanNetwork.scala 1421:42]
  wire  _GEN_127 = w_vn_lvl_0_valid_23 & ~w_vn_lvl_0_valid_22 ? 1'h0 : _T_147; // @[FanNetwork.scala 340:70 344:31]
  wire  _GEN_130 = w_vn_lvl_0_valid_23 & w_vn_lvl_0_valid_22 | _T_143; // @[FanNetwork.scala 335:63 338:31]
  wire  _GEN_131 = w_vn_lvl_0_valid_23 & w_vn_lvl_0_valid_22 | _GEN_127; // @[FanNetwork.scala 335:63 339:31]
  wire  w_vn_lvl_0_valid_25 = my_adder_24_io_o_vn_valid[1]; // @[FanNetwork.scala 1459:54]
  wire  w_vn_lvl_0_valid_24 = my_adder_24_io_o_vn_valid[0]; // @[FanNetwork.scala 1458:54]
  wire  _T_154 = w_vn_lvl_0_valid_25 & ~w_vn_lvl_0_valid_24; // @[FanNetwork.scala 363:41]
  wire  _T_158 = ~w_vn_lvl_0_valid_25 & w_vn_lvl_0_valid_24; // @[FanNetwork.scala 368:42]
  wire [31:0] w_vn_lvl_0_24 = my_adder_24_io_o_vn[31:0]; // @[FanNetwork.scala 1455:42]
  wire [31:0] w_vn_lvl_0_25 = my_adder_24_io_o_vn[63:32]; // @[FanNetwork.scala 1456:42]
  wire  _GEN_138 = w_vn_lvl_0_valid_25 & ~w_vn_lvl_0_valid_24 ? 1'h0 : _T_158; // @[FanNetwork.scala 363:70 367:31]
  wire  _GEN_141 = w_vn_lvl_0_valid_25 & w_vn_lvl_0_valid_24 | _T_154; // @[FanNetwork.scala 358:63 361:31]
  wire  _GEN_142 = w_vn_lvl_0_valid_25 & w_vn_lvl_0_valid_24 | _GEN_138; // @[FanNetwork.scala 358:63 362:31]
  wire  w_vn_lvl_0_valid_27 = my_adder_26_io_o_vn_valid[1]; // @[FanNetwork.scala 1498:54]
  wire  w_vn_lvl_0_valid_26 = my_adder_26_io_o_vn_valid[0]; // @[FanNetwork.scala 1497:54]
  wire  _T_165 = w_vn_lvl_0_valid_27 & ~w_vn_lvl_0_valid_26; // @[FanNetwork.scala 386:41]
  wire  _T_169 = ~w_vn_lvl_0_valid_27 & w_vn_lvl_0_valid_26; // @[FanNetwork.scala 391:42]
  wire [31:0] w_vn_lvl_0_26 = my_adder_26_io_o_vn[31:0]; // @[FanNetwork.scala 1494:42]
  wire [31:0] w_vn_lvl_0_27 = my_adder_26_io_o_vn[63:32]; // @[FanNetwork.scala 1495:42]
  wire  _GEN_149 = w_vn_lvl_0_valid_27 & ~w_vn_lvl_0_valid_26 ? 1'h0 : _T_169; // @[FanNetwork.scala 386:70 390:31]
  wire  _GEN_152 = w_vn_lvl_0_valid_27 & w_vn_lvl_0_valid_26 | _T_165; // @[FanNetwork.scala 381:63 384:31]
  wire  _GEN_153 = w_vn_lvl_0_valid_27 & w_vn_lvl_0_valid_26 | _GEN_149; // @[FanNetwork.scala 381:63 385:31]
  wire  w_vn_lvl_0_valid_29 = my_adder_28_io_o_vn_valid[1]; // @[FanNetwork.scala 1537:54]
  wire  w_vn_lvl_0_valid_28 = my_adder_28_io_o_vn_valid[0]; // @[FanNetwork.scala 1536:54]
  wire  _T_176 = w_vn_lvl_0_valid_29 & ~w_vn_lvl_0_valid_28; // @[FanNetwork.scala 409:41]
  wire  _T_180 = ~w_vn_lvl_0_valid_29 & w_vn_lvl_0_valid_28; // @[FanNetwork.scala 414:42]
  wire [31:0] w_vn_lvl_0_28 = my_adder_28_io_o_vn[31:0]; // @[FanNetwork.scala 1533:42]
  wire [31:0] w_vn_lvl_0_29 = my_adder_28_io_o_vn[63:32]; // @[FanNetwork.scala 1534:46]
  wire  _GEN_160 = w_vn_lvl_0_valid_29 & ~w_vn_lvl_0_valid_28 ? 1'h0 : _T_180; // @[FanNetwork.scala 409:70 413:31]
  wire  _GEN_163 = w_vn_lvl_0_valid_29 & w_vn_lvl_0_valid_28 | _T_176; // @[FanNetwork.scala 404:63 407:31]
  wire  _GEN_164 = w_vn_lvl_0_valid_29 & w_vn_lvl_0_valid_28 | _GEN_160; // @[FanNetwork.scala 404:63 408:31]
  wire  w_vn_lvl_0_valid_31 = my_adder_30_io_o_vn_valid[1]; // @[FanNetwork.scala 1574:54]
  wire  w_vn_lvl_0_valid_30 = my_adder_30_io_o_vn_valid[0]; // @[FanNetwork.scala 1573:54]
  wire  _T_187 = w_vn_lvl_0_valid_31 & ~w_vn_lvl_0_valid_30; // @[FanNetwork.scala 432:40]
  wire  _T_191 = ~w_vn_lvl_0_valid_31 & w_vn_lvl_0_valid_30; // @[FanNetwork.scala 437:41]
  wire [31:0] w_vn_lvl_0_30 = my_adder_30_io_o_vn[31:0]; // @[FanNetwork.scala 1570:42]
  wire [31:0] w_vn_lvl_0_31 = my_adder_30_io_o_vn[63:32]; // @[FanNetwork.scala 1571:42]
  wire  _GEN_171 = w_vn_lvl_0_valid_31 & ~w_vn_lvl_0_valid_30 ? 1'h0 : _T_191; // @[FanNetwork.scala 432:69 436:31]
  wire  _GEN_174 = w_vn_lvl_0_valid_31 & w_vn_lvl_0_valid_30 | _T_187; // @[FanNetwork.scala 427:62 430:31]
  wire  _GEN_175 = w_vn_lvl_0_valid_31 & w_vn_lvl_0_valid_30 | _GEN_171; // @[FanNetwork.scala 427:62 431:31]
  wire  w_vn_lvl_1_valid_0 = my_adder_1_io_o_vn_valid[0]; // @[FanNetwork.scala 1041:52]
  wire [31:0] w_vn_lvl_1_0 = my_adder_1_io_o_vn[31:0]; // @[FanNetwork.scala 1039:40]
  wire  _GEN_177 = w_vn_lvl_1_valid_0 | r_lvl_output_ff_valid_1; // @[FanNetwork.scala 455:34 457:35 460:35]
  wire  w_vn_lvl_1_valid_1 = my_adder_1_io_o_vn_valid[1]; // @[FanNetwork.scala 1042:52]
  wire [31:0] w_vn_lvl_1_1 = my_adder_1_io_o_vn[63:32]; // @[FanNetwork.scala 1040:40]
  wire  _GEN_179 = w_vn_lvl_1_valid_1 | r_lvl_output_ff_valid_2; // @[FanNetwork.scala 463:34 465:35 468:35]
  wire  w_vn_lvl_1_valid_2 = my_adder_5_io_o_vn_valid[0]; // @[FanNetwork.scala 1110:52]
  wire [31:0] w_vn_lvl_1_2 = my_adder_5_io_o_vn[31:0]; // @[FanNetwork.scala 1107:40]
  wire  _GEN_181 = w_vn_lvl_1_valid_2 | r_lvl_output_ff_valid_5; // @[FanNetwork.scala 477:34 479:35 482:35]
  wire  w_vn_lvl_1_valid_3 = my_adder_5_io_o_vn_valid[1]; // @[FanNetwork.scala 1111:52]
  wire [31:0] w_vn_lvl_1_3 = my_adder_5_io_o_vn[63:32]; // @[FanNetwork.scala 1108:40]
  wire  _GEN_183 = w_vn_lvl_1_valid_3 | r_lvl_output_ff_valid_6; // @[FanNetwork.scala 485:34 487:35 490:35]
  wire  w_vn_lvl_1_valid_4 = my_adder_9_io_o_vn_valid[0]; // @[FanNetwork.scala 1180:52]
  wire [31:0] w_vn_lvl_1_4 = my_adder_9_io_o_vn[31:0]; // @[FanNetwork.scala 1177:40]
  wire  _GEN_185 = w_vn_lvl_1_valid_4 | r_lvl_output_ff_valid_9; // @[FanNetwork.scala 501:34 503:35 506:35]
  wire  w_vn_lvl_1_valid_5 = my_adder_9_io_o_vn_valid[1]; // @[FanNetwork.scala 1181:56]
  wire [31:0] w_vn_lvl_1_5 = my_adder_9_io_o_vn[63:32]; // @[FanNetwork.scala 1178:44]
  wire  _GEN_187 = w_vn_lvl_1_valid_5 | r_lvl_output_ff_valid_10; // @[FanNetwork.scala 508:34 510:35 513:35]
  wire  w_vn_lvl_1_valid_6 = my_adder_13_io_o_vn_valid[0]; // @[FanNetwork.scala 1254:53]
  wire [31:0] w_vn_lvl_1_6 = my_adder_13_io_o_vn[31:0]; // @[FanNetwork.scala 1251:41]
  wire  _GEN_189 = w_vn_lvl_1_valid_6 | r_lvl_output_ff_valid_13; // @[FanNetwork.scala 522:34 524:35 527:35]
  wire  w_vn_lvl_1_valid_7 = my_adder_13_io_o_vn_valid[1]; // @[FanNetwork.scala 1255:57]
  wire [31:0] w_vn_lvl_1_7 = my_adder_13_io_o_vn[63:32]; // @[FanNetwork.scala 1252:45]
  wire  _GEN_191 = w_vn_lvl_1_valid_7 | r_lvl_output_ff_valid_14; // @[FanNetwork.scala 530:34 532:35 535:35]
  wire  w_vn_lvl_1_valid_8 = my_adder_17_io_o_vn_valid[0]; // @[FanNetwork.scala 1328:53]
  wire [31:0] w_vn_lvl_1_8 = my_adder_17_io_o_vn[31:0]; // @[FanNetwork.scala 1325:41]
  wire  _GEN_193 = w_vn_lvl_1_valid_8 | r_lvl_output_ff_valid_17; // @[FanNetwork.scala 543:34 545:35 548:35]
  wire  w_vn_lvl_1_valid_9 = my_adder_17_io_o_vn_valid[1]; // @[FanNetwork.scala 1329:53]
  wire [31:0] w_vn_lvl_1_9 = my_adder_17_io_o_vn[63:32]; // @[FanNetwork.scala 1326:41]
  wire  _GEN_195 = w_vn_lvl_1_valid_9 | r_lvl_output_ff_valid_18; // @[FanNetwork.scala 551:34 553:35 556:35]
  wire  w_vn_lvl_1_valid_10 = my_adder_21_io_o_vn_valid[0]; // @[FanNetwork.scala 1405:54]
  wire [31:0] w_vn_lvl_1_10 = my_adder_21_io_o_vn[31:0]; // @[FanNetwork.scala 1402:42]
  wire  _GEN_197 = w_vn_lvl_1_valid_10 | r_lvl_output_ff_valid_21; // @[FanNetwork.scala 567:35 569:35 572:35]
  wire  w_vn_lvl_1_valid_11 = my_adder_21_io_o_vn_valid[1]; // @[FanNetwork.scala 1406:54]
  wire [31:0] w_vn_lvl_1_11 = my_adder_21_io_o_vn[63:32]; // @[FanNetwork.scala 1403:42]
  wire  _GEN_199 = w_vn_lvl_1_valid_11 | r_lvl_output_ff_valid_22; // @[FanNetwork.scala 575:35 577:35 580:35]
  wire  w_vn_lvl_1_valid_12 = my_adder_25_io_o_vn_valid[0]; // @[FanNetwork.scala 1477:54]
  wire [31:0] w_vn_lvl_1_12 = my_adder_25_io_o_vn[31:0];
  wire  _GEN_201 = w_vn_lvl_1_valid_12 | r_lvl_output_ff_valid_25; // @[FanNetwork.scala 589:35 591:35 594:35]
  wire  w_vn_lvl_1_valid_13 = my_adder_25_io_o_vn_valid[1]; // @[FanNetwork.scala 1478:54]
  wire [31:0] w_vn_lvl_1_13 = my_adder_25_io_o_vn[63:32]; // @[FanNetwork.scala 1475:42]
  wire  _GEN_203 = w_vn_lvl_1_valid_13 | r_lvl_output_ff_valid_26; // @[FanNetwork.scala 597:35 599:35 602:35]
  wire  w_vn_lvl_1_valid_14 = my_adder_29_io_o_vn_valid[0]; // @[FanNetwork.scala 1555:54]
  wire [31:0] w_vn_lvl_1_14 = my_adder_29_io_o_vn[31:0]; // @[FanNetwork.scala 1552:42]
  wire  _GEN_205 = w_vn_lvl_1_valid_14 | r_lvl_output_ff_valid_29; // @[FanNetwork.scala 611:43 613:35 616:31]
  wire  w_vn_lvl_1_valid_15 = my_adder_29_io_o_vn_valid[1]; // @[FanNetwork.scala 1556:54]
  wire [31:0] w_vn_lvl_1_15 = my_adder_29_io_o_vn[63:32]; // @[FanNetwork.scala 1553:42]
  wire  _GEN_207 = w_vn_lvl_1_valid_15 | r_lvl_output_ff_valid_30; // @[FanNetwork.scala 619:43 621:35 624:35]
  wire  w_vn_lvl_2_valid_0 = my_adder_3_io_o_vn_valid[0]; // @[FanNetwork.scala 1076:52]
  wire [31:0] w_vn_lvl_2_0 = my_adder_3_io_o_vn[31:0]; // @[FanNetwork.scala 1073:40]
  wire  _GEN_209 = w_vn_lvl_2_valid_0 | r_lvl_output_ff_valid_35; // @[FanNetwork.scala 645:43 647:35 650:39]
  wire  w_vn_lvl_2_valid_1 = my_adder_3_io_o_vn_valid[1]; // @[FanNetwork.scala 1077:52]
  wire [31:0] w_vn_lvl_2_1 = my_adder_3_io_o_vn[63:32]; // @[FanNetwork.scala 1074:40]
  wire  _GEN_211 = w_vn_lvl_2_valid_1 | r_lvl_output_ff_valid_36; // @[FanNetwork.scala 653:43 655:35 658:35]
  wire  w_vn_lvl_2_valid_2 = my_adder_11_io_o_vn_valid[0]; // @[FanNetwork.scala 1218:53]
  wire [31:0] w_vn_lvl_2_2 = my_adder_11_io_o_vn[31:0]; // @[FanNetwork.scala 1215:41]
  wire  _GEN_213 = w_vn_lvl_2_valid_2 | r_lvl_output_ff_valid_43; // @[FanNetwork.scala 679:43 681:35 684:35]
  wire  w_vn_lvl_2_valid_3 = my_adder_11_io_o_vn_valid[1]; // @[FanNetwork.scala 1219:57]
  wire [31:0] w_vn_lvl_2_3 = my_adder_11_io_o_vn[63:32]; // @[FanNetwork.scala 1216:45]
  wire  _GEN_215 = w_vn_lvl_2_valid_3 | r_lvl_output_ff_valid_44; // @[FanNetwork.scala 687:43 689:35 692:35]
  wire  w_vn_lvl_2_valid_4 = my_adder_19_io_o_vn_valid[0]; // @[FanNetwork.scala 1365:53]
  wire [31:0] w_vn_lvl_2_4 = my_adder_19_io_o_vn[31:0]; // @[FanNetwork.scala 1362:41]
  wire  _GEN_217 = w_vn_lvl_2_valid_4 | r_lvl_output_ff_valid_51; // @[FanNetwork.scala 713:43 715:35 718:35]
  wire  w_vn_lvl_2_valid_5 = my_adder_19_io_o_vn_valid[1]; // @[FanNetwork.scala 1366:53]
  wire [31:0] w_vn_lvl_2_5 = my_adder_19_io_o_vn[63:32]; // @[FanNetwork.scala 1363:41]
  wire  _GEN_219 = w_vn_lvl_2_valid_5 | r_lvl_output_ff_valid_52; // @[FanNetwork.scala 721:40 723:35 726:31]
  wire  w_vn_lvl_2_valid_6 = my_adder_27_io_o_vn_valid[0]; // @[FanNetwork.scala 1516:53]
  wire [31:0] w_vn_lvl_2_6 = my_adder_27_io_o_vn[31:0]; // @[FanNetwork.scala 1513:41]
  wire  _GEN_221 = w_vn_lvl_2_valid_6 | r_lvl_output_ff_valid_59; // @[FanNetwork.scala 747:40 749:35 752:35]
  wire  w_vn_lvl_2_valid_7 = my_adder_27_io_o_vn_valid[1]; // @[FanNetwork.scala 1517:53]
  wire [31:0] w_vn_lvl_2_7 = my_adder_27_io_o_vn[63:32]; // @[FanNetwork.scala 1514:41]
  wire  _GEN_223 = w_vn_lvl_2_valid_7 | r_lvl_output_ff_valid_60; // @[FanNetwork.scala 755:40 757:35 760:35]
  wire  w_vn_lvl_3_valid_0 = my_adder_7_io_o_vn_valid[0]; // @[FanNetwork.scala 1147:53]
  wire [31:0] w_vn_lvl_3_0 = my_adder_7_io_o_vn[31:0]; // @[FanNetwork.scala 1144:40]
  wire  _GEN_225 = w_vn_lvl_3_valid_0 | r_lvl_output_ff_valid_71; // @[FanNetwork.scala 795:40 797:34 800:34]
  wire  w_vn_lvl_3_valid_1 = my_adder_7_io_o_vn_valid[1]; // @[FanNetwork.scala 1148:53]
  wire [31:0] w_vn_lvl_3_1 = my_adder_7_io_o_vn[63:32]; // @[FanNetwork.scala 1145:40]
  wire  _GEN_227 = w_vn_lvl_3_valid_1 | r_lvl_output_ff_valid_72; // @[FanNetwork.scala 803:40 805:34 808:34]
  wire  w_vn_lvl_3_valid_2 = my_adder_23_io_o_vn_valid[0]; // @[FanNetwork.scala 1442:53]
  wire [31:0] w_vn_lvl_3_2 = my_adder_23_io_o_vn[31:0]; // @[FanNetwork.scala 1439:41]
  wire  _GEN_229 = w_vn_lvl_3_valid_2 | r_lvl_output_ff_valid_87; // @[FanNetwork.scala 853:40 855:36 858:36]
  wire  w_vn_lvl_3_valid_3 = my_adder_23_io_o_vn_valid[1]; // @[FanNetwork.scala 1443:53]
  wire [31:0] w_vn_lvl_3_3 = my_adder_23_io_o_vn[63:32]; // @[FanNetwork.scala 1440:41]
  wire  _GEN_231 = w_vn_lvl_3_valid_3 | r_lvl_output_ff_valid_88; // @[FanNetwork.scala 861:41 863:36 866:36]
  wire  w_vn_lvl_4_valid_0 = my_adder_15_io_o_vn_valid[0]; // @[FanNetwork.scala 1293:53]
  wire [31:0] w_vn_lvl_4_0 = my_adder_15_io_o_vn[31:0]; // @[FanNetwork.scala 1290:41]
  wire  _GEN_233 = w_vn_lvl_4_valid_0 | r_lvl_output_ff_valid_111; // @[FanNetwork.scala 944:40 946:36 949:36]
  wire  w_vn_lvl_4_valid_1 = my_adder_15_io_o_vn_valid[1]; // @[FanNetwork.scala 1294:53]
  wire [31:0] w_vn_lvl_4_1 = my_adder_15_io_o_vn[63:32]; // @[FanNetwork.scala 1291:41]
  wire  _GEN_235 = w_vn_lvl_4_valid_1 | r_lvl_output_ff_valid_112; // @[FanNetwork.scala 952:40 954:36 957:36]
  wire [1:0] my_adder_7_io_i_sel_lo = {io_i_sel_bus_9,io_i_sel_bus_8}; // @[Cat.scala 33:92]
  wire [1:0] my_adder_7_io_i_sel_hi = {io_i_sel_bus_11,io_i_sel_bus_10}; // @[Cat.scala 33:92]
  wire [1:0] _my_adder_15_io_i_sel_T = {io_i_sel_bus_19,io_i_sel_bus_16}; // @[Cat.scala 33:92]
  wire [1:0] _my_adder_23_io_i_sel_T = {io_i_sel_bus_15,io_i_sel_bus_12}; // @[Cat.scala 33:92]
  wire [959:0] w_fan_lvl_0_0 = {{928'd0}, my_adder_0_io_o_adder};
  wire [959:0] w_fan_lvl_0_1 = {{928'd0}, my_adder_2_io_o_adder_0};
  wire [959:0] w_fan_lvl_0_2 = {{928'd0}, my_adder_2_io_o_adder_1};
  wire [959:0] w_fan_lvl_0_3 = {{928'd0}, my_adder_4_io_o_adder_0};
  wire [959:0] w_fan_lvl_0_4 = {{928'd0}, my_adder_4_io_o_adder_1};
  wire [959:0] w_fan_lvl_0_5 = {{928'd0}, my_adder_6_io_o_adder_0};
  wire [959:0] w_fan_lvl_0_6 = {{928'd0}, my_adder_6_io_o_adder_1};
  wire [959:0] w_fan_lvl_0_7 = {{928'd0}, my_adder_8_io_o_adder_0};
  wire [959:0] w_fan_lvl_0_8 = {{928'd0}, my_adder_8_io_o_adder_1};
  wire [959:0] w_fan_lvl_0_9 = {{928'd0}, my_adder_10_io_o_adder_0};
  wire [959:0] w_fan_lvl_0_10 = {{928'd0}, my_adder_10_io_o_adder_1};
  wire [959:0] w_fan_lvl_0_11 = {{928'd0}, my_adder_12_io_o_adder_0};
  wire [959:0] w_fan_lvl_0_12 = {{928'd0}, my_adder_12_io_o_adder_1};
  wire [959:0] w_fan_lvl_0_14 = {{928'd0}, my_adder_14_io_o_adder_1};
  wire [959:0] w_fan_lvl_0_15 = {{928'd0}, my_adder_16_io_o_adder_0};
  wire [959:0] w_fan_lvl_0_16 = {{928'd0}, my_adder_16_io_o_adder_1};
  wire [959:0] w_fan_lvl_0_18 = {{928'd0}, my_adder_18_io_o_adder_1};
  wire [959:0] w_fan_lvl_0_19 = {{928'd0}, my_adder_20_io_o_adder_0};
  wire [959:0] w_fan_lvl_0_20 = {{928'd0}, my_adder_20_io_o_adder_1};
  wire [959:0] w_fan_lvl_0_22 = {{928'd0}, my_adder_22_io_o_adder_1};
  wire [959:0] w_fan_lvl_0_23 = {{928'd0}, my_adder_24_io_o_adder_0};
  wire [959:0] w_fan_lvl_0_24 = {{928'd0}, my_adder_24_io_o_adder_1};
  wire [959:0] w_fan_lvl_0_26 = {{928'd0}, my_adder_26_io_o_adder_1};
  wire [959:0] w_fan_lvl_0_27 = {{928'd0}, my_adder_28_io_o_adder_0};
  wire [959:0] w_fan_lvl_0_28 = {{928'd0}, my_adder_28_io_o_adder_1};
  wire [479:0] w_fan_lvl_1_0 = {{448'd0}, my_adder_1_io_o_adder};
  wire [479:0] w_fan_lvl_1_1 = {{448'd0}, my_adder_5_io_o_adder_0};
  wire [479:0] w_fan_lvl_1_2 = {{448'd0}, my_adder_5_io_o_adder_1};
  wire [479:0] w_fan_lvl_1_3 = {{448'd0}, my_adder_9_io_o_adder_0};
  wire [479:0] w_fan_lvl_1_4 = {{448'd0}, my_adder_9_io_o_adder_1};
  wire [479:0] w_fan_lvl_1_5 = {{448'd0}, my_adder_13_io_o_adder_0};
  wire [479:0] w_fan_lvl_1_6 = {{448'd0}, my_adder_13_io_o_adder_1};
  wire [479:0] w_fan_lvl_1_7 = {{448'd0}, my_adder_17_io_o_adder_0};
  wire [479:0] w_fan_lvl_1_8 = {{448'd0}, my_adder_17_io_o_adder_1};
  wire [479:0] w_fan_lvl_1_9 = {{448'd0}, my_adder_21_io_o_adder_0};
  wire [479:0] w_fan_lvl_1_10 = {{448'd0}, my_adder_21_io_o_adder_1};
  wire [479:0] w_fan_lvl_1_11 = {{448'd0}, my_adder_25_io_o_adder_0};
  wire [479:0] w_fan_lvl_1_12 = {{448'd0}, my_adder_25_io_o_adder_1};
  wire [479:0] w_fan_lvl_1_13 = {{448'd0}, my_adder_29_io_o_adder};
  wire [191:0] w_fan_lvl_2_0 = {{160'd0}, my_adder_3_io_o_adder};
  wire [191:0] w_fan_lvl_2_1 = {{160'd0}, my_adder_11_io_o_adder_0};
  wire [191:0] w_fan_lvl_2_2 = {{160'd0}, my_adder_11_io_o_adder_1};
  wire [191:0] w_fan_lvl_2_3 = {{160'd0}, my_adder_19_io_o_adder_0};
  wire [191:0] w_fan_lvl_2_4 = {{160'd0}, my_adder_19_io_o_adder_1};
  wire [191:0] w_fan_lvl_2_5 = {{160'd0}, my_adder_27_io_o_adder};
  wire [31:0] w_fan_lvl_4_0 = my_adder_15_io_o_adder;
  wire [479:0] _WIRE_9_1 = {{448'd0}, r_fan_ff_lvl_0_to_2_1}; // @[FanNetwork.scala 1067:{42,42}]
  wire [479:0] _WIRE_9_2 = {{448'd0}, r_fan_ff_lvl_0_to_2_0}; // @[FanNetwork.scala 1067:{42,42}]
  wire [191:0] _WIRE_13_1 = {{160'd0}, r_fan_ff_lvl_1_to_3_1}; // @[FanNetwork.scala 1138:{40,40}]
  wire [191:0] _WIRE_13_2 = {{160'd0}, r_fan_ff_lvl_0_to_3_1}; // @[FanNetwork.scala 1138:{40,40}]
  wire [191:0] _WIRE_13_3 = {{160'd0}, r_fan_ff_lvl_0_to_3_0}; // @[FanNetwork.scala 1138:{40,40}]
  wire [191:0] _WIRE_13_4 = {{160'd0}, r_fan_ff_lvl_1_to_3_0}; // @[FanNetwork.scala 1138:{40,40}]
  wire [479:0] _WIRE_17_1 = {{448'd0}, r_fan_ff_lvl_0_to_2_5}; // @[FanNetwork.scala 1208:{41,41}]
  wire [479:0] _WIRE_17_2 = {{448'd0}, r_fan_ff_lvl_0_to_2_4}; // @[FanNetwork.scala 1208:{41,41}]
  wire [479:0] _WIRE_25_1 = {{448'd0}, r_fan_ff_lvl_0_to_2_9}; // @[FanNetwork.scala 1357:{42,42}]
  wire [479:0] _WIRE_25_2 = {{448'd0}, r_fan_ff_lvl_0_to_2_8}; // @[FanNetwork.scala 1357:{42,42}]
  wire [191:0] _WIRE_29_1 = {{160'd0}, r_fan_ff_lvl_1_to_3_5}; // @[FanNetwork.scala 1434:{41,41}]
  wire [191:0] _WIRE_29_2 = {{160'd0}, r_fan_ff_lvl_0_to_3_5}; // @[FanNetwork.scala 1434:{41,41}]
  wire [191:0] _WIRE_29_3 = {{160'd0}, r_fan_ff_lvl_0_to_3_4}; // @[FanNetwork.scala 1434:{41,41}]
  wire [191:0] _WIRE_29_4 = {{160'd0}, r_fan_ff_lvl_1_to_3_4}; // @[FanNetwork.scala 1434:{41,41}]
  wire [479:0] _WIRE_33_1 = {{448'd0}, r_fan_ff_lvl_0_to_2_13}; // @[FanNetwork.scala 1508:{41,41}]
  wire [479:0] _WIRE_33_2 = {{448'd0}, r_fan_ff_lvl_0_to_2_12}; // @[FanNetwork.scala 1508:{41,41}]
  wire [959:0] _GEN_239 = reset ? 960'h0 : w_fan_lvl_0_2; // @[FanNetwork.scala 34:{38,38} 73:25]
  wire [959:0] _GEN_240 = reset ? 960'h0 : w_fan_lvl_0_3; // @[FanNetwork.scala 34:{38,38} 73:25]
  wire [959:0] _GEN_241 = reset ? 960'h0 : w_fan_lvl_0_6; // @[FanNetwork.scala 34:{38,38} 73:25]
  wire [959:0] _GEN_242 = reset ? 960'h0 : w_fan_lvl_0_7; // @[FanNetwork.scala 34:{38,38} 73:25]
  wire [959:0] _GEN_243 = reset ? 960'h0 : w_fan_lvl_0_10; // @[FanNetwork.scala 34:{38,38} 73:25]
  wire [959:0] _GEN_244 = reset ? 960'h0 : w_fan_lvl_0_11; // @[FanNetwork.scala 34:{38,38} 73:25]
  wire [959:0] _GEN_245 = reset ? 960'h0 : w_fan_lvl_0_14; // @[FanNetwork.scala 34:{38,38} 73:25]
  wire [959:0] _GEN_246 = reset ? 960'h0 : w_fan_lvl_0_15; // @[FanNetwork.scala 34:{38,38} 73:25]
  wire [959:0] _GEN_247 = reset ? 960'h0 : w_fan_lvl_0_18; // @[FanNetwork.scala 34:{38,38} 73:25]
  wire [959:0] _GEN_248 = reset ? 960'h0 : w_fan_lvl_0_19; // @[FanNetwork.scala 34:{38,38} 73:25]
  wire [959:0] _GEN_249 = reset ? 960'h0 : w_fan_lvl_0_22; // @[FanNetwork.scala 34:{38,38} 73:25]
  wire [959:0] _GEN_250 = reset ? 960'h0 : w_fan_lvl_0_23; // @[FanNetwork.scala 34:{38,38} 73:25]
  wire [959:0] _GEN_251 = reset ? 960'h0 : w_fan_lvl_0_26; // @[FanNetwork.scala 34:{38,38} 73:25]
  wire [959:0] _GEN_252 = reset ? 960'h0 : w_fan_lvl_0_27; // @[FanNetwork.scala 34:{38,38} 73:25]
  wire [479:0] _GEN_253 = reset ? 480'h0 : w_fan_lvl_1_2; // @[FanNetwork.scala 36:{38,38} 77:25]
  wire [479:0] _GEN_254 = reset ? 480'h0 : w_fan_lvl_1_3; // @[FanNetwork.scala 36:{38,38} 77:25]
  wire [479:0] _GEN_255 = reset ? 480'h0 : w_fan_lvl_1_6; // @[FanNetwork.scala 36:{38,38} 77:25]
  wire [479:0] _GEN_256 = reset ? 480'h0 : w_fan_lvl_1_7; // @[FanNetwork.scala 36:{38,38} 77:25]
  wire [479:0] _GEN_257 = reset ? 480'h0 : w_fan_lvl_1_10; // @[FanNetwork.scala 36:{38,38} 77:25]
  wire [479:0] _GEN_258 = reset ? 480'h0 : w_fan_lvl_1_11; // @[FanNetwork.scala 36:{38,38} 77:25]
  wire [191:0] _GEN_259 = reset ? 192'h0 : w_fan_lvl_2_2; // @[FanNetwork.scala 37:{38,38} 78:25]
  wire [191:0] _GEN_260 = reset ? 192'h0 : w_fan_lvl_2_3; // @[FanNetwork.scala 37:{38,38} 78:25]
  EdgeAdderSwitch my_adder_0 ( // @[FanNetwork.scala 1018:28]
    .clock(my_adder_0_clock),
    .reset(my_adder_0_reset),
    .io_i_valid(my_adder_0_io_i_valid),
    .io_i_data_bus_0(my_adder_0_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_0_io_i_data_bus_1),
    .io_i_add_en(my_adder_0_io_i_add_en),
    .io_i_cmd(my_adder_0_io_i_cmd),
    .io_o_vn(my_adder_0_io_o_vn),
    .io_o_vn_valid(my_adder_0_io_o_vn_valid),
    .io_o_adder(my_adder_0_io_o_adder)
  );
  EdgeAdderSwitch my_adder_1 ( // @[FanNetwork.scala 1031:28]
    .clock(my_adder_1_clock),
    .reset(my_adder_1_reset),
    .io_i_valid(my_adder_1_io_i_valid),
    .io_i_data_bus_0(my_adder_1_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_1_io_i_data_bus_1),
    .io_i_add_en(my_adder_1_io_i_add_en),
    .io_i_cmd(my_adder_1_io_i_cmd),
    .io_o_vn(my_adder_1_io_o_vn),
    .io_o_vn_valid(my_adder_1_io_o_vn_valid),
    .io_o_adder(my_adder_1_io_o_adder)
  );
  AdderSwitch my_adder_2 ( // @[FanNetwork.scala 1045:28]
    .clock(my_adder_2_clock),
    .reset(my_adder_2_reset),
    .io_i_valid(my_adder_2_io_i_valid),
    .io_i_data_bus_0(my_adder_2_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_2_io_i_data_bus_1),
    .io_i_add_en(my_adder_2_io_i_add_en),
    .io_i_cmd(my_adder_2_io_i_cmd),
    .io_o_vn_valid(my_adder_2_io_o_vn_valid),
    .io_o_vn(my_adder_2_io_o_vn),
    .io_o_adder_0(my_adder_2_io_o_adder_0),
    .io_o_adder_1(my_adder_2_io_o_adder_1)
  );
  EdgeAdderSwitch_2 my_adder_3 ( // @[FanNetwork.scala 1064:28]
    .clock(my_adder_3_clock),
    .reset(my_adder_3_reset),
    .io_i_valid(my_adder_3_io_i_valid),
    .io_i_data_bus_0(my_adder_3_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_3_io_i_data_bus_1),
    .io_i_data_bus_2(my_adder_3_io_i_data_bus_2),
    .io_i_data_bus_3(my_adder_3_io_i_data_bus_3),
    .io_i_add_en(my_adder_3_io_i_add_en),
    .io_i_cmd(my_adder_3_io_i_cmd),
    .io_i_sel(my_adder_3_io_i_sel),
    .io_o_vn(my_adder_3_io_o_vn),
    .io_o_vn_valid(my_adder_3_io_o_vn_valid),
    .io_o_adder(my_adder_3_io_o_adder)
  );
  AdderSwitch my_adder_4 ( // @[FanNetwork.scala 1081:28]
    .clock(my_adder_4_clock),
    .reset(my_adder_4_reset),
    .io_i_valid(my_adder_4_io_i_valid),
    .io_i_data_bus_0(my_adder_4_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_4_io_i_data_bus_1),
    .io_i_add_en(my_adder_4_io_i_add_en),
    .io_i_cmd(my_adder_4_io_i_cmd),
    .io_o_vn_valid(my_adder_4_io_o_vn_valid),
    .io_o_vn(my_adder_4_io_o_vn),
    .io_o_adder_0(my_adder_4_io_o_adder_0),
    .io_o_adder_1(my_adder_4_io_o_adder_1)
  );
  AdderSwitch my_adder_5 ( // @[FanNetwork.scala 1099:28]
    .clock(my_adder_5_clock),
    .reset(my_adder_5_reset),
    .io_i_valid(my_adder_5_io_i_valid),
    .io_i_data_bus_0(my_adder_5_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_5_io_i_data_bus_1),
    .io_i_add_en(my_adder_5_io_i_add_en),
    .io_i_cmd(my_adder_5_io_i_cmd),
    .io_o_vn_valid(my_adder_5_io_o_vn_valid),
    .io_o_vn(my_adder_5_io_o_vn),
    .io_o_adder_0(my_adder_5_io_o_adder_0),
    .io_o_adder_1(my_adder_5_io_o_adder_1)
  );
  AdderSwitch my_adder_6 ( // @[FanNetwork.scala 1116:28]
    .clock(my_adder_6_clock),
    .reset(my_adder_6_reset),
    .io_i_valid(my_adder_6_io_i_valid),
    .io_i_data_bus_0(my_adder_6_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_6_io_i_data_bus_1),
    .io_i_add_en(my_adder_6_io_i_add_en),
    .io_i_cmd(my_adder_6_io_i_cmd),
    .io_o_vn_valid(my_adder_6_io_o_vn_valid),
    .io_o_vn(my_adder_6_io_o_vn),
    .io_o_adder_0(my_adder_6_io_o_adder_0),
    .io_o_adder_1(my_adder_6_io_o_adder_1)
  );
  EdgeAdderSwitch_3 my_adder_7 ( // @[FanNetwork.scala 1133:28]
    .clock(my_adder_7_clock),
    .reset(my_adder_7_reset),
    .io_i_valid(my_adder_7_io_i_valid),
    .io_i_data_bus_0(my_adder_7_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_7_io_i_data_bus_1),
    .io_i_data_bus_2(my_adder_7_io_i_data_bus_2),
    .io_i_data_bus_3(my_adder_7_io_i_data_bus_3),
    .io_i_data_bus_4(my_adder_7_io_i_data_bus_4),
    .io_i_data_bus_5(my_adder_7_io_i_data_bus_5),
    .io_i_add_en(my_adder_7_io_i_add_en),
    .io_i_cmd(my_adder_7_io_i_cmd),
    .io_i_sel(my_adder_7_io_i_sel),
    .io_o_vn(my_adder_7_io_o_vn),
    .io_o_vn_valid(my_adder_7_io_o_vn_valid),
    .io_o_adder(my_adder_7_io_o_adder)
  );
  AdderSwitch my_adder_8 ( // @[FanNetwork.scala 1152:28]
    .clock(my_adder_8_clock),
    .reset(my_adder_8_reset),
    .io_i_valid(my_adder_8_io_i_valid),
    .io_i_data_bus_0(my_adder_8_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_8_io_i_data_bus_1),
    .io_i_add_en(my_adder_8_io_i_add_en),
    .io_i_cmd(my_adder_8_io_i_cmd),
    .io_o_vn_valid(my_adder_8_io_o_vn_valid),
    .io_o_vn(my_adder_8_io_o_vn),
    .io_o_adder_0(my_adder_8_io_o_adder_0),
    .io_o_adder_1(my_adder_8_io_o_adder_1)
  );
  AdderSwitch my_adder_9 ( // @[FanNetwork.scala 1169:28]
    .clock(my_adder_9_clock),
    .reset(my_adder_9_reset),
    .io_i_valid(my_adder_9_io_i_valid),
    .io_i_data_bus_0(my_adder_9_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_9_io_i_data_bus_1),
    .io_i_add_en(my_adder_9_io_i_add_en),
    .io_i_cmd(my_adder_9_io_i_cmd),
    .io_o_vn_valid(my_adder_9_io_o_vn_valid),
    .io_o_vn(my_adder_9_io_o_vn),
    .io_o_adder_0(my_adder_9_io_o_adder_0),
    .io_o_adder_1(my_adder_9_io_o_adder_1)
  );
  AdderSwitch my_adder_10 ( // @[FanNetwork.scala 1186:29]
    .clock(my_adder_10_clock),
    .reset(my_adder_10_reset),
    .io_i_valid(my_adder_10_io_i_valid),
    .io_i_data_bus_0(my_adder_10_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_10_io_i_data_bus_1),
    .io_i_add_en(my_adder_10_io_i_add_en),
    .io_i_cmd(my_adder_10_io_i_cmd),
    .io_o_vn_valid(my_adder_10_io_o_vn_valid),
    .io_o_vn(my_adder_10_io_o_vn),
    .io_o_adder_0(my_adder_10_io_o_adder_0),
    .io_o_adder_1(my_adder_10_io_o_adder_1)
  );
  AdderSwitch_7 my_adder_11 ( // @[FanNetwork.scala 1204:29]
    .clock(my_adder_11_clock),
    .reset(my_adder_11_reset),
    .io_i_valid(my_adder_11_io_i_valid),
    .io_i_data_bus_0(my_adder_11_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_11_io_i_data_bus_1),
    .io_i_data_bus_2(my_adder_11_io_i_data_bus_2),
    .io_i_data_bus_3(my_adder_11_io_i_data_bus_3),
    .io_i_add_en(my_adder_11_io_i_add_en),
    .io_i_cmd(my_adder_11_io_i_cmd),
    .io_i_sel(my_adder_11_io_i_sel),
    .io_o_vn_valid(my_adder_11_io_o_vn_valid),
    .io_o_vn(my_adder_11_io_o_vn),
    .io_o_adder_0(my_adder_11_io_o_adder_0),
    .io_o_adder_1(my_adder_11_io_o_adder_1)
  );
  AdderSwitch my_adder_12 ( // @[FanNetwork.scala 1225:29]
    .clock(my_adder_12_clock),
    .reset(my_adder_12_reset),
    .io_i_valid(my_adder_12_io_i_valid),
    .io_i_data_bus_0(my_adder_12_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_12_io_i_data_bus_1),
    .io_i_add_en(my_adder_12_io_i_add_en),
    .io_i_cmd(my_adder_12_io_i_cmd),
    .io_o_vn_valid(my_adder_12_io_o_vn_valid),
    .io_o_vn(my_adder_12_io_o_vn),
    .io_o_adder_0(my_adder_12_io_o_adder_0),
    .io_o_adder_1(my_adder_12_io_o_adder_1)
  );
  AdderSwitch my_adder_13 ( // @[FanNetwork.scala 1243:29]
    .clock(my_adder_13_clock),
    .reset(my_adder_13_reset),
    .io_i_valid(my_adder_13_io_i_valid),
    .io_i_data_bus_0(my_adder_13_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_13_io_i_data_bus_1),
    .io_i_add_en(my_adder_13_io_i_add_en),
    .io_i_cmd(my_adder_13_io_i_cmd),
    .io_o_vn_valid(my_adder_13_io_o_vn_valid),
    .io_o_vn(my_adder_13_io_o_vn),
    .io_o_adder_0(my_adder_13_io_o_adder_0),
    .io_o_adder_1(my_adder_13_io_o_adder_1)
  );
  AdderSwitch my_adder_14 ( // @[FanNetwork.scala 1261:29]
    .clock(my_adder_14_clock),
    .reset(my_adder_14_reset),
    .io_i_valid(my_adder_14_io_i_valid),
    .io_i_data_bus_0(my_adder_14_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_14_io_i_data_bus_1),
    .io_i_add_en(my_adder_14_io_i_add_en),
    .io_i_cmd(my_adder_14_io_i_cmd),
    .io_o_vn_valid(my_adder_14_io_o_vn_valid),
    .io_o_vn(my_adder_14_io_o_vn),
    .io_o_adder_0(my_adder_14_io_o_adder_0),
    .io_o_adder_1(my_adder_14_io_o_adder_1)
  );
  EdgeAdderSwitch_4 my_adder_15 ( // @[FanNetwork.scala 1279:29]
    .clock(my_adder_15_clock),
    .reset(my_adder_15_reset),
    .io_i_valid(my_adder_15_io_i_valid),
    .io_i_data_bus_0(my_adder_15_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_15_io_i_data_bus_1),
    .io_i_data_bus_2(my_adder_15_io_i_data_bus_2),
    .io_i_data_bus_3(my_adder_15_io_i_data_bus_3),
    .io_i_data_bus_4(my_adder_15_io_i_data_bus_4),
    .io_i_data_bus_5(my_adder_15_io_i_data_bus_5),
    .io_i_data_bus_6(my_adder_15_io_i_data_bus_6),
    .io_i_data_bus_7(my_adder_15_io_i_data_bus_7),
    .io_i_add_en(my_adder_15_io_i_add_en),
    .io_i_cmd(my_adder_15_io_i_cmd),
    .io_i_sel(my_adder_15_io_i_sel),
    .io_o_vn(my_adder_15_io_o_vn),
    .io_o_vn_valid(my_adder_15_io_o_vn_valid),
    .io_o_adder(my_adder_15_io_o_adder)
  );
  AdderSwitch my_adder_16 ( // @[FanNetwork.scala 1299:29]
    .clock(my_adder_16_clock),
    .reset(my_adder_16_reset),
    .io_i_valid(my_adder_16_io_i_valid),
    .io_i_data_bus_0(my_adder_16_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_16_io_i_data_bus_1),
    .io_i_add_en(my_adder_16_io_i_add_en),
    .io_i_cmd(my_adder_16_io_i_cmd),
    .io_o_vn_valid(my_adder_16_io_o_vn_valid),
    .io_o_vn(my_adder_16_io_o_vn),
    .io_o_adder_0(my_adder_16_io_o_adder_0),
    .io_o_adder_1(my_adder_16_io_o_adder_1)
  );
  AdderSwitch my_adder_17 ( // @[FanNetwork.scala 1317:29]
    .clock(my_adder_17_clock),
    .reset(my_adder_17_reset),
    .io_i_valid(my_adder_17_io_i_valid),
    .io_i_data_bus_0(my_adder_17_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_17_io_i_data_bus_1),
    .io_i_add_en(my_adder_17_io_i_add_en),
    .io_i_cmd(my_adder_17_io_i_cmd),
    .io_o_vn_valid(my_adder_17_io_o_vn_valid),
    .io_o_vn(my_adder_17_io_o_vn),
    .io_o_adder_0(my_adder_17_io_o_adder_0),
    .io_o_adder_1(my_adder_17_io_o_adder_1)
  );
  AdderSwitch my_adder_18 ( // @[FanNetwork.scala 1335:29]
    .clock(my_adder_18_clock),
    .reset(my_adder_18_reset),
    .io_i_valid(my_adder_18_io_i_valid),
    .io_i_data_bus_0(my_adder_18_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_18_io_i_data_bus_1),
    .io_i_add_en(my_adder_18_io_i_add_en),
    .io_i_cmd(my_adder_18_io_i_cmd),
    .io_o_vn_valid(my_adder_18_io_o_vn_valid),
    .io_o_vn(my_adder_18_io_o_vn),
    .io_o_adder_0(my_adder_18_io_o_adder_0),
    .io_o_adder_1(my_adder_18_io_o_adder_1)
  );
  AdderSwitch_7 my_adder_19 ( // @[FanNetwork.scala 1353:29]
    .clock(my_adder_19_clock),
    .reset(my_adder_19_reset),
    .io_i_valid(my_adder_19_io_i_valid),
    .io_i_data_bus_0(my_adder_19_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_19_io_i_data_bus_1),
    .io_i_data_bus_2(my_adder_19_io_i_data_bus_2),
    .io_i_data_bus_3(my_adder_19_io_i_data_bus_3),
    .io_i_add_en(my_adder_19_io_i_add_en),
    .io_i_cmd(my_adder_19_io_i_cmd),
    .io_i_sel(my_adder_19_io_i_sel),
    .io_o_vn_valid(my_adder_19_io_o_vn_valid),
    .io_o_vn(my_adder_19_io_o_vn),
    .io_o_adder_0(my_adder_19_io_o_adder_0),
    .io_o_adder_1(my_adder_19_io_o_adder_1)
  );
  AdderSwitch my_adder_20 ( // @[FanNetwork.scala 1373:29]
    .clock(my_adder_20_clock),
    .reset(my_adder_20_reset),
    .io_i_valid(my_adder_20_io_i_valid),
    .io_i_data_bus_0(my_adder_20_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_20_io_i_data_bus_1),
    .io_i_add_en(my_adder_20_io_i_add_en),
    .io_i_cmd(my_adder_20_io_i_cmd),
    .io_o_vn_valid(my_adder_20_io_o_vn_valid),
    .io_o_vn(my_adder_20_io_o_vn),
    .io_o_adder_0(my_adder_20_io_o_adder_0),
    .io_o_adder_1(my_adder_20_io_o_adder_1)
  );
  AdderSwitch my_adder_21 ( // @[FanNetwork.scala 1393:29]
    .clock(my_adder_21_clock),
    .reset(my_adder_21_reset),
    .io_i_valid(my_adder_21_io_i_valid),
    .io_i_data_bus_0(my_adder_21_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_21_io_i_data_bus_1),
    .io_i_add_en(my_adder_21_io_i_add_en),
    .io_i_cmd(my_adder_21_io_i_cmd),
    .io_o_vn_valid(my_adder_21_io_o_vn_valid),
    .io_o_vn(my_adder_21_io_o_vn),
    .io_o_adder_0(my_adder_21_io_o_adder_0),
    .io_o_adder_1(my_adder_21_io_o_adder_1)
  );
  AdderSwitch my_adder_22 ( // @[FanNetwork.scala 1412:29]
    .clock(my_adder_22_clock),
    .reset(my_adder_22_reset),
    .io_i_valid(my_adder_22_io_i_valid),
    .io_i_data_bus_0(my_adder_22_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_22_io_i_data_bus_1),
    .io_i_add_en(my_adder_22_io_i_add_en),
    .io_i_cmd(my_adder_22_io_i_cmd),
    .io_o_vn_valid(my_adder_22_io_o_vn_valid),
    .io_o_vn(my_adder_22_io_o_vn),
    .io_o_adder_0(my_adder_22_io_o_adder_0),
    .io_o_adder_1(my_adder_22_io_o_adder_1)
  );
  EdgeAdderSwitch_3 my_adder_23 ( // @[FanNetwork.scala 1430:29]
    .clock(my_adder_23_clock),
    .reset(my_adder_23_reset),
    .io_i_valid(my_adder_23_io_i_valid),
    .io_i_data_bus_0(my_adder_23_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_23_io_i_data_bus_1),
    .io_i_data_bus_2(my_adder_23_io_i_data_bus_2),
    .io_i_data_bus_3(my_adder_23_io_i_data_bus_3),
    .io_i_data_bus_4(my_adder_23_io_i_data_bus_4),
    .io_i_data_bus_5(my_adder_23_io_i_data_bus_5),
    .io_i_add_en(my_adder_23_io_i_add_en),
    .io_i_cmd(my_adder_23_io_i_cmd),
    .io_i_sel(my_adder_23_io_i_sel),
    .io_o_vn(my_adder_23_io_o_vn),
    .io_o_vn_valid(my_adder_23_io_o_vn_valid),
    .io_o_adder(my_adder_23_io_o_adder)
  );
  AdderSwitch my_adder_24 ( // @[FanNetwork.scala 1447:29]
    .clock(my_adder_24_clock),
    .reset(my_adder_24_reset),
    .io_i_valid(my_adder_24_io_i_valid),
    .io_i_data_bus_0(my_adder_24_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_24_io_i_data_bus_1),
    .io_i_add_en(my_adder_24_io_i_add_en),
    .io_i_cmd(my_adder_24_io_i_cmd),
    .io_o_vn_valid(my_adder_24_io_o_vn_valid),
    .io_o_vn(my_adder_24_io_o_vn),
    .io_o_adder_0(my_adder_24_io_o_adder_0),
    .io_o_adder_1(my_adder_24_io_o_adder_1)
  );
  AdderSwitch my_adder_25 ( // @[FanNetwork.scala 1466:29]
    .clock(my_adder_25_clock),
    .reset(my_adder_25_reset),
    .io_i_valid(my_adder_25_io_i_valid),
    .io_i_data_bus_0(my_adder_25_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_25_io_i_data_bus_1),
    .io_i_add_en(my_adder_25_io_i_add_en),
    .io_i_cmd(my_adder_25_io_i_cmd),
    .io_o_vn_valid(my_adder_25_io_o_vn_valid),
    .io_o_vn(my_adder_25_io_o_vn),
    .io_o_adder_0(my_adder_25_io_o_adder_0),
    .io_o_adder_1(my_adder_25_io_o_adder_1)
  );
  AdderSwitch my_adder_26 ( // @[FanNetwork.scala 1486:29]
    .clock(my_adder_26_clock),
    .reset(my_adder_26_reset),
    .io_i_valid(my_adder_26_io_i_valid),
    .io_i_data_bus_0(my_adder_26_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_26_io_i_data_bus_1),
    .io_i_add_en(my_adder_26_io_i_add_en),
    .io_i_cmd(my_adder_26_io_i_cmd),
    .io_o_vn_valid(my_adder_26_io_o_vn_valid),
    .io_o_vn(my_adder_26_io_o_vn),
    .io_o_adder_0(my_adder_26_io_o_adder_0),
    .io_o_adder_1(my_adder_26_io_o_adder_1)
  );
  EdgeAdderSwitch_2 my_adder_27 ( // @[FanNetwork.scala 1504:29]
    .clock(my_adder_27_clock),
    .reset(my_adder_27_reset),
    .io_i_valid(my_adder_27_io_i_valid),
    .io_i_data_bus_0(my_adder_27_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_27_io_i_data_bus_1),
    .io_i_data_bus_2(my_adder_27_io_i_data_bus_2),
    .io_i_data_bus_3(my_adder_27_io_i_data_bus_3),
    .io_i_add_en(my_adder_27_io_i_add_en),
    .io_i_cmd(my_adder_27_io_i_cmd),
    .io_i_sel(my_adder_27_io_i_sel),
    .io_o_vn(my_adder_27_io_o_vn),
    .io_o_vn_valid(my_adder_27_io_o_vn_valid),
    .io_o_adder(my_adder_27_io_o_adder)
  );
  AdderSwitch my_adder_28 ( // @[FanNetwork.scala 1525:29]
    .clock(my_adder_28_clock),
    .reset(my_adder_28_reset),
    .io_i_valid(my_adder_28_io_i_valid),
    .io_i_data_bus_0(my_adder_28_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_28_io_i_data_bus_1),
    .io_i_add_en(my_adder_28_io_i_add_en),
    .io_i_cmd(my_adder_28_io_i_cmd),
    .io_o_vn_valid(my_adder_28_io_o_vn_valid),
    .io_o_vn(my_adder_28_io_o_vn),
    .io_o_adder_0(my_adder_28_io_o_adder_0),
    .io_o_adder_1(my_adder_28_io_o_adder_1)
  );
  EdgeAdderSwitch my_adder_29 ( // @[FanNetwork.scala 1544:29]
    .clock(my_adder_29_clock),
    .reset(my_adder_29_reset),
    .io_i_valid(my_adder_29_io_i_valid),
    .io_i_data_bus_0(my_adder_29_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_29_io_i_data_bus_1),
    .io_i_add_en(my_adder_29_io_i_add_en),
    .io_i_cmd(my_adder_29_io_i_cmd),
    .io_o_vn(my_adder_29_io_o_vn),
    .io_o_vn_valid(my_adder_29_io_o_vn_valid),
    .io_o_adder(my_adder_29_io_o_adder)
  );
  EdgeAdderSwitch my_adder_30 ( // @[FanNetwork.scala 1562:29]
    .clock(my_adder_30_clock),
    .reset(my_adder_30_reset),
    .io_i_valid(my_adder_30_io_i_valid),
    .io_i_data_bus_0(my_adder_30_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_30_io_i_data_bus_1),
    .io_i_add_en(my_adder_30_io_i_add_en),
    .io_i_cmd(my_adder_30_io_i_cmd),
    .io_o_vn(my_adder_30_io_o_vn),
    .io_o_vn_valid(my_adder_30_io_o_vn_valid),
    .io_o_adder(my_adder_30_io_o_adder)
  );
  assign io_o_valid_0 = r_lvl_output_ff_valid_128; // @[FanNetwork.scala 1710:19]
  assign io_o_valid_1 = r_lvl_output_ff_valid_129; // @[FanNetwork.scala 1711:19]
  assign io_o_valid_2 = r_lvl_output_ff_valid_130; // @[FanNetwork.scala 1712:19]
  assign io_o_valid_3 = r_lvl_output_ff_valid_131; // @[FanNetwork.scala 1713:19]
  assign io_o_valid_4 = r_lvl_output_ff_valid_132; // @[FanNetwork.scala 1714:19]
  assign io_o_valid_5 = r_lvl_output_ff_valid_133; // @[FanNetwork.scala 1715:19]
  assign io_o_valid_6 = r_lvl_output_ff_valid_134; // @[FanNetwork.scala 1716:19]
  assign io_o_valid_7 = r_lvl_output_ff_valid_135; // @[FanNetwork.scala 1717:19]
  assign io_o_valid_8 = r_lvl_output_ff_valid_136; // @[FanNetwork.scala 1718:19]
  assign io_o_valid_9 = r_lvl_output_ff_valid_137; // @[FanNetwork.scala 1719:19]
  assign io_o_valid_10 = r_lvl_output_ff_valid_138; // @[FanNetwork.scala 1720:20]
  assign io_o_valid_11 = r_lvl_output_ff_valid_139; // @[FanNetwork.scala 1721:20]
  assign io_o_valid_12 = r_lvl_output_ff_valid_140; // @[FanNetwork.scala 1722:20]
  assign io_o_valid_13 = r_lvl_output_ff_valid_141; // @[FanNetwork.scala 1723:20]
  assign io_o_valid_14 = r_lvl_output_ff_valid_142; // @[FanNetwork.scala 1724:20]
  assign io_o_valid_15 = r_final_add2 | r_lvl_output_ff_valid_143; // @[FanNetwork.scala 1725:33 1726:24 1728:25]
  assign io_o_valid_16 = r_lvl_output_ff_valid_144; // @[FanNetwork.scala 1730:20]
  assign io_o_valid_17 = r_lvl_output_ff_valid_145; // @[FanNetwork.scala 1731:20]
  assign io_o_valid_18 = r_lvl_output_ff_valid_146; // @[FanNetwork.scala 1732:20]
  assign io_o_valid_19 = r_lvl_output_ff_valid_147; // @[FanNetwork.scala 1733:20]
  assign io_o_valid_20 = r_lvl_output_ff_valid_148; // @[FanNetwork.scala 1734:20]
  assign io_o_valid_21 = r_lvl_output_ff_valid_149; // @[FanNetwork.scala 1735:20]
  assign io_o_valid_22 = r_lvl_output_ff_valid_150; // @[FanNetwork.scala 1736:20]
  assign io_o_valid_23 = r_lvl_output_ff_valid_151; // @[FanNetwork.scala 1737:20]
  assign io_o_valid_24 = r_lvl_output_ff_valid_152; // @[FanNetwork.scala 1738:20]
  assign io_o_valid_25 = r_lvl_output_ff_valid_153; // @[FanNetwork.scala 1739:20]
  assign io_o_valid_26 = r_lvl_output_ff_valid_154; // @[FanNetwork.scala 1740:20]
  assign io_o_valid_27 = r_lvl_output_ff_valid_155; // @[FanNetwork.scala 1741:20]
  assign io_o_valid_28 = r_lvl_output_ff_valid_156; // @[FanNetwork.scala 1742:20]
  assign io_o_valid_29 = r_lvl_output_ff_valid_157; // @[FanNetwork.scala 1743:20]
  assign io_o_valid_30 = r_lvl_output_ff_valid_158; // @[FanNetwork.scala 1744:20]
  assign io_o_valid_31 = r_lvl_output_ff_valid_159; // @[FanNetwork.scala 1745:20]
  assign io_o_data_bus_0 = r_lvl_output_ff_128; // @[FanNetwork.scala 1629:22]
  assign io_o_data_bus_1 = r_lvl_output_ff_129; // @[FanNetwork.scala 1630:22]
  assign io_o_data_bus_2 = r_lvl_output_ff_130; // @[FanNetwork.scala 1631:22]
  assign io_o_data_bus_3 = r_lvl_output_ff_131; // @[FanNetwork.scala 1632:22]
  assign io_o_data_bus_4 = r_lvl_output_ff_132; // @[FanNetwork.scala 1633:22]
  assign io_o_data_bus_5 = r_lvl_output_ff_133; // @[FanNetwork.scala 1634:22]
  assign io_o_data_bus_6 = r_lvl_output_ff_134; // @[FanNetwork.scala 1635:22]
  assign io_o_data_bus_7 = r_lvl_output_ff_135; // @[FanNetwork.scala 1636:22]
  assign io_o_data_bus_8 = r_lvl_output_ff_136; // @[FanNetwork.scala 1637:22]
  assign io_o_data_bus_9 = r_lvl_output_ff_137; // @[FanNetwork.scala 1638:22]
  assign io_o_data_bus_10 = r_lvl_output_ff_138; // @[FanNetwork.scala 1639:23]
  assign io_o_data_bus_11 = r_lvl_output_ff_139; // @[FanNetwork.scala 1640:23]
  assign io_o_data_bus_12 = r_lvl_output_ff_140; // @[FanNetwork.scala 1641:23]
  assign io_o_data_bus_13 = r_lvl_output_ff_141; // @[FanNetwork.scala 1642:23]
  assign io_o_data_bus_14 = r_lvl_output_ff_142; // @[FanNetwork.scala 1643:23]
  assign io_o_data_bus_15 = r_final_add2 ? r_final_sum : r_lvl_output_ff_143; // @[FanNetwork.scala 1645:33 1646:27 1648:27]
  assign io_o_data_bus_16 = r_lvl_output_ff_144; // @[FanNetwork.scala 1650:23]
  assign io_o_data_bus_17 = r_lvl_output_ff_145; // @[FanNetwork.scala 1651:23]
  assign io_o_data_bus_18 = r_lvl_output_ff_146; // @[FanNetwork.scala 1652:23]
  assign io_o_data_bus_19 = r_lvl_output_ff_147; // @[FanNetwork.scala 1653:23]
  assign io_o_data_bus_20 = r_lvl_output_ff_148; // @[FanNetwork.scala 1654:23]
  assign io_o_data_bus_21 = r_lvl_output_ff_149; // @[FanNetwork.scala 1655:23]
  assign io_o_data_bus_22 = r_lvl_output_ff_150; // @[FanNetwork.scala 1656:23]
  assign io_o_data_bus_23 = r_lvl_output_ff_151; // @[FanNetwork.scala 1657:23]
  assign io_o_data_bus_24 = r_lvl_output_ff_152; // @[FanNetwork.scala 1658:23]
  assign io_o_data_bus_25 = r_lvl_output_ff_153; // @[FanNetwork.scala 1659:23]
  assign io_o_data_bus_26 = r_lvl_output_ff_154; // @[FanNetwork.scala 1660:23]
  assign io_o_data_bus_27 = r_lvl_output_ff_155; // @[FanNetwork.scala 1661:23]
  assign io_o_data_bus_28 = r_lvl_output_ff_156; // @[FanNetwork.scala 1662:23]
  assign io_o_data_bus_29 = r_lvl_output_ff_157; // @[FanNetwork.scala 1663:23]
  assign io_o_data_bus_30 = r_lvl_output_ff_158; // @[FanNetwork.scala 1664:23]
  assign io_o_data_bus_31 = r_lvl_output_ff_159; // @[FanNetwork.scala 1665:23]
  assign my_adder_0_clock = clock;
  assign my_adder_0_reset = reset;
  assign my_adder_0_io_i_valid = r_valid_0; // @[FanNetwork.scala 1020:27]
  assign my_adder_0_io_i_data_bus_0 = {{32'd0}, io_i_data_bus_1}; // @[FanNetwork.scala 1021:30]
  assign my_adder_0_io_i_data_bus_1 = {{32'd0}, io_i_data_bus_0}; // @[FanNetwork.scala 1021:30]
  assign my_adder_0_io_i_add_en = {{2'd0}, io_i_add_en_bus_0}; // @[FanNetwork.scala 1022:28]
  assign my_adder_0_io_i_cmd = {{2'd0}, io_i_cmd_bus_0}; // @[FanNetwork.scala 1023:25]
  assign my_adder_1_clock = clock;
  assign my_adder_1_reset = reset;
  assign my_adder_1_io_i_valid = r_valid_1; // @[FanNetwork.scala 1033:27]
  assign my_adder_1_io_i_data_bus_0 = w_fan_lvl_0_1[63:0]; // @[FanNetwork.scala 1034:30]
  assign my_adder_1_io_i_data_bus_1 = w_fan_lvl_0_0[63:0]; // @[FanNetwork.scala 1034:30]
  assign my_adder_1_io_i_add_en = {{2'd0}, io_i_add_en_bus_16}; // @[FanNetwork.scala 1035:28]
  assign my_adder_1_io_i_cmd = {{2'd0}, io_i_cmd_bus_16}; // @[FanNetwork.scala 1037:26]
  assign my_adder_2_clock = clock;
  assign my_adder_2_reset = reset;
  assign my_adder_2_io_i_valid = r_valid_0; // @[FanNetwork.scala 1047:27]
  assign my_adder_2_io_i_data_bus_0 = io_i_data_bus_3; // @[FanNetwork.scala 1048:{40,40}]
  assign my_adder_2_io_i_data_bus_1 = io_i_data_bus_2; // @[FanNetwork.scala 1048:{40,40}]
  assign my_adder_2_io_i_add_en = {{2'd0}, io_i_add_en_bus_1}; // @[FanNetwork.scala 1049:28]
  assign my_adder_2_io_i_cmd = io_i_cmd_bus_1; // @[FanNetwork.scala 1051:25]
  assign my_adder_3_clock = clock;
  assign my_adder_3_reset = reset;
  assign my_adder_3_io_i_valid = r_valid_2; // @[FanNetwork.scala 1066:27]
  assign my_adder_3_io_i_data_bus_0 = w_fan_lvl_1_1[63:0]; // @[FanNetwork.scala 1067:32]
  assign my_adder_3_io_i_data_bus_1 = _WIRE_9_1[63:0]; // @[FanNetwork.scala 1067:32]
  assign my_adder_3_io_i_data_bus_2 = _WIRE_9_2[63:0]; // @[FanNetwork.scala 1067:32]
  assign my_adder_3_io_i_data_bus_3 = w_fan_lvl_1_0[63:0]; // @[FanNetwork.scala 1067:32]
  assign my_adder_3_io_i_add_en = {{2'd0}, io_i_add_en_bus_24}; // @[FanNetwork.scala 1069:28]
  assign my_adder_3_io_i_cmd = {{2'd0}, io_i_cmd_bus_24}; // @[FanNetwork.scala 1071:27]
  assign my_adder_3_io_i_sel = {{1'd0}, io_i_sel_bus_1}; // @[FanNetwork.scala 1072:25]
  assign my_adder_4_clock = clock;
  assign my_adder_4_reset = reset;
  assign my_adder_4_io_i_valid = r_valid_0; // @[FanNetwork.scala 1083:27]
  assign my_adder_4_io_i_data_bus_0 = io_i_data_bus_5; // @[FanNetwork.scala 1084:{40,40}]
  assign my_adder_4_io_i_data_bus_1 = io_i_data_bus_4; // @[FanNetwork.scala 1084:{40,40}]
  assign my_adder_4_io_i_add_en = {{2'd0}, io_i_add_en_bus_2}; // @[FanNetwork.scala 1085:28]
  assign my_adder_4_io_i_cmd = io_i_cmd_bus_2; // @[FanNetwork.scala 1086:26]
  assign my_adder_5_clock = clock;
  assign my_adder_5_reset = reset;
  assign my_adder_5_io_i_valid = r_valid_1; // @[FanNetwork.scala 1101:27]
  assign my_adder_5_io_i_data_bus_0 = w_fan_lvl_0_5[31:0]; // @[FanNetwork.scala 1102:30]
  assign my_adder_5_io_i_data_bus_1 = w_fan_lvl_0_4[31:0]; // @[FanNetwork.scala 1102:30]
  assign my_adder_5_io_i_add_en = {{2'd0}, io_i_add_en_bus_17}; // @[FanNetwork.scala 1103:28]
  assign my_adder_5_io_i_cmd = io_i_cmd_bus_17; // @[FanNetwork.scala 1105:26]
  assign my_adder_6_clock = clock;
  assign my_adder_6_reset = reset;
  assign my_adder_6_io_i_valid = r_valid_0; // @[FanNetwork.scala 1118:27]
  assign my_adder_6_io_i_data_bus_0 = io_i_data_bus_7; // @[FanNetwork.scala 1119:{40,40}]
  assign my_adder_6_io_i_data_bus_1 = io_i_data_bus_6; // @[FanNetwork.scala 1119:{40,40}]
  assign my_adder_6_io_i_add_en = {{2'd0}, io_i_add_en_bus_3}; // @[FanNetwork.scala 1120:28]
  assign my_adder_6_io_i_cmd = io_i_cmd_bus_3; // @[FanNetwork.scala 1121:25]
  assign my_adder_7_clock = clock;
  assign my_adder_7_reset = reset;
  assign my_adder_7_io_i_valid = r_valid_3; // @[FanNetwork.scala 1135:27]
  assign my_adder_7_io_i_data_bus_0 = w_fan_lvl_2_1[63:0]; // @[FanNetwork.scala 1138:30]
  assign my_adder_7_io_i_data_bus_1 = _WIRE_13_1[63:0]; // @[FanNetwork.scala 1138:30]
  assign my_adder_7_io_i_data_bus_2 = _WIRE_13_2[63:0]; // @[FanNetwork.scala 1138:30]
  assign my_adder_7_io_i_data_bus_3 = _WIRE_13_3[63:0]; // @[FanNetwork.scala 1138:30]
  assign my_adder_7_io_i_data_bus_4 = _WIRE_13_4[63:0]; // @[FanNetwork.scala 1138:30]
  assign my_adder_7_io_i_data_bus_5 = w_fan_lvl_2_0[63:0]; // @[FanNetwork.scala 1138:30]
  assign my_adder_7_io_i_add_en = {{2'd0}, io_i_add_en_bus_28}; // @[FanNetwork.scala 1139:28]
  assign my_adder_7_io_i_cmd = {{2'd0}, io_i_cmd_bus_28}; // @[FanNetwork.scala 1141:25]
  assign my_adder_7_io_i_sel = {my_adder_7_io_i_sel_hi,my_adder_7_io_i_sel_lo}; // @[Cat.scala 33:92]
  assign my_adder_8_clock = clock;
  assign my_adder_8_reset = reset;
  assign my_adder_8_io_i_valid = r_valid_0; // @[FanNetwork.scala 1154:27]
  assign my_adder_8_io_i_data_bus_0 = io_i_data_bus_9; // @[FanNetwork.scala 1155:{40,40}]
  assign my_adder_8_io_i_data_bus_1 = io_i_data_bus_8; // @[FanNetwork.scala 1155:{40,40}]
  assign my_adder_8_io_i_add_en = {{2'd0}, io_i_add_en_bus_4}; // @[FanNetwork.scala 1156:28]
  assign my_adder_8_io_i_cmd = io_i_cmd_bus_4; // @[FanNetwork.scala 1158:25]
  assign my_adder_9_clock = clock;
  assign my_adder_9_reset = reset;
  assign my_adder_9_io_i_valid = r_valid_1; // @[FanNetwork.scala 1171:27]
  assign my_adder_9_io_i_data_bus_0 = w_fan_lvl_0_9[31:0]; // @[FanNetwork.scala 1172:30]
  assign my_adder_9_io_i_data_bus_1 = w_fan_lvl_0_8[31:0]; // @[FanNetwork.scala 1172:30]
  assign my_adder_9_io_i_add_en = {{2'd0}, io_i_add_en_bus_18}; // @[FanNetwork.scala 1173:28]
  assign my_adder_9_io_i_cmd = io_i_cmd_bus_18; // @[FanNetwork.scala 1175:25]
  assign my_adder_10_clock = clock;
  assign my_adder_10_reset = reset;
  assign my_adder_10_io_i_valid = r_valid_0; // @[FanNetwork.scala 1188:28]
  assign my_adder_10_io_i_data_bus_0 = io_i_data_bus_11; // @[FanNetwork.scala 1189:{41,41}]
  assign my_adder_10_io_i_data_bus_1 = io_i_data_bus_10; // @[FanNetwork.scala 1189:{41,41}]
  assign my_adder_10_io_i_add_en = {{2'd0}, io_i_add_en_bus_5}; // @[FanNetwork.scala 1190:29]
  assign my_adder_10_io_i_cmd = io_i_cmd_bus_5; // @[FanNetwork.scala 1191:27]
  assign my_adder_11_clock = clock;
  assign my_adder_11_reset = reset;
  assign my_adder_11_io_i_valid = r_valid_2; // @[FanNetwork.scala 1206:28]
  assign my_adder_11_io_i_data_bus_0 = w_fan_lvl_1_5[31:0]; // @[FanNetwork.scala 1208:31]
  assign my_adder_11_io_i_data_bus_1 = _WIRE_17_1[31:0]; // @[FanNetwork.scala 1208:31]
  assign my_adder_11_io_i_data_bus_2 = _WIRE_17_2[31:0]; // @[FanNetwork.scala 1208:31]
  assign my_adder_11_io_i_data_bus_3 = w_fan_lvl_1_4[31:0]; // @[FanNetwork.scala 1208:31]
  assign my_adder_11_io_i_add_en = {{2'd0}, io_i_add_en_bus_25}; // @[FanNetwork.scala 1210:29]
  assign my_adder_11_io_i_cmd = io_i_cmd_bus_25; // @[FanNetwork.scala 1212:26]
  assign my_adder_11_io_i_sel = {io_i_sel_bus_3,io_i_sel_bus_2}; // @[Cat.scala 33:92]
  assign my_adder_12_clock = clock;
  assign my_adder_12_reset = reset;
  assign my_adder_12_io_i_valid = r_valid_0; // @[FanNetwork.scala 1227:28]
  assign my_adder_12_io_i_data_bus_0 = io_i_data_bus_13; // @[FanNetwork.scala 1228:{41,41}]
  assign my_adder_12_io_i_data_bus_1 = io_i_data_bus_12; // @[FanNetwork.scala 1228:{41,41}]
  assign my_adder_12_io_i_add_en = {{2'd0}, io_i_add_en_bus_6}; // @[FanNetwork.scala 1229:29]
  assign my_adder_12_io_i_cmd = io_i_cmd_bus_6; // @[FanNetwork.scala 1231:27]
  assign my_adder_13_clock = clock;
  assign my_adder_13_reset = reset;
  assign my_adder_13_io_i_valid = r_valid_1; // @[FanNetwork.scala 1245:28]
  assign my_adder_13_io_i_data_bus_0 = w_fan_lvl_0_12[31:0]; // @[FanNetwork.scala 1246:31]
  assign my_adder_13_io_i_data_bus_1 = w_fan_lvl_0_11[31:0]; // @[FanNetwork.scala 1246:31]
  assign my_adder_13_io_i_add_en = {{2'd0}, io_i_add_en_bus_19}; // @[FanNetwork.scala 1247:29]
  assign my_adder_13_io_i_cmd = io_i_cmd_bus_19; // @[FanNetwork.scala 1249:26]
  assign my_adder_14_clock = clock;
  assign my_adder_14_reset = reset;
  assign my_adder_14_io_i_valid = r_valid_0; // @[FanNetwork.scala 1263:28]
  assign my_adder_14_io_i_data_bus_0 = io_i_data_bus_15; // @[FanNetwork.scala 1264:{41,41}]
  assign my_adder_14_io_i_data_bus_1 = io_i_data_bus_14; // @[FanNetwork.scala 1264:{41,41}]
  assign my_adder_14_io_i_add_en = {{2'd0}, io_i_add_en_bus_7}; // @[FanNetwork.scala 1265:29]
  assign my_adder_14_io_i_cmd = io_i_cmd_bus_7; // @[FanNetwork.scala 1267:26]
  assign my_adder_15_clock = clock;
  assign my_adder_15_reset = reset;
  assign my_adder_15_io_i_valid = r_valid_4; // @[FanNetwork.scala 1281:28]
  assign my_adder_15_io_i_data_bus_0 = {{32'd0}, my_adder_23_io_o_adder}; // @[FanNetwork.scala 1283:{41,41}]
  assign my_adder_15_io_i_data_bus_1 = {{32'd0}, r_fan_ff_lvl_2_to_4_1}; // @[FanNetwork.scala 1283:{41,41}]
  assign my_adder_15_io_i_data_bus_2 = {{32'd0}, r_fan_ff_lvl_1_to_4_1}; // @[FanNetwork.scala 1283:{41,41}]
  assign my_adder_15_io_i_data_bus_3 = {{32'd0}, r_fan_ff_lvl_0_to_4_1}; // @[FanNetwork.scala 1283:{41,41}]
  assign my_adder_15_io_i_data_bus_4 = {{32'd0}, r_fan_ff_lvl_0_to_4_0}; // @[FanNetwork.scala 1283:{41,41}]
  assign my_adder_15_io_i_data_bus_5 = {{32'd0}, r_fan_ff_lvl_1_to_4_0}; // @[FanNetwork.scala 1283:{41,41}]
  assign my_adder_15_io_i_data_bus_6 = {{32'd0}, r_fan_ff_lvl_2_to_4_0}; // @[FanNetwork.scala 1283:{41,41}]
  assign my_adder_15_io_i_data_bus_7 = {{32'd0}, my_adder_7_io_o_adder}; // @[FanNetwork.scala 1283:{41,41}]
  assign my_adder_15_io_i_add_en = {{2'd0}, io_i_add_en_bus_30}; // @[FanNetwork.scala 1285:29]
  assign my_adder_15_io_i_cmd = {{2'd0}, io_i_cmd_bus_30}; // @[FanNetwork.scala 1287:26]
  assign my_adder_15_io_i_sel = {{2'd0}, _my_adder_15_io_i_sel_T}; // @[FanNetwork.scala 1288:26]
  assign my_adder_16_clock = clock;
  assign my_adder_16_reset = reset;
  assign my_adder_16_io_i_valid = r_valid_0; // @[FanNetwork.scala 1301:28]
  assign my_adder_16_io_i_data_bus_0 = io_i_data_bus_17; // @[FanNetwork.scala 1302:{41,41}]
  assign my_adder_16_io_i_data_bus_1 = io_i_data_bus_16; // @[FanNetwork.scala 1302:{41,41}]
  assign my_adder_16_io_i_add_en = {{2'd0}, io_i_add_en_bus_8}; // @[FanNetwork.scala 1303:29]
  assign my_adder_16_io_i_cmd = io_i_cmd_bus_8; // @[FanNetwork.scala 1305:26]
  assign my_adder_17_clock = clock;
  assign my_adder_17_reset = reset;
  assign my_adder_17_io_i_valid = r_valid_1; // @[FanNetwork.scala 1319:28]
  assign my_adder_17_io_i_data_bus_0 = w_fan_lvl_0_16[31:0]; // @[FanNetwork.scala 1320:31]
  assign my_adder_17_io_i_data_bus_1 = w_fan_lvl_0_15[31:0]; // @[FanNetwork.scala 1320:31]
  assign my_adder_17_io_i_add_en = {{2'd0}, io_i_add_en_bus_20}; // @[FanNetwork.scala 1321:29]
  assign my_adder_17_io_i_cmd = io_i_cmd_bus_20; // @[FanNetwork.scala 1322:26]
  assign my_adder_18_clock = clock;
  assign my_adder_18_reset = reset;
  assign my_adder_18_io_i_valid = r_valid_0; // @[FanNetwork.scala 1337:28]
  assign my_adder_18_io_i_data_bus_0 = io_i_data_bus_19; // @[FanNetwork.scala 1338:{41,41}]
  assign my_adder_18_io_i_data_bus_1 = io_i_data_bus_18; // @[FanNetwork.scala 1338:{41,41}]
  assign my_adder_18_io_i_add_en = {{2'd0}, io_i_add_en_bus_9}; // @[FanNetwork.scala 1339:29]
  assign my_adder_18_io_i_cmd = io_i_cmd_bus_9; // @[FanNetwork.scala 1341:26]
  assign my_adder_19_clock = clock;
  assign my_adder_19_reset = reset;
  assign my_adder_19_io_i_valid = r_valid_2; // @[FanNetwork.scala 1355:28]
  assign my_adder_19_io_i_data_bus_0 = w_fan_lvl_1_9[31:0]; // @[FanNetwork.scala 1357:32]
  assign my_adder_19_io_i_data_bus_1 = _WIRE_25_1[31:0]; // @[FanNetwork.scala 1357:32]
  assign my_adder_19_io_i_data_bus_2 = _WIRE_25_2[31:0]; // @[FanNetwork.scala 1357:32]
  assign my_adder_19_io_i_data_bus_3 = w_fan_lvl_1_8[31:0]; // @[FanNetwork.scala 1357:32]
  assign my_adder_19_io_i_add_en = {{2'd0}, io_i_add_en_bus_26}; // @[FanNetwork.scala 1358:29]
  assign my_adder_19_io_i_cmd = io_i_cmd_bus_26; // @[FanNetwork.scala 1359:26]
  assign my_adder_19_io_i_sel = {io_i_sel_bus_5,io_i_sel_bus_4}; // @[Cat.scala 33:92]
  assign my_adder_20_clock = clock;
  assign my_adder_20_reset = reset;
  assign my_adder_20_io_i_valid = r_valid_0; // @[FanNetwork.scala 1375:28]
  assign my_adder_20_io_i_data_bus_0 = io_i_data_bus_21; // @[FanNetwork.scala 1376:{41,41}]
  assign my_adder_20_io_i_data_bus_1 = io_i_data_bus_20; // @[FanNetwork.scala 1376:{41,41}]
  assign my_adder_20_io_i_add_en = {{2'd0}, io_i_add_en_bus_10}; // @[FanNetwork.scala 1377:29]
  assign my_adder_20_io_i_cmd = io_i_cmd_bus_10; // @[FanNetwork.scala 1379:26]
  assign my_adder_21_clock = clock;
  assign my_adder_21_reset = reset;
  assign my_adder_21_io_i_valid = r_valid_1; // @[FanNetwork.scala 1395:28]
  assign my_adder_21_io_i_data_bus_0 = w_fan_lvl_0_20[31:0]; // @[FanNetwork.scala 1396:31]
  assign my_adder_21_io_i_data_bus_1 = w_fan_lvl_0_19[31:0]; // @[FanNetwork.scala 1396:31]
  assign my_adder_21_io_i_add_en = {{2'd0}, io_i_add_en_bus_21}; // @[FanNetwork.scala 1397:29]
  assign my_adder_21_io_i_cmd = io_i_cmd_bus_21; // @[FanNetwork.scala 1398:27]
  assign my_adder_22_clock = clock;
  assign my_adder_22_reset = reset;
  assign my_adder_22_io_i_valid = r_valid_0; // @[FanNetwork.scala 1414:28]
  assign my_adder_22_io_i_data_bus_0 = io_i_data_bus_23; // @[FanNetwork.scala 1415:{41,41}]
  assign my_adder_22_io_i_data_bus_1 = io_i_data_bus_22; // @[FanNetwork.scala 1415:{41,41}]
  assign my_adder_22_io_i_add_en = {{2'd0}, io_i_add_en_bus_11}; // @[FanNetwork.scala 1416:29]
  assign my_adder_22_io_i_cmd = io_i_cmd_bus_11; // @[FanNetwork.scala 1417:26]
  assign my_adder_23_clock = clock;
  assign my_adder_23_reset = reset;
  assign my_adder_23_io_i_valid = r_valid_3; // @[FanNetwork.scala 1432:28]
  assign my_adder_23_io_i_data_bus_0 = w_fan_lvl_2_5[63:0]; // @[FanNetwork.scala 1434:31]
  assign my_adder_23_io_i_data_bus_1 = _WIRE_29_1[63:0]; // @[FanNetwork.scala 1434:31]
  assign my_adder_23_io_i_data_bus_2 = _WIRE_29_2[63:0]; // @[FanNetwork.scala 1434:31]
  assign my_adder_23_io_i_data_bus_3 = _WIRE_29_3[63:0]; // @[FanNetwork.scala 1434:31]
  assign my_adder_23_io_i_data_bus_4 = _WIRE_29_4[63:0]; // @[FanNetwork.scala 1434:31]
  assign my_adder_23_io_i_data_bus_5 = w_fan_lvl_2_4[63:0]; // @[FanNetwork.scala 1434:31]
  assign my_adder_23_io_i_add_en = {{2'd0}, io_i_add_en_bus_29}; // @[FanNetwork.scala 1435:29]
  assign my_adder_23_io_i_cmd = {{2'd0}, io_i_cmd_bus_29}; // @[FanNetwork.scala 1437:26]
  assign my_adder_23_io_i_sel = {{2'd0}, _my_adder_23_io_i_sel_T}; // @[FanNetwork.scala 1438:26]
  assign my_adder_24_clock = clock;
  assign my_adder_24_reset = reset;
  assign my_adder_24_io_i_valid = r_valid_0; // @[FanNetwork.scala 1449:28]
  assign my_adder_24_io_i_data_bus_0 = io_i_data_bus_25; // @[FanNetwork.scala 1450:{41,41}]
  assign my_adder_24_io_i_data_bus_1 = io_i_data_bus_24; // @[FanNetwork.scala 1450:{41,41}]
  assign my_adder_24_io_i_add_en = {{2'd0}, io_i_add_en_bus_12}; // @[FanNetwork.scala 1451:29]
  assign my_adder_24_io_i_cmd = io_i_cmd_bus_12; // @[FanNetwork.scala 1453:26]
  assign my_adder_25_clock = clock;
  assign my_adder_25_reset = reset;
  assign my_adder_25_io_i_valid = r_valid_1; // @[FanNetwork.scala 1468:28]
  assign my_adder_25_io_i_data_bus_0 = w_fan_lvl_0_24[31:0]; // @[FanNetwork.scala 1469:31]
  assign my_adder_25_io_i_data_bus_1 = w_fan_lvl_0_23[31:0]; // @[FanNetwork.scala 1469:31]
  assign my_adder_25_io_i_add_en = {{2'd0}, io_i_add_en_bus_22}; // @[FanNetwork.scala 1470:29]
  assign my_adder_25_io_i_cmd = io_i_cmd_bus_22; // @[FanNetwork.scala 1472:26]
  assign my_adder_26_clock = clock;
  assign my_adder_26_reset = reset;
  assign my_adder_26_io_i_valid = r_valid_0; // @[FanNetwork.scala 1488:28]
  assign my_adder_26_io_i_data_bus_0 = io_i_data_bus_27; // @[FanNetwork.scala 1489:{41,41}]
  assign my_adder_26_io_i_data_bus_1 = io_i_data_bus_26; // @[FanNetwork.scala 1489:{41,41}]
  assign my_adder_26_io_i_add_en = {{2'd0}, io_i_add_en_bus_13}; // @[FanNetwork.scala 1490:29]
  assign my_adder_26_io_i_cmd = io_i_cmd_bus_13; // @[FanNetwork.scala 1491:26]
  assign my_adder_27_clock = clock;
  assign my_adder_27_reset = reset;
  assign my_adder_27_io_i_valid = r_valid_2; // @[FanNetwork.scala 1506:28]
  assign my_adder_27_io_i_data_bus_0 = w_fan_lvl_1_13[63:0]; // @[FanNetwork.scala 1508:31]
  assign my_adder_27_io_i_data_bus_1 = _WIRE_33_1[63:0]; // @[FanNetwork.scala 1508:31]
  assign my_adder_27_io_i_data_bus_2 = _WIRE_33_2[63:0]; // @[FanNetwork.scala 1508:31]
  assign my_adder_27_io_i_data_bus_3 = w_fan_lvl_1_12[63:0]; // @[FanNetwork.scala 1508:31]
  assign my_adder_27_io_i_add_en = {{2'd0}, io_i_add_en_bus_27}; // @[FanNetwork.scala 1509:29]
  assign my_adder_27_io_i_cmd = {{2'd0}, io_i_cmd_bus_27}; // @[FanNetwork.scala 1511:26]
  assign my_adder_27_io_i_sel = {io_i_sel_bus_7,io_i_sel_bus_6}; // @[Cat.scala 33:92]
  assign my_adder_28_clock = clock;
  assign my_adder_28_reset = reset;
  assign my_adder_28_io_i_valid = r_valid_0; // @[FanNetwork.scala 1527:28]
  assign my_adder_28_io_i_data_bus_0 = io_i_data_bus_29; // @[FanNetwork.scala 1528:{41,41}]
  assign my_adder_28_io_i_data_bus_1 = io_i_data_bus_28; // @[FanNetwork.scala 1528:{41,41}]
  assign my_adder_28_io_i_add_en = {{2'd0}, io_i_add_en_bus_14}; // @[FanNetwork.scala 1529:29]
  assign my_adder_28_io_i_cmd = io_i_cmd_bus_14; // @[FanNetwork.scala 1531:27]
  assign my_adder_29_clock = clock;
  assign my_adder_29_reset = reset;
  assign my_adder_29_io_i_valid = r_valid_1; // @[FanNetwork.scala 1546:28]
  assign my_adder_29_io_i_data_bus_0 = w_fan_lvl_0_28[63:0]; // @[FanNetwork.scala 1547:31]
  assign my_adder_29_io_i_data_bus_1 = w_fan_lvl_0_27[63:0]; // @[FanNetwork.scala 1547:31]
  assign my_adder_29_io_i_add_en = {{2'd0}, io_i_add_en_bus_23}; // @[FanNetwork.scala 1548:29]
  assign my_adder_29_io_i_cmd = {{2'd0}, io_i_cmd_bus_23}; // @[FanNetwork.scala 1550:26]
  assign my_adder_30_clock = clock;
  assign my_adder_30_reset = reset;
  assign my_adder_30_io_i_valid = r_valid_0; // @[FanNetwork.scala 1564:28]
  assign my_adder_30_io_i_data_bus_0 = {{32'd0}, io_i_data_bus_31}; // @[FanNetwork.scala 1565:31]
  assign my_adder_30_io_i_data_bus_1 = {{32'd0}, io_i_data_bus_30}; // @[FanNetwork.scala 1565:31]
  assign my_adder_30_io_i_add_en = {{2'd0}, io_i_add_en_bus_15}; // @[FanNetwork.scala 1566:29]
  assign my_adder_30_io_i_cmd = {{2'd0}, io_i_cmd_bus_15}; // @[FanNetwork.scala 1568:26]
  always @(posedge clock) begin
    if (reset) begin // @[FanNetwork.scala 32:38]
      r_fan_ff_lvl_0_to_4_0 <= 32'h0; // @[FanNetwork.scala 32:38]
    end else begin
      r_fan_ff_lvl_0_to_4_0 <= r_fan_ff_lvl_0_to_3_2; // @[FanNetwork.scala 75:25]
    end
    if (reset) begin // @[FanNetwork.scala 32:38]
      r_fan_ff_lvl_0_to_4_1 <= 32'h0; // @[FanNetwork.scala 32:38]
    end else begin
      r_fan_ff_lvl_0_to_4_1 <= r_fan_ff_lvl_0_to_3_3; // @[FanNetwork.scala 75:25]
    end
    if (reset) begin // @[FanNetwork.scala 33:38]
      r_fan_ff_lvl_0_to_3_0 <= 32'h0; // @[FanNetwork.scala 33:38]
    end else begin
      r_fan_ff_lvl_0_to_3_0 <= r_fan_ff_lvl_0_to_2_2; // @[FanNetwork.scala 74:25]
    end
    if (reset) begin // @[FanNetwork.scala 33:38]
      r_fan_ff_lvl_0_to_3_1 <= 32'h0; // @[FanNetwork.scala 33:38]
    end else begin
      r_fan_ff_lvl_0_to_3_1 <= r_fan_ff_lvl_0_to_2_3; // @[FanNetwork.scala 74:25]
    end
    if (reset) begin // @[FanNetwork.scala 33:38]
      r_fan_ff_lvl_0_to_3_2 <= 32'h0; // @[FanNetwork.scala 33:38]
    end else begin
      r_fan_ff_lvl_0_to_3_2 <= r_fan_ff_lvl_0_to_2_6; // @[FanNetwork.scala 74:25]
    end
    if (reset) begin // @[FanNetwork.scala 33:38]
      r_fan_ff_lvl_0_to_3_3 <= 32'h0; // @[FanNetwork.scala 33:38]
    end else begin
      r_fan_ff_lvl_0_to_3_3 <= r_fan_ff_lvl_0_to_2_7; // @[FanNetwork.scala 74:25]
    end
    if (reset) begin // @[FanNetwork.scala 33:38]
      r_fan_ff_lvl_0_to_3_4 <= 32'h0; // @[FanNetwork.scala 33:38]
    end else begin
      r_fan_ff_lvl_0_to_3_4 <= r_fan_ff_lvl_0_to_2_10; // @[FanNetwork.scala 74:25]
    end
    if (reset) begin // @[FanNetwork.scala 33:38]
      r_fan_ff_lvl_0_to_3_5 <= 32'h0; // @[FanNetwork.scala 33:38]
    end else begin
      r_fan_ff_lvl_0_to_3_5 <= r_fan_ff_lvl_0_to_2_11; // @[FanNetwork.scala 74:25]
    end
    r_fan_ff_lvl_0_to_2_0 <= _GEN_239[31:0]; // @[FanNetwork.scala 34:{38,38} 73:25]
    r_fan_ff_lvl_0_to_2_1 <= _GEN_240[31:0]; // @[FanNetwork.scala 34:{38,38} 73:25]
    r_fan_ff_lvl_0_to_2_2 <= _GEN_241[31:0]; // @[FanNetwork.scala 34:{38,38} 73:25]
    r_fan_ff_lvl_0_to_2_3 <= _GEN_242[31:0]; // @[FanNetwork.scala 34:{38,38} 73:25]
    r_fan_ff_lvl_0_to_2_4 <= _GEN_243[31:0]; // @[FanNetwork.scala 34:{38,38} 73:25]
    r_fan_ff_lvl_0_to_2_5 <= _GEN_244[31:0]; // @[FanNetwork.scala 34:{38,38} 73:25]
    r_fan_ff_lvl_0_to_2_6 <= _GEN_245[31:0]; // @[FanNetwork.scala 34:{38,38} 73:25]
    r_fan_ff_lvl_0_to_2_7 <= _GEN_246[31:0]; // @[FanNetwork.scala 34:{38,38} 73:25]
    r_fan_ff_lvl_0_to_2_8 <= _GEN_247[31:0]; // @[FanNetwork.scala 34:{38,38} 73:25]
    r_fan_ff_lvl_0_to_2_9 <= _GEN_248[31:0]; // @[FanNetwork.scala 34:{38,38} 73:25]
    r_fan_ff_lvl_0_to_2_10 <= _GEN_249[31:0]; // @[FanNetwork.scala 34:{38,38} 73:25]
    r_fan_ff_lvl_0_to_2_11 <= _GEN_250[31:0]; // @[FanNetwork.scala 34:{38,38} 73:25]
    r_fan_ff_lvl_0_to_2_12 <= _GEN_251[31:0]; // @[FanNetwork.scala 34:{38,38} 73:25]
    r_fan_ff_lvl_0_to_2_13 <= _GEN_252[31:0]; // @[FanNetwork.scala 34:{38,38} 73:25]
    if (reset) begin // @[FanNetwork.scala 35:38]
      r_fan_ff_lvl_1_to_4_0 <= 32'h0; // @[FanNetwork.scala 35:38]
    end else begin
      r_fan_ff_lvl_1_to_4_0 <= r_fan_ff_lvl_1_to_3_2; // @[FanNetwork.scala 76:25]
    end
    if (reset) begin // @[FanNetwork.scala 35:38]
      r_fan_ff_lvl_1_to_4_1 <= 32'h0; // @[FanNetwork.scala 35:38]
    end else begin
      r_fan_ff_lvl_1_to_4_1 <= r_fan_ff_lvl_1_to_3_3; // @[FanNetwork.scala 76:25]
    end
    r_fan_ff_lvl_1_to_3_0 <= _GEN_253[31:0]; // @[FanNetwork.scala 36:{38,38} 77:25]
    r_fan_ff_lvl_1_to_3_1 <= _GEN_254[31:0]; // @[FanNetwork.scala 36:{38,38} 77:25]
    r_fan_ff_lvl_1_to_3_2 <= _GEN_255[31:0]; // @[FanNetwork.scala 36:{38,38} 77:25]
    r_fan_ff_lvl_1_to_3_3 <= _GEN_256[31:0]; // @[FanNetwork.scala 36:{38,38} 77:25]
    r_fan_ff_lvl_1_to_3_4 <= _GEN_257[31:0]; // @[FanNetwork.scala 36:{38,38} 77:25]
    r_fan_ff_lvl_1_to_3_5 <= _GEN_258[31:0]; // @[FanNetwork.scala 36:{38,38} 77:25]
    r_fan_ff_lvl_2_to_4_0 <= _GEN_259[31:0]; // @[FanNetwork.scala 37:{38,38} 78:25]
    r_fan_ff_lvl_2_to_4_1 <= _GEN_260[31:0]; // @[FanNetwork.scala 37:{38,38} 78:25]
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_0 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_0_valid_1 & w_vn_lvl_0_valid_0) begin // @[FanNetwork.scala 83:77]
      r_lvl_output_ff_0 <= w_vn_lvl_0_0; // @[FanNetwork.scala 85:24]
    end else if (w_vn_lvl_0_valid_1 & ~w_vn_lvl_0_valid_0) begin // @[FanNetwork.scala 88:83]
      r_lvl_output_ff_0 <= 32'h0; // @[FanNetwork.scala 90:24]
    end else if (~w_vn_lvl_0_valid_1 & w_vn_lvl_0_valid_0) begin // @[FanNetwork.scala 93:83]
      r_lvl_output_ff_0 <= w_vn_lvl_0_0; // @[FanNetwork.scala 95:24]
    end else begin
      r_lvl_output_ff_0 <= 32'h0; // @[FanNetwork.scala 100:24]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_1 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_0_valid_1 & w_vn_lvl_0_valid_0) begin // @[FanNetwork.scala 83:77]
      r_lvl_output_ff_1 <= w_vn_lvl_0_1; // @[FanNetwork.scala 84:24]
    end else if (w_vn_lvl_0_valid_1 & ~w_vn_lvl_0_valid_0) begin // @[FanNetwork.scala 88:83]
      r_lvl_output_ff_1 <= w_vn_lvl_0_1; // @[FanNetwork.scala 89:24]
    end else begin
      r_lvl_output_ff_1 <= 32'h0;
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_2 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_0_valid_3 & w_vn_lvl_0_valid_2) begin // @[FanNetwork.scala 106:77]
      r_lvl_output_ff_2 <= w_vn_lvl_0_2; // @[FanNetwork.scala 108:24]
    end else if (w_vn_lvl_0_valid_3 & ~w_vn_lvl_0_valid_2) begin // @[FanNetwork.scala 111:83]
      r_lvl_output_ff_2 <= 32'h0; // @[FanNetwork.scala 113:24]
    end else if (~w_vn_lvl_0_valid_3 & w_vn_lvl_0_valid_2) begin // @[FanNetwork.scala 116:83]
      r_lvl_output_ff_2 <= w_vn_lvl_0_2; // @[FanNetwork.scala 118:24]
    end else begin
      r_lvl_output_ff_2 <= 32'h0; // @[FanNetwork.scala 123:24]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_3 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_0_valid_3 & w_vn_lvl_0_valid_2) begin // @[FanNetwork.scala 106:77]
      r_lvl_output_ff_3 <= w_vn_lvl_0_3; // @[FanNetwork.scala 107:24]
    end else if (w_vn_lvl_0_valid_3 & ~w_vn_lvl_0_valid_2) begin // @[FanNetwork.scala 111:83]
      r_lvl_output_ff_3 <= w_vn_lvl_0_3; // @[FanNetwork.scala 112:24]
    end else begin
      r_lvl_output_ff_3 <= 32'h0;
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_6 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_0_valid_7 & w_vn_lvl_0_valid_6) begin // @[FanNetwork.scala 151:77]
      r_lvl_output_ff_6 <= w_vn_lvl_0_6; // @[FanNetwork.scala 153:24]
    end else if (w_vn_lvl_0_valid_7 & ~w_vn_lvl_0_valid_6) begin // @[FanNetwork.scala 156:83]
      r_lvl_output_ff_6 <= 32'h0; // @[FanNetwork.scala 158:24]
    end else if (~w_vn_lvl_0_valid_7 & w_vn_lvl_0_valid_6) begin // @[FanNetwork.scala 161:83]
      r_lvl_output_ff_6 <= w_vn_lvl_0_6; // @[FanNetwork.scala 163:24]
    end else begin
      r_lvl_output_ff_6 <= 32'h0; // @[FanNetwork.scala 168:24]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_7 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_0_valid_7 & w_vn_lvl_0_valid_6) begin // @[FanNetwork.scala 151:77]
      r_lvl_output_ff_7 <= w_vn_lvl_0_7; // @[FanNetwork.scala 152:24]
    end else if (w_vn_lvl_0_valid_7 & ~w_vn_lvl_0_valid_6) begin // @[FanNetwork.scala 156:83]
      r_lvl_output_ff_7 <= w_vn_lvl_0_7; // @[FanNetwork.scala 157:24]
    end else begin
      r_lvl_output_ff_7 <= 32'h0;
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_8 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_0_valid_9 & w_vn_lvl_0_valid_8) begin // @[FanNetwork.scala 174:61]
      r_lvl_output_ff_8 <= w_vn_lvl_0_8; // @[FanNetwork.scala 176:24]
    end else if (w_vn_lvl_0_valid_9 & ~w_vn_lvl_0_valid_8) begin // @[FanNetwork.scala 179:68]
      r_lvl_output_ff_8 <= 32'h0; // @[FanNetwork.scala 181:24]
    end else if (~w_vn_lvl_0_valid_9 & w_vn_lvl_0_valid_8) begin // @[FanNetwork.scala 184:68]
      r_lvl_output_ff_8 <= w_vn_lvl_0_8; // @[FanNetwork.scala 186:24]
    end else begin
      r_lvl_output_ff_8 <= 32'h0; // @[FanNetwork.scala 191:24]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_9 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_0_valid_9 & w_vn_lvl_0_valid_8) begin // @[FanNetwork.scala 174:61]
      r_lvl_output_ff_9 <= w_vn_lvl_0_9; // @[FanNetwork.scala 175:24]
    end else if (w_vn_lvl_0_valid_9 & ~w_vn_lvl_0_valid_8) begin // @[FanNetwork.scala 179:68]
      r_lvl_output_ff_9 <= w_vn_lvl_0_9; // @[FanNetwork.scala 180:24]
    end else begin
      r_lvl_output_ff_9 <= 32'h0;
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_10 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_0_valid_11 & w_vn_lvl_0_valid_10) begin // @[FanNetwork.scala 197:63]
      r_lvl_output_ff_10 <= w_vn_lvl_0_10; // @[FanNetwork.scala 199:25]
    end else if (w_vn_lvl_0_valid_11 & ~w_vn_lvl_0_valid_10) begin // @[FanNetwork.scala 202:70]
      r_lvl_output_ff_10 <= 32'h0; // @[FanNetwork.scala 204:25]
    end else if (~w_vn_lvl_0_valid_11 & w_vn_lvl_0_valid_10) begin // @[FanNetwork.scala 207:70]
      r_lvl_output_ff_10 <= w_vn_lvl_0_10; // @[FanNetwork.scala 209:25]
    end else begin
      r_lvl_output_ff_10 <= 32'h0; // @[FanNetwork.scala 214:25]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_11 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_11 <= r_lvl_output_ff_79; // @[FanNetwork.scala 829:25]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_12 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_0_valid_13 & w_vn_lvl_0_valid_12) begin // @[FanNetwork.scala 220:63]
      r_lvl_output_ff_12 <= w_vn_lvl_0_12; // @[FanNetwork.scala 222:25]
    end else if (w_vn_lvl_0_valid_13 & ~w_vn_lvl_0_valid_12) begin // @[FanNetwork.scala 225:70]
      r_lvl_output_ff_12 <= 32'h0; // @[FanNetwork.scala 227:25]
    end else if (~w_vn_lvl_0_valid_13 & w_vn_lvl_0_valid_12) begin // @[FanNetwork.scala 230:70]
      r_lvl_output_ff_12 <= w_vn_lvl_0_12; // @[FanNetwork.scala 232:25]
    end else begin
      r_lvl_output_ff_12 <= 32'h0; // @[FanNetwork.scala 237:25]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_13 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_0_valid_13 & w_vn_lvl_0_valid_12) begin // @[FanNetwork.scala 220:63]
      r_lvl_output_ff_13 <= w_vn_lvl_0_13; // @[FanNetwork.scala 221:25]
    end else if (w_vn_lvl_0_valid_13 & ~w_vn_lvl_0_valid_12) begin // @[FanNetwork.scala 225:70]
      r_lvl_output_ff_13 <= w_vn_lvl_0_13; // @[FanNetwork.scala 226:25]
    end else begin
      r_lvl_output_ff_13 <= 32'h0;
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_14 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_0_valid_15 & w_vn_lvl_0_valid_14) begin // @[FanNetwork.scala 243:63]
      r_lvl_output_ff_14 <= w_vn_lvl_0_14; // @[FanNetwork.scala 245:25]
    end else if (w_vn_lvl_0_valid_15 & ~w_vn_lvl_0_valid_14) begin // @[FanNetwork.scala 248:70]
      r_lvl_output_ff_14 <= 32'h0; // @[FanNetwork.scala 250:25]
    end else if (~w_vn_lvl_0_valid_15 & w_vn_lvl_0_valid_14) begin // @[FanNetwork.scala 253:70]
      r_lvl_output_ff_14 <= w_vn_lvl_0_14; // @[FanNetwork.scala 255:25]
    end else begin
      r_lvl_output_ff_14 <= 32'h0; // @[FanNetwork.scala 260:25]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_15 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_0_valid_15 & w_vn_lvl_0_valid_14) begin // @[FanNetwork.scala 243:63]
      r_lvl_output_ff_15 <= w_vn_lvl_0_15; // @[FanNetwork.scala 244:25]
    end else if (w_vn_lvl_0_valid_15 & ~w_vn_lvl_0_valid_14) begin // @[FanNetwork.scala 248:70]
      r_lvl_output_ff_15 <= w_vn_lvl_0_15; // @[FanNetwork.scala 249:25]
    end else begin
      r_lvl_output_ff_15 <= 32'h0;
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_16 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_0_valid_17 & w_vn_lvl_0_valid_16) begin // @[FanNetwork.scala 266:63]
      r_lvl_output_ff_16 <= w_vn_lvl_0_16; // @[FanNetwork.scala 268:25]
    end else if (w_vn_lvl_0_valid_17 & ~w_vn_lvl_0_valid_16) begin // @[FanNetwork.scala 271:70]
      r_lvl_output_ff_16 <= 32'h0; // @[FanNetwork.scala 273:25]
    end else if (~w_vn_lvl_0_valid_17 & w_vn_lvl_0_valid_16) begin // @[FanNetwork.scala 276:70]
      r_lvl_output_ff_16 <= w_vn_lvl_0_16; // @[FanNetwork.scala 278:25]
    end else begin
      r_lvl_output_ff_16 <= 32'h0; // @[FanNetwork.scala 283:25]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_17 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_0_valid_17 & w_vn_lvl_0_valid_16) begin // @[FanNetwork.scala 266:63]
      r_lvl_output_ff_17 <= w_vn_lvl_0_17; // @[FanNetwork.scala 267:25]
    end else if (w_vn_lvl_0_valid_17 & ~w_vn_lvl_0_valid_16) begin // @[FanNetwork.scala 271:70]
      r_lvl_output_ff_17 <= w_vn_lvl_0_17; // @[FanNetwork.scala 272:25]
    end else begin
      r_lvl_output_ff_17 <= 32'h0;
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_18 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_0_valid_19 & w_vn_lvl_0_valid_18) begin // @[FanNetwork.scala 289:63]
      r_lvl_output_ff_18 <= w_vn_lvl_0_18; // @[FanNetwork.scala 291:25]
    end else if (w_vn_lvl_0_valid_19 & ~w_vn_lvl_0_valid_18) begin // @[FanNetwork.scala 294:70]
      r_lvl_output_ff_18 <= 32'h0; // @[FanNetwork.scala 296:25]
    end else if (~w_vn_lvl_0_valid_19 & w_vn_lvl_0_valid_18) begin // @[FanNetwork.scala 299:70]
      r_lvl_output_ff_18 <= w_vn_lvl_0_18; // @[FanNetwork.scala 301:25]
    end else begin
      r_lvl_output_ff_18 <= 32'h0; // @[FanNetwork.scala 306:25]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_19 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_0_valid_19 & w_vn_lvl_0_valid_18) begin // @[FanNetwork.scala 289:63]
      r_lvl_output_ff_19 <= w_vn_lvl_0_19; // @[FanNetwork.scala 290:25]
    end else if (w_vn_lvl_0_valid_19 & ~w_vn_lvl_0_valid_18) begin // @[FanNetwork.scala 294:70]
      r_lvl_output_ff_19 <= w_vn_lvl_0_19; // @[FanNetwork.scala 295:25]
    end else begin
      r_lvl_output_ff_19 <= 32'h0;
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_20 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_0_valid_21 & w_vn_lvl_0_valid_20) begin // @[FanNetwork.scala 312:63]
      r_lvl_output_ff_20 <= w_vn_lvl_0_20; // @[FanNetwork.scala 314:25]
    end else if (w_vn_lvl_0_valid_21 & ~w_vn_lvl_0_valid_20) begin // @[FanNetwork.scala 317:70]
      r_lvl_output_ff_20 <= 32'h0; // @[FanNetwork.scala 319:25]
    end else if (~w_vn_lvl_0_valid_21 & w_vn_lvl_0_valid_20) begin // @[FanNetwork.scala 322:70]
      r_lvl_output_ff_20 <= w_vn_lvl_0_20; // @[FanNetwork.scala 324:25]
    end else begin
      r_lvl_output_ff_20 <= 32'h0; // @[FanNetwork.scala 329:25]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_21 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_0_valid_21 & w_vn_lvl_0_valid_20) begin // @[FanNetwork.scala 312:63]
      r_lvl_output_ff_21 <= w_vn_lvl_0_21; // @[FanNetwork.scala 313:25]
    end else if (w_vn_lvl_0_valid_21 & ~w_vn_lvl_0_valid_20) begin // @[FanNetwork.scala 317:70]
      r_lvl_output_ff_21 <= w_vn_lvl_0_21; // @[FanNetwork.scala 318:25]
    end else begin
      r_lvl_output_ff_21 <= 32'h0;
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_22 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_0_valid_23 & w_vn_lvl_0_valid_22) begin // @[FanNetwork.scala 335:63]
      r_lvl_output_ff_22 <= w_vn_lvl_0_22; // @[FanNetwork.scala 337:25]
    end else if (w_vn_lvl_0_valid_23 & ~w_vn_lvl_0_valid_22) begin // @[FanNetwork.scala 340:70]
      r_lvl_output_ff_22 <= 32'h0; // @[FanNetwork.scala 342:25]
    end else if (~w_vn_lvl_0_valid_23 & w_vn_lvl_0_valid_22) begin // @[FanNetwork.scala 345:70]
      r_lvl_output_ff_22 <= w_vn_lvl_0_22; // @[FanNetwork.scala 347:25]
    end else begin
      r_lvl_output_ff_22 <= 32'h0; // @[FanNetwork.scala 352:25]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_23 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_0_valid_23 & w_vn_lvl_0_valid_22) begin // @[FanNetwork.scala 335:63]
      r_lvl_output_ff_23 <= w_vn_lvl_0_23; // @[FanNetwork.scala 336:25]
    end else if (w_vn_lvl_0_valid_23 & ~w_vn_lvl_0_valid_22) begin // @[FanNetwork.scala 340:70]
      r_lvl_output_ff_23 <= w_vn_lvl_0_23; // @[FanNetwork.scala 341:25]
    end else begin
      r_lvl_output_ff_23 <= 32'h0;
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_24 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_0_valid_25 & w_vn_lvl_0_valid_24) begin // @[FanNetwork.scala 358:63]
      r_lvl_output_ff_24 <= w_vn_lvl_0_24; // @[FanNetwork.scala 360:25]
    end else if (w_vn_lvl_0_valid_25 & ~w_vn_lvl_0_valid_24) begin // @[FanNetwork.scala 363:70]
      r_lvl_output_ff_24 <= 32'h0; // @[FanNetwork.scala 365:25]
    end else if (~w_vn_lvl_0_valid_25 & w_vn_lvl_0_valid_24) begin // @[FanNetwork.scala 368:70]
      r_lvl_output_ff_24 <= w_vn_lvl_0_24; // @[FanNetwork.scala 370:25]
    end else begin
      r_lvl_output_ff_24 <= 32'h0; // @[FanNetwork.scala 375:25]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_25 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_0_valid_25 & w_vn_lvl_0_valid_24) begin // @[FanNetwork.scala 358:63]
      r_lvl_output_ff_25 <= w_vn_lvl_0_25; // @[FanNetwork.scala 359:25]
    end else if (w_vn_lvl_0_valid_25 & ~w_vn_lvl_0_valid_24) begin // @[FanNetwork.scala 363:70]
      r_lvl_output_ff_25 <= w_vn_lvl_0_25; // @[FanNetwork.scala 364:25]
    end else begin
      r_lvl_output_ff_25 <= 32'h0;
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_26 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_0_valid_27 & w_vn_lvl_0_valid_26) begin // @[FanNetwork.scala 381:63]
      r_lvl_output_ff_26 <= w_vn_lvl_0_26; // @[FanNetwork.scala 383:25]
    end else if (w_vn_lvl_0_valid_27 & ~w_vn_lvl_0_valid_26) begin // @[FanNetwork.scala 386:70]
      r_lvl_output_ff_26 <= 32'h0; // @[FanNetwork.scala 388:25]
    end else if (~w_vn_lvl_0_valid_27 & w_vn_lvl_0_valid_26) begin // @[FanNetwork.scala 391:70]
      r_lvl_output_ff_26 <= w_vn_lvl_0_26; // @[FanNetwork.scala 393:25]
    end else begin
      r_lvl_output_ff_26 <= 32'h0; // @[FanNetwork.scala 398:25]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_27 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_0_valid_27 & w_vn_lvl_0_valid_26) begin // @[FanNetwork.scala 381:63]
      r_lvl_output_ff_27 <= w_vn_lvl_0_27; // @[FanNetwork.scala 382:25]
    end else if (w_vn_lvl_0_valid_27 & ~w_vn_lvl_0_valid_26) begin // @[FanNetwork.scala 386:70]
      r_lvl_output_ff_27 <= w_vn_lvl_0_27; // @[FanNetwork.scala 387:25]
    end else begin
      r_lvl_output_ff_27 <= 32'h0;
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_28 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_0_valid_29 & w_vn_lvl_0_valid_28) begin // @[FanNetwork.scala 404:63]
      r_lvl_output_ff_28 <= w_vn_lvl_0_28; // @[FanNetwork.scala 406:25]
    end else if (w_vn_lvl_0_valid_29 & ~w_vn_lvl_0_valid_28) begin // @[FanNetwork.scala 409:70]
      r_lvl_output_ff_28 <= 32'h0; // @[FanNetwork.scala 411:25]
    end else if (~w_vn_lvl_0_valid_29 & w_vn_lvl_0_valid_28) begin // @[FanNetwork.scala 414:70]
      r_lvl_output_ff_28 <= w_vn_lvl_0_28; // @[FanNetwork.scala 416:25]
    end else begin
      r_lvl_output_ff_28 <= 32'h0; // @[FanNetwork.scala 421:25]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_29 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_0_valid_29 & w_vn_lvl_0_valid_28) begin // @[FanNetwork.scala 404:63]
      r_lvl_output_ff_29 <= w_vn_lvl_0_29; // @[FanNetwork.scala 405:25]
    end else if (w_vn_lvl_0_valid_29 & ~w_vn_lvl_0_valid_28) begin // @[FanNetwork.scala 409:70]
      r_lvl_output_ff_29 <= w_vn_lvl_0_29; // @[FanNetwork.scala 410:25]
    end else begin
      r_lvl_output_ff_29 <= 32'h0;
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_30 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_0_valid_31 & w_vn_lvl_0_valid_30) begin // @[FanNetwork.scala 427:62]
      r_lvl_output_ff_30 <= w_vn_lvl_0_30; // @[FanNetwork.scala 429:25]
    end else if (w_vn_lvl_0_valid_31 & ~w_vn_lvl_0_valid_30) begin // @[FanNetwork.scala 432:69]
      r_lvl_output_ff_30 <= 32'h0; // @[FanNetwork.scala 434:25]
    end else if (~w_vn_lvl_0_valid_31 & w_vn_lvl_0_valid_30) begin // @[FanNetwork.scala 437:69]
      r_lvl_output_ff_30 <= w_vn_lvl_0_30; // @[FanNetwork.scala 439:25]
    end else begin
      r_lvl_output_ff_30 <= 32'h0; // @[FanNetwork.scala 444:25]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_31 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_0_valid_31 & w_vn_lvl_0_valid_30) begin // @[FanNetwork.scala 427:62]
      r_lvl_output_ff_31 <= w_vn_lvl_0_31; // @[FanNetwork.scala 428:25]
    end else if (w_vn_lvl_0_valid_31 & ~w_vn_lvl_0_valid_30) begin // @[FanNetwork.scala 432:69]
      r_lvl_output_ff_31 <= w_vn_lvl_0_31; // @[FanNetwork.scala 433:25]
    end else begin
      r_lvl_output_ff_31 <= 32'h0;
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_32 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_32 <= r_lvl_output_ff_0; // @[FanNetwork.scala 452:25]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_33 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_1_valid_0) begin // @[FanNetwork.scala 455:34]
      r_lvl_output_ff_33 <= w_vn_lvl_1_0; // @[FanNetwork.scala 456:29]
    end else begin
      r_lvl_output_ff_33 <= r_lvl_output_ff_1; // @[FanNetwork.scala 459:29]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_34 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_1_valid_1) begin // @[FanNetwork.scala 463:34]
      r_lvl_output_ff_34 <= w_vn_lvl_1_1; // @[FanNetwork.scala 464:29]
    end else begin
      r_lvl_output_ff_34 <= r_lvl_output_ff_2; // @[FanNetwork.scala 467:29]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_35 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_35 <= r_lvl_output_ff_3; // @[FanNetwork.scala 471:25]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_37 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_1_valid_2) begin // @[FanNetwork.scala 477:34]
      r_lvl_output_ff_37 <= w_vn_lvl_1_2; // @[FanNetwork.scala 478:29]
    end else begin
      r_lvl_output_ff_37 <= 32'h0; // @[FanNetwork.scala 481:29]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_38 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_1_valid_3) begin // @[FanNetwork.scala 485:34]
      r_lvl_output_ff_38 <= w_vn_lvl_1_3; // @[FanNetwork.scala 486:29]
    end else begin
      r_lvl_output_ff_38 <= r_lvl_output_ff_6; // @[FanNetwork.scala 489:29]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_39 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_39 <= r_lvl_output_ff_7; // @[FanNetwork.scala 495:25]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_40 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_40 <= r_lvl_output_ff_8; // @[FanNetwork.scala 498:25]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_41 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_1_valid_4) begin // @[FanNetwork.scala 501:34]
      r_lvl_output_ff_41 <= w_vn_lvl_1_4; // @[FanNetwork.scala 502:29]
    end else begin
      r_lvl_output_ff_41 <= r_lvl_output_ff_9; // @[FanNetwork.scala 505:29]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_42 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_1_valid_5) begin // @[FanNetwork.scala 508:34]
      r_lvl_output_ff_42 <= w_vn_lvl_1_5; // @[FanNetwork.scala 509:29]
    end else begin
      r_lvl_output_ff_42 <= r_lvl_output_ff_10; // @[FanNetwork.scala 512:29]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_43 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_43 <= r_lvl_output_ff_11; // @[FanNetwork.scala 516:25]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_44 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_44 <= r_lvl_output_ff_12; // @[FanNetwork.scala 519:25]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_45 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_1_valid_6) begin // @[FanNetwork.scala 522:34]
      r_lvl_output_ff_45 <= w_vn_lvl_1_6; // @[FanNetwork.scala 523:29]
    end else begin
      r_lvl_output_ff_45 <= r_lvl_output_ff_13; // @[FanNetwork.scala 526:29]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_46 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_1_valid_7) begin // @[FanNetwork.scala 530:34]
      r_lvl_output_ff_46 <= w_vn_lvl_1_7; // @[FanNetwork.scala 531:29]
    end else begin
      r_lvl_output_ff_46 <= r_lvl_output_ff_14; // @[FanNetwork.scala 534:29]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_47 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_47 <= r_lvl_output_ff_15; // @[FanNetwork.scala 537:25]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_48 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_48 <= r_lvl_output_ff_16; // @[FanNetwork.scala 540:25]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_49 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_1_valid_8) begin // @[FanNetwork.scala 543:34]
      r_lvl_output_ff_49 <= w_vn_lvl_1_8; // @[FanNetwork.scala 544:29]
    end else begin
      r_lvl_output_ff_49 <= r_lvl_output_ff_17; // @[FanNetwork.scala 547:29]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_50 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_1_valid_9) begin // @[FanNetwork.scala 551:34]
      r_lvl_output_ff_50 <= w_vn_lvl_1_9; // @[FanNetwork.scala 552:29]
    end else begin
      r_lvl_output_ff_50 <= r_lvl_output_ff_18; // @[FanNetwork.scala 555:29]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_51 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_51 <= r_lvl_output_ff_19; // @[FanNetwork.scala 561:25]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_52 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_52 <= r_lvl_output_ff_20; // @[FanNetwork.scala 564:25]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_53 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_1_valid_10) begin // @[FanNetwork.scala 567:35]
      r_lvl_output_ff_53 <= w_vn_lvl_1_10; // @[FanNetwork.scala 568:29]
    end else begin
      r_lvl_output_ff_53 <= r_lvl_output_ff_21; // @[FanNetwork.scala 571:29]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_54 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_1_valid_11) begin // @[FanNetwork.scala 575:35]
      r_lvl_output_ff_54 <= w_vn_lvl_1_11; // @[FanNetwork.scala 576:29]
    end else begin
      r_lvl_output_ff_54 <= r_lvl_output_ff_22; // @[FanNetwork.scala 579:29]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_55 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_55 <= r_lvl_output_ff_23; // @[FanNetwork.scala 583:25]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_56 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_56 <= r_lvl_output_ff_24; // @[FanNetwork.scala 586:25]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_57 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_1_valid_12) begin // @[FanNetwork.scala 589:35]
      r_lvl_output_ff_57 <= w_vn_lvl_1_12; // @[FanNetwork.scala 590:29]
    end else begin
      r_lvl_output_ff_57 <= r_lvl_output_ff_25; // @[FanNetwork.scala 593:29]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_58 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_1_valid_13) begin // @[FanNetwork.scala 597:35]
      r_lvl_output_ff_58 <= w_vn_lvl_1_13; // @[FanNetwork.scala 598:29]
    end else begin
      r_lvl_output_ff_58 <= r_lvl_output_ff_26; // @[FanNetwork.scala 601:29]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_59 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_59 <= r_lvl_output_ff_27; // @[FanNetwork.scala 605:25]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_60 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_60 <= r_lvl_output_ff_28; // @[FanNetwork.scala 608:25]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_61 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_1_valid_14) begin // @[FanNetwork.scala 611:43]
      r_lvl_output_ff_61 <= w_vn_lvl_1_14; // @[FanNetwork.scala 612:29]
    end else begin
      r_lvl_output_ff_61 <= r_lvl_output_ff_29; // @[FanNetwork.scala 615:29]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_62 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_1_valid_15) begin // @[FanNetwork.scala 619:43]
      r_lvl_output_ff_62 <= w_vn_lvl_1_15; // @[FanNetwork.scala 620:29]
    end else begin
      r_lvl_output_ff_62 <= r_lvl_output_ff_30; // @[FanNetwork.scala 623:29]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_63 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_63 <= r_lvl_output_ff_31; // @[FanNetwork.scala 627:25]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_64 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_64 <= r_lvl_output_ff_32; // @[FanNetwork.scala 636:26]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_65 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_65 <= r_lvl_output_ff_33; // @[FanNetwork.scala 639:25]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_66 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_66 <= r_lvl_output_ff_34; // @[FanNetwork.scala 642:25]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_67 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_2_valid_0) begin // @[FanNetwork.scala 645:43]
      r_lvl_output_ff_67 <= w_vn_lvl_2_0; // @[FanNetwork.scala 646:29]
    end else begin
      r_lvl_output_ff_67 <= r_lvl_output_ff_35; // @[FanNetwork.scala 649:33]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_68 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_2_valid_1) begin // @[FanNetwork.scala 653:43]
      r_lvl_output_ff_68 <= w_vn_lvl_2_1; // @[FanNetwork.scala 654:29]
    end else begin
      r_lvl_output_ff_68 <= 32'h0; // @[FanNetwork.scala 657:29]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_69 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_69 <= r_lvl_output_ff_37; // @[FanNetwork.scala 661:25]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_70 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_70 <= r_lvl_output_ff_38; // @[FanNetwork.scala 664:25]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_71 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_71 <= r_lvl_output_ff_39; // @[FanNetwork.scala 667:25]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_72 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_72 <= r_lvl_output_ff_40; // @[FanNetwork.scala 670:25]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_73 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_73 <= r_lvl_output_ff_41; // @[FanNetwork.scala 673:25]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_74 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_74 <= r_lvl_output_ff_42; // @[FanNetwork.scala 676:25]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_75 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_2_valid_2) begin // @[FanNetwork.scala 679:43]
      r_lvl_output_ff_75 <= w_vn_lvl_2_2; // @[FanNetwork.scala 680:29]
    end else begin
      r_lvl_output_ff_75 <= r_lvl_output_ff_43; // @[FanNetwork.scala 683:29]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_76 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_2_valid_3) begin // @[FanNetwork.scala 687:43]
      r_lvl_output_ff_76 <= w_vn_lvl_2_3; // @[FanNetwork.scala 688:29]
    end else begin
      r_lvl_output_ff_76 <= r_lvl_output_ff_44; // @[FanNetwork.scala 691:29]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_77 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_77 <= r_lvl_output_ff_45; // @[FanNetwork.scala 695:25]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_78 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_78 <= r_lvl_output_ff_46; // @[FanNetwork.scala 698:25]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_79 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_79 <= r_lvl_output_ff_47; // @[FanNetwork.scala 701:25]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_80 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_80 <= r_lvl_output_ff_48; // @[FanNetwork.scala 704:25]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_81 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_81 <= r_lvl_output_ff_49; // @[FanNetwork.scala 707:25]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_82 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_82 <= r_lvl_output_ff_50; // @[FanNetwork.scala 710:25]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_83 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_2_valid_4) begin // @[FanNetwork.scala 713:43]
      r_lvl_output_ff_83 <= w_vn_lvl_2_4; // @[FanNetwork.scala 714:29]
    end else begin
      r_lvl_output_ff_83 <= r_lvl_output_ff_51; // @[FanNetwork.scala 717:29]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_84 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_2_valid_5) begin // @[FanNetwork.scala 721:40]
      r_lvl_output_ff_84 <= w_vn_lvl_2_5; // @[FanNetwork.scala 722:29]
    end else begin
      r_lvl_output_ff_84 <= r_lvl_output_ff_52; // @[FanNetwork.scala 725:29]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_85 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_85 <= r_lvl_output_ff_53; // @[FanNetwork.scala 729:25]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_86 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_86 <= r_lvl_output_ff_54; // @[FanNetwork.scala 732:25]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_87 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_87 <= r_lvl_output_ff_55; // @[FanNetwork.scala 735:25]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_88 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_88 <= r_lvl_output_ff_56; // @[FanNetwork.scala 738:25]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_89 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_89 <= r_lvl_output_ff_57; // @[FanNetwork.scala 741:25]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_90 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_90 <= r_lvl_output_ff_58; // @[FanNetwork.scala 744:25]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_91 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_2_valid_6) begin // @[FanNetwork.scala 747:40]
      r_lvl_output_ff_91 <= w_vn_lvl_2_6; // @[FanNetwork.scala 748:29]
    end else begin
      r_lvl_output_ff_91 <= r_lvl_output_ff_59; // @[FanNetwork.scala 751:29]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_92 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_2_valid_7) begin // @[FanNetwork.scala 755:40]
      r_lvl_output_ff_92 <= w_vn_lvl_2_7; // @[FanNetwork.scala 756:29]
    end else begin
      r_lvl_output_ff_92 <= r_lvl_output_ff_60; // @[FanNetwork.scala 759:29]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_93 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_93 <= r_lvl_output_ff_61; // @[FanNetwork.scala 763:25]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_94 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_94 <= r_lvl_output_ff_62; // @[FanNetwork.scala 766:25]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_95 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_95 <= r_lvl_output_ff_63; // @[FanNetwork.scala 769:25]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_96 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_96 <= r_lvl_output_ff_64; // @[FanNetwork.scala 774:25]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_97 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_97 <= r_lvl_output_ff_65; // @[FanNetwork.scala 777:25]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_98 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_98 <= r_lvl_output_ff_66; // @[FanNetwork.scala 780:25]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_99 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_99 <= r_lvl_output_ff_67; // @[FanNetwork.scala 783:25]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_100 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_100 <= r_lvl_output_ff_68; // @[FanNetwork.scala 786:26]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_101 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_101 <= r_lvl_output_ff_69; // @[FanNetwork.scala 789:26]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_102 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_102 <= r_lvl_output_ff_70; // @[FanNetwork.scala 792:26]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_103 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_3_valid_0) begin // @[FanNetwork.scala 795:40]
      r_lvl_output_ff_103 <= w_vn_lvl_3_0; // @[FanNetwork.scala 796:28]
    end else begin
      r_lvl_output_ff_103 <= r_lvl_output_ff_71; // @[FanNetwork.scala 799:28]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_104 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_3_valid_1) begin // @[FanNetwork.scala 803:40]
      r_lvl_output_ff_104 <= w_vn_lvl_3_1; // @[FanNetwork.scala 804:28]
    end else begin
      r_lvl_output_ff_104 <= r_lvl_output_ff_72; // @[FanNetwork.scala 807:28]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_105 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_105 <= r_lvl_output_ff_73; // @[FanNetwork.scala 811:26]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_106 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_106 <= r_lvl_output_ff_74; // @[FanNetwork.scala 814:26]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_107 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_107 <= r_lvl_output_ff_75; // @[FanNetwork.scala 817:26]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_108 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_108 <= r_lvl_output_ff_76; // @[FanNetwork.scala 820:26]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_109 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_109 <= r_lvl_output_ff_77; // @[FanNetwork.scala 823:26]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_110 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_110 <= r_lvl_output_ff_78; // @[FanNetwork.scala 826:26]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_112 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_112 <= r_lvl_output_ff_80; // @[FanNetwork.scala 832:26]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_113 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_113 <= r_lvl_output_ff_81; // @[FanNetwork.scala 835:26]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_114 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_114 <= r_lvl_output_ff_82; // @[FanNetwork.scala 838:26]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_115 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_115 <= r_lvl_output_ff_83; // @[FanNetwork.scala 841:26]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_116 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_116 <= r_lvl_output_ff_84; // @[FanNetwork.scala 844:26]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_117 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_117 <= r_lvl_output_ff_85; // @[FanNetwork.scala 847:26]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_118 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_118 <= r_lvl_output_ff_86; // @[FanNetwork.scala 850:26]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_119 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_3_valid_2) begin // @[FanNetwork.scala 853:40]
      r_lvl_output_ff_119 <= w_vn_lvl_3_2; // @[FanNetwork.scala 854:30]
    end else begin
      r_lvl_output_ff_119 <= r_lvl_output_ff_87; // @[FanNetwork.scala 857:30]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_120 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_3_valid_3) begin // @[FanNetwork.scala 861:41]
      r_lvl_output_ff_120 <= w_vn_lvl_3_3; // @[FanNetwork.scala 862:30]
    end else begin
      r_lvl_output_ff_120 <= r_lvl_output_ff_88; // @[FanNetwork.scala 865:30]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_121 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_121 <= r_lvl_output_ff_89; // @[FanNetwork.scala 869:26]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_122 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_122 <= r_lvl_output_ff_90; // @[FanNetwork.scala 872:26]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_123 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_123 <= r_lvl_output_ff_91; // @[FanNetwork.scala 875:26]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_124 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_124 <= r_lvl_output_ff_92; // @[FanNetwork.scala 878:26]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_125 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_125 <= r_lvl_output_ff_93; // @[FanNetwork.scala 881:26]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_126 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_126 <= r_lvl_output_ff_94; // @[FanNetwork.scala 884:26]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_127 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_127 <= r_lvl_output_ff_95; // @[FanNetwork.scala 887:26]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_128 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_128 <= r_lvl_output_ff_96; // @[FanNetwork.scala 899:26]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_129 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_129 <= r_lvl_output_ff_97; // @[FanNetwork.scala 902:26]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_130 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_130 <= r_lvl_output_ff_98; // @[FanNetwork.scala 905:26]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_131 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_131 <= r_lvl_output_ff_99; // @[FanNetwork.scala 908:26]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_132 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_132 <= r_lvl_output_ff_100; // @[FanNetwork.scala 911:26]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_133 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_133 <= r_lvl_output_ff_101; // @[FanNetwork.scala 914:26]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_134 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_134 <= r_lvl_output_ff_102; // @[FanNetwork.scala 917:26]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_135 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_135 <= r_lvl_output_ff_103; // @[FanNetwork.scala 920:26]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_136 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_136 <= r_lvl_output_ff_104; // @[FanNetwork.scala 923:26]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_137 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_137 <= r_lvl_output_ff_105; // @[FanNetwork.scala 926:26]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_138 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_138 <= r_lvl_output_ff_106; // @[FanNetwork.scala 929:26]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_139 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_139 <= r_lvl_output_ff_107; // @[FanNetwork.scala 932:26]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_140 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_140 <= r_lvl_output_ff_108; // @[FanNetwork.scala 935:26]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_141 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_141 <= r_lvl_output_ff_109; // @[FanNetwork.scala 938:26]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_142 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_142 <= r_lvl_output_ff_110; // @[FanNetwork.scala 941:26]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_143 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_4_valid_0) begin // @[FanNetwork.scala 944:40]
      r_lvl_output_ff_143 <= w_vn_lvl_4_0; // @[FanNetwork.scala 945:30]
    end else begin
      r_lvl_output_ff_143 <= 32'h0; // @[FanNetwork.scala 948:30]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_144 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else if (w_vn_lvl_4_valid_1) begin // @[FanNetwork.scala 952:40]
      r_lvl_output_ff_144 <= w_vn_lvl_4_1; // @[FanNetwork.scala 953:30]
    end else begin
      r_lvl_output_ff_144 <= r_lvl_output_ff_112; // @[FanNetwork.scala 956:30]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_145 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_145 <= r_lvl_output_ff_113; // @[FanNetwork.scala 960:26]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_146 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_146 <= r_lvl_output_ff_114; // @[FanNetwork.scala 963:26]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_147 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_147 <= r_lvl_output_ff_115; // @[FanNetwork.scala 966:26]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_148 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_148 <= r_lvl_output_ff_116; // @[FanNetwork.scala 969:26]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_149 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_149 <= r_lvl_output_ff_117; // @[FanNetwork.scala 972:26]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_150 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_150 <= r_lvl_output_ff_118; // @[FanNetwork.scala 975:26]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_151 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_151 <= r_lvl_output_ff_119; // @[FanNetwork.scala 978:26]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_152 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_152 <= r_lvl_output_ff_120; // @[FanNetwork.scala 981:26]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_153 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_153 <= r_lvl_output_ff_121; // @[FanNetwork.scala 984:26]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_154 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_154 <= r_lvl_output_ff_122; // @[FanNetwork.scala 987:26]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_155 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_155 <= r_lvl_output_ff_123; // @[FanNetwork.scala 990:26]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_156 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_156 <= r_lvl_output_ff_124; // @[FanNetwork.scala 993:26]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_157 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_157 <= r_lvl_output_ff_125; // @[FanNetwork.scala 996:26]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_158 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_158 <= r_lvl_output_ff_126; // @[FanNetwork.scala 999:26]
    end
    if (reset) begin // @[FanNetwork.scala 50:34]
      r_lvl_output_ff_159 <= 32'h0; // @[FanNetwork.scala 50:34]
    end else begin
      r_lvl_output_ff_159 <= r_lvl_output_ff_127; // @[FanNetwork.scala 1002:26]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_0 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_0 <= _GEN_10;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_1 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_1 <= _GEN_9;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_2 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_2 <= _GEN_21;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_3 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_3 <= _GEN_20;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_4 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_4 <= _GEN_32;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_5 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_5 <= _GEN_31;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_6 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_6 <= _GEN_43;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_7 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_7 <= _GEN_42;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_8 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_8 <= _GEN_54;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_9 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_9 <= _GEN_53;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_10 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_10 <= _GEN_65;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_11 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_11 <= _GEN_64;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_12 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_12 <= _GEN_76;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_13 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_13 <= _GEN_75;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_14 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_14 <= _GEN_87;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_15 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_15 <= _GEN_86;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_16 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_16 <= _GEN_98;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_17 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_17 <= _GEN_97;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_18 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_18 <= _GEN_109;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_19 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_19 <= _GEN_108;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_20 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_20 <= _GEN_120;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_21 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_21 <= _GEN_119;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_22 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_22 <= _GEN_131;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_23 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_23 <= _GEN_130;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_24 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_24 <= _GEN_142;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_25 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_25 <= _GEN_141;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_26 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_26 <= _GEN_153;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_27 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_27 <= _GEN_152;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_28 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_28 <= _GEN_164;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_29 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_29 <= _GEN_163;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_30 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_30 <= _GEN_175;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_31 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_31 <= _GEN_174;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_32 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_32 <= r_lvl_output_ff_valid_0; // @[FanNetwork.scala 453:31]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_33 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_33 <= _GEN_177;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_34 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_34 <= _GEN_179;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_35 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_35 <= r_lvl_output_ff_valid_3; // @[FanNetwork.scala 472:31]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_36 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_36 <= r_lvl_output_ff_valid_4; // @[FanNetwork.scala 475:31]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_37 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_37 <= _GEN_181;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_38 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_38 <= _GEN_183;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_39 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_39 <= r_lvl_output_ff_valid_7; // @[FanNetwork.scala 496:31]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_40 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_40 <= r_lvl_output_ff_valid_8; // @[FanNetwork.scala 499:31]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_41 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_41 <= _GEN_185;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_42 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_42 <= _GEN_187;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_43 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_43 <= r_lvl_output_ff_valid_11; // @[FanNetwork.scala 517:31]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_44 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_44 <= r_lvl_output_ff_valid_12; // @[FanNetwork.scala 520:31]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_45 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_45 <= _GEN_189;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_46 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_46 <= _GEN_191;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_47 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_47 <= r_lvl_output_ff_valid_15; // @[FanNetwork.scala 538:31]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_48 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_48 <= r_lvl_output_ff_valid_16; // @[FanNetwork.scala 541:31]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_49 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_49 <= _GEN_193;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_50 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_50 <= _GEN_195;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_51 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_51 <= r_lvl_output_ff_valid_19; // @[FanNetwork.scala 562:31]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_52 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_52 <= r_lvl_output_ff_valid_20; // @[FanNetwork.scala 565:31]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_53 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_53 <= _GEN_197;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_54 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_54 <= _GEN_199;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_55 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_55 <= r_lvl_output_ff_valid_23; // @[FanNetwork.scala 584:31]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_56 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_56 <= r_lvl_output_ff_valid_24; // @[FanNetwork.scala 587:31]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_57 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_57 <= _GEN_201;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_58 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_58 <= _GEN_203;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_59 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_59 <= r_lvl_output_ff_valid_27; // @[FanNetwork.scala 606:31]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_60 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_60 <= r_lvl_output_ff_valid_28; // @[FanNetwork.scala 609:31]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_61 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_61 <= _GEN_205;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_62 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_62 <= _GEN_207;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_63 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_63 <= r_lvl_output_ff_valid_31; // @[FanNetwork.scala 628:31]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_64 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_64 <= r_lvl_output_ff_valid_32; // @[FanNetwork.scala 637:31]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_65 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_65 <= r_lvl_output_ff_valid_33; // @[FanNetwork.scala 640:31]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_66 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_66 <= r_lvl_output_ff_valid_34; // @[FanNetwork.scala 643:31]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_67 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_67 <= _GEN_209;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_68 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_68 <= _GEN_211;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_69 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_69 <= r_lvl_output_ff_valid_37; // @[FanNetwork.scala 662:31]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_70 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_70 <= r_lvl_output_ff_valid_38; // @[FanNetwork.scala 665:31]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_71 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_71 <= r_lvl_output_ff_valid_39; // @[FanNetwork.scala 668:31]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_72 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_72 <= r_lvl_output_ff_valid_40; // @[FanNetwork.scala 671:31]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_73 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_73 <= r_lvl_output_ff_valid_41; // @[FanNetwork.scala 674:31]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_74 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_74 <= r_lvl_output_ff_valid_42; // @[FanNetwork.scala 677:31]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_75 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_75 <= _GEN_213;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_76 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_76 <= _GEN_215;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_77 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_77 <= r_lvl_output_ff_valid_45; // @[FanNetwork.scala 696:31]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_78 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_78 <= r_lvl_output_ff_valid_46; // @[FanNetwork.scala 699:31]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_79 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_79 <= r_lvl_output_ff_valid_47; // @[FanNetwork.scala 702:31]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_80 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_80 <= r_lvl_output_ff_valid_48; // @[FanNetwork.scala 705:31]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_81 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_81 <= r_lvl_output_ff_valid_49; // @[FanNetwork.scala 708:31]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_82 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_82 <= r_lvl_output_ff_valid_50; // @[FanNetwork.scala 711:31]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_83 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_83 <= _GEN_217;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_84 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_84 <= _GEN_219;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_85 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_85 <= r_lvl_output_ff_valid_53; // @[FanNetwork.scala 730:31]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_86 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_86 <= r_lvl_output_ff_valid_54; // @[FanNetwork.scala 733:31]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_87 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_87 <= r_lvl_output_ff_valid_55; // @[FanNetwork.scala 736:31]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_88 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_88 <= r_lvl_output_ff_valid_56; // @[FanNetwork.scala 739:31]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_89 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_89 <= r_lvl_output_ff_valid_57; // @[FanNetwork.scala 742:31]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_90 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_90 <= r_lvl_output_ff_valid_58; // @[FanNetwork.scala 745:31]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_91 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_91 <= _GEN_221;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_92 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_92 <= _GEN_223;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_93 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_93 <= r_lvl_output_ff_valid_61; // @[FanNetwork.scala 764:31]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_94 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_94 <= r_lvl_output_ff_valid_62; // @[FanNetwork.scala 767:31]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_95 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_95 <= r_lvl_output_ff_valid_63; // @[FanNetwork.scala 770:31]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_96 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_96 <= r_lvl_output_ff_valid_64; // @[FanNetwork.scala 775:31]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_97 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_97 <= r_lvl_output_ff_valid_65; // @[FanNetwork.scala 778:31]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_98 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_98 <= r_lvl_output_ff_valid_66; // @[FanNetwork.scala 781:31]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_99 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_99 <= r_lvl_output_ff_valid_67; // @[FanNetwork.scala 784:31]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_100 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_100 <= r_lvl_output_ff_valid_68; // @[FanNetwork.scala 787:32]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_101 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_101 <= r_lvl_output_ff_valid_69; // @[FanNetwork.scala 790:32]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_102 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_102 <= r_lvl_output_ff_valid_70; // @[FanNetwork.scala 793:32]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_103 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_103 <= _GEN_225;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_104 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_104 <= _GEN_227;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_105 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_105 <= r_lvl_output_ff_valid_73; // @[FanNetwork.scala 812:32]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_106 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_106 <= r_lvl_output_ff_valid_74; // @[FanNetwork.scala 815:32]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_107 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_107 <= r_lvl_output_ff_valid_75; // @[FanNetwork.scala 818:32]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_108 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_108 <= r_lvl_output_ff_valid_76; // @[FanNetwork.scala 821:32]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_109 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_109 <= r_lvl_output_ff_valid_77; // @[FanNetwork.scala 824:32]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_110 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_110 <= r_lvl_output_ff_valid_78; // @[FanNetwork.scala 827:32]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_111 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_111 <= r_lvl_output_ff_valid_79; // @[FanNetwork.scala 830:32]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_112 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_112 <= r_lvl_output_ff_valid_80; // @[FanNetwork.scala 833:32]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_113 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_113 <= r_lvl_output_ff_valid_81; // @[FanNetwork.scala 836:32]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_114 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_114 <= r_lvl_output_ff_valid_82; // @[FanNetwork.scala 839:32]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_115 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_115 <= r_lvl_output_ff_valid_83; // @[FanNetwork.scala 842:32]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_116 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_116 <= r_lvl_output_ff_valid_84; // @[FanNetwork.scala 845:32]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_117 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_117 <= r_lvl_output_ff_valid_85; // @[FanNetwork.scala 848:32]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_118 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_118 <= r_lvl_output_ff_valid_86; // @[FanNetwork.scala 851:32]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_119 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_119 <= _GEN_229;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_120 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_120 <= _GEN_231;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_121 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_121 <= r_lvl_output_ff_valid_89; // @[FanNetwork.scala 870:32]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_122 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_122 <= r_lvl_output_ff_valid_90; // @[FanNetwork.scala 873:32]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_123 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_123 <= r_lvl_output_ff_valid_91; // @[FanNetwork.scala 876:32]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_124 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_124 <= r_lvl_output_ff_valid_92; // @[FanNetwork.scala 879:32]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_125 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_125 <= r_lvl_output_ff_valid_93; // @[FanNetwork.scala 882:32]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_126 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_126 <= r_lvl_output_ff_valid_94; // @[FanNetwork.scala 885:32]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_127 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_127 <= r_lvl_output_ff_valid_95; // @[FanNetwork.scala 888:32]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_128 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_128 <= r_lvl_output_ff_valid_96; // @[FanNetwork.scala 900:32]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_129 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_129 <= r_lvl_output_ff_valid_97; // @[FanNetwork.scala 903:32]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_130 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_130 <= r_lvl_output_ff_valid_98; // @[FanNetwork.scala 906:32]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_131 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_131 <= r_lvl_output_ff_valid_99; // @[FanNetwork.scala 909:32]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_132 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_132 <= r_lvl_output_ff_valid_100; // @[FanNetwork.scala 912:32]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_133 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_133 <= r_lvl_output_ff_valid_101; // @[FanNetwork.scala 915:32]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_134 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_134 <= r_lvl_output_ff_valid_102; // @[FanNetwork.scala 918:32]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_135 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_135 <= r_lvl_output_ff_valid_103; // @[FanNetwork.scala 921:32]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_136 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_136 <= r_lvl_output_ff_valid_104; // @[FanNetwork.scala 924:32]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_137 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_137 <= r_lvl_output_ff_valid_105; // @[FanNetwork.scala 927:32]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_138 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_138 <= r_lvl_output_ff_valid_106; // @[FanNetwork.scala 930:32]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_139 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_139 <= r_lvl_output_ff_valid_107; // @[FanNetwork.scala 933:32]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_140 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_140 <= r_lvl_output_ff_valid_108; // @[FanNetwork.scala 936:32]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_141 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_141 <= r_lvl_output_ff_valid_109; // @[FanNetwork.scala 939:32]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_142 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_142 <= r_lvl_output_ff_valid_110; // @[FanNetwork.scala 942:32]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_143 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_143 <= _GEN_233;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_144 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_144 <= _GEN_235;
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_145 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_145 <= r_lvl_output_ff_valid_113; // @[FanNetwork.scala 961:32]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_146 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_146 <= r_lvl_output_ff_valid_114; // @[FanNetwork.scala 964:32]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_147 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_147 <= r_lvl_output_ff_valid_115; // @[FanNetwork.scala 967:32]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_148 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_148 <= r_lvl_output_ff_valid_116; // @[FanNetwork.scala 970:32]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_149 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_149 <= r_lvl_output_ff_valid_117; // @[FanNetwork.scala 973:32]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_150 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_150 <= r_lvl_output_ff_valid_118; // @[FanNetwork.scala 976:32]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_151 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_151 <= r_lvl_output_ff_valid_119; // @[FanNetwork.scala 979:32]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_152 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_152 <= r_lvl_output_ff_valid_120; // @[FanNetwork.scala 982:32]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_153 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_153 <= r_lvl_output_ff_valid_121; // @[FanNetwork.scala 985:32]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_154 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_154 <= r_lvl_output_ff_valid_122; // @[FanNetwork.scala 988:32]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_155 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_155 <= r_lvl_output_ff_valid_123; // @[FanNetwork.scala 991:32]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_156 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_156 <= r_lvl_output_ff_valid_124; // @[FanNetwork.scala 994:32]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_157 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_157 <= r_lvl_output_ff_valid_125; // @[FanNetwork.scala 997:32]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_158 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_158 <= r_lvl_output_ff_valid_126; // @[FanNetwork.scala 1000:32]
    end
    if (reset) begin // @[FanNetwork.scala 51:40]
      r_lvl_output_ff_valid_159 <= 1'h0; // @[FanNetwork.scala 51:40]
    end else begin
      r_lvl_output_ff_valid_159 <= r_lvl_output_ff_valid_127; // @[FanNetwork.scala 1003:32]
    end
    if (reset) begin // @[FanNetwork.scala 52:26]
      r_valid_0 <= 1'h0; // @[FanNetwork.scala 52:26]
    end else begin
      r_valid_0 <= io_i_valid;
    end
    if (reset) begin // @[FanNetwork.scala 52:26]
      r_valid_1 <= 1'h0; // @[FanNetwork.scala 52:26]
    end else begin
      r_valid_1 <= r_valid_0; // @[FanNetwork.scala 1014:24]
    end
    if (reset) begin // @[FanNetwork.scala 52:26]
      r_valid_2 <= 1'h0; // @[FanNetwork.scala 52:26]
    end else begin
      r_valid_2 <= r_valid_1; // @[FanNetwork.scala 1014:24]
    end
    if (reset) begin // @[FanNetwork.scala 52:26]
      r_valid_3 <= 1'h0; // @[FanNetwork.scala 52:26]
    end else begin
      r_valid_3 <= r_valid_2; // @[FanNetwork.scala 1014:24]
    end
    if (reset) begin // @[FanNetwork.scala 52:26]
      r_valid_4 <= 1'h0; // @[FanNetwork.scala 52:26]
    end else begin
      r_valid_4 <= r_valid_3; // @[FanNetwork.scala 1014:24]
    end
    if (reset) begin // @[FanNetwork.scala 54:30]
      r_final_sum <= 32'h0; // @[FanNetwork.scala 54:30]
    end else begin
      r_final_sum <= w_fan_lvl_4_0; // @[FanNetwork.scala 1585:17]
    end
    if (reset) begin // @[FanNetwork.scala 55:30]
      r_final_add <= 1'h0; // @[FanNetwork.scala 55:30]
    end else begin
      r_final_add <= io_i_add_en_bus_30; // @[FanNetwork.scala 1583:17]
    end
    if (reset) begin // @[FanNetwork.scala 56:31]
      r_final_add2 <= 1'h0; // @[FanNetwork.scala 56:31]
    end else begin
      r_final_add2 <= r_final_add; // @[FanNetwork.scala 1584:18]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_fan_ff_lvl_0_to_4_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  r_fan_ff_lvl_0_to_4_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  r_fan_ff_lvl_0_to_3_0 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  r_fan_ff_lvl_0_to_3_1 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  r_fan_ff_lvl_0_to_3_2 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  r_fan_ff_lvl_0_to_3_3 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  r_fan_ff_lvl_0_to_3_4 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  r_fan_ff_lvl_0_to_3_5 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  r_fan_ff_lvl_0_to_2_0 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  r_fan_ff_lvl_0_to_2_1 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  r_fan_ff_lvl_0_to_2_2 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  r_fan_ff_lvl_0_to_2_3 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  r_fan_ff_lvl_0_to_2_4 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  r_fan_ff_lvl_0_to_2_5 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  r_fan_ff_lvl_0_to_2_6 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  r_fan_ff_lvl_0_to_2_7 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  r_fan_ff_lvl_0_to_2_8 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  r_fan_ff_lvl_0_to_2_9 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  r_fan_ff_lvl_0_to_2_10 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  r_fan_ff_lvl_0_to_2_11 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  r_fan_ff_lvl_0_to_2_12 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  r_fan_ff_lvl_0_to_2_13 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  r_fan_ff_lvl_1_to_4_0 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  r_fan_ff_lvl_1_to_4_1 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  r_fan_ff_lvl_1_to_3_0 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  r_fan_ff_lvl_1_to_3_1 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  r_fan_ff_lvl_1_to_3_2 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  r_fan_ff_lvl_1_to_3_3 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  r_fan_ff_lvl_1_to_3_4 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  r_fan_ff_lvl_1_to_3_5 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  r_fan_ff_lvl_2_to_4_0 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  r_fan_ff_lvl_2_to_4_1 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  r_lvl_output_ff_0 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  r_lvl_output_ff_1 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  r_lvl_output_ff_2 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  r_lvl_output_ff_3 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  r_lvl_output_ff_6 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  r_lvl_output_ff_7 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  r_lvl_output_ff_8 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  r_lvl_output_ff_9 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  r_lvl_output_ff_10 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  r_lvl_output_ff_11 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  r_lvl_output_ff_12 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  r_lvl_output_ff_13 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  r_lvl_output_ff_14 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  r_lvl_output_ff_15 = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  r_lvl_output_ff_16 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  r_lvl_output_ff_17 = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  r_lvl_output_ff_18 = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  r_lvl_output_ff_19 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  r_lvl_output_ff_20 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  r_lvl_output_ff_21 = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  r_lvl_output_ff_22 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  r_lvl_output_ff_23 = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  r_lvl_output_ff_24 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  r_lvl_output_ff_25 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  r_lvl_output_ff_26 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  r_lvl_output_ff_27 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  r_lvl_output_ff_28 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  r_lvl_output_ff_29 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  r_lvl_output_ff_30 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  r_lvl_output_ff_31 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  r_lvl_output_ff_32 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  r_lvl_output_ff_33 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  r_lvl_output_ff_34 = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  r_lvl_output_ff_35 = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  r_lvl_output_ff_37 = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  r_lvl_output_ff_38 = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  r_lvl_output_ff_39 = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  r_lvl_output_ff_40 = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  r_lvl_output_ff_41 = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  r_lvl_output_ff_42 = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  r_lvl_output_ff_43 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  r_lvl_output_ff_44 = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  r_lvl_output_ff_45 = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  r_lvl_output_ff_46 = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  r_lvl_output_ff_47 = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  r_lvl_output_ff_48 = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  r_lvl_output_ff_49 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  r_lvl_output_ff_50 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  r_lvl_output_ff_51 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  r_lvl_output_ff_52 = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  r_lvl_output_ff_53 = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  r_lvl_output_ff_54 = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  r_lvl_output_ff_55 = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  r_lvl_output_ff_56 = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  r_lvl_output_ff_57 = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  r_lvl_output_ff_58 = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  r_lvl_output_ff_59 = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  r_lvl_output_ff_60 = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  r_lvl_output_ff_61 = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  r_lvl_output_ff_62 = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  r_lvl_output_ff_63 = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  r_lvl_output_ff_64 = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  r_lvl_output_ff_65 = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  r_lvl_output_ff_66 = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  r_lvl_output_ff_67 = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  r_lvl_output_ff_68 = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  r_lvl_output_ff_69 = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  r_lvl_output_ff_70 = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  r_lvl_output_ff_71 = _RAND_100[31:0];
  _RAND_101 = {1{`RANDOM}};
  r_lvl_output_ff_72 = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  r_lvl_output_ff_73 = _RAND_102[31:0];
  _RAND_103 = {1{`RANDOM}};
  r_lvl_output_ff_74 = _RAND_103[31:0];
  _RAND_104 = {1{`RANDOM}};
  r_lvl_output_ff_75 = _RAND_104[31:0];
  _RAND_105 = {1{`RANDOM}};
  r_lvl_output_ff_76 = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  r_lvl_output_ff_77 = _RAND_106[31:0];
  _RAND_107 = {1{`RANDOM}};
  r_lvl_output_ff_78 = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  r_lvl_output_ff_79 = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  r_lvl_output_ff_80 = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  r_lvl_output_ff_81 = _RAND_110[31:0];
  _RAND_111 = {1{`RANDOM}};
  r_lvl_output_ff_82 = _RAND_111[31:0];
  _RAND_112 = {1{`RANDOM}};
  r_lvl_output_ff_83 = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  r_lvl_output_ff_84 = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  r_lvl_output_ff_85 = _RAND_114[31:0];
  _RAND_115 = {1{`RANDOM}};
  r_lvl_output_ff_86 = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  r_lvl_output_ff_87 = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  r_lvl_output_ff_88 = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  r_lvl_output_ff_89 = _RAND_118[31:0];
  _RAND_119 = {1{`RANDOM}};
  r_lvl_output_ff_90 = _RAND_119[31:0];
  _RAND_120 = {1{`RANDOM}};
  r_lvl_output_ff_91 = _RAND_120[31:0];
  _RAND_121 = {1{`RANDOM}};
  r_lvl_output_ff_92 = _RAND_121[31:0];
  _RAND_122 = {1{`RANDOM}};
  r_lvl_output_ff_93 = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  r_lvl_output_ff_94 = _RAND_123[31:0];
  _RAND_124 = {1{`RANDOM}};
  r_lvl_output_ff_95 = _RAND_124[31:0];
  _RAND_125 = {1{`RANDOM}};
  r_lvl_output_ff_96 = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  r_lvl_output_ff_97 = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  r_lvl_output_ff_98 = _RAND_127[31:0];
  _RAND_128 = {1{`RANDOM}};
  r_lvl_output_ff_99 = _RAND_128[31:0];
  _RAND_129 = {1{`RANDOM}};
  r_lvl_output_ff_100 = _RAND_129[31:0];
  _RAND_130 = {1{`RANDOM}};
  r_lvl_output_ff_101 = _RAND_130[31:0];
  _RAND_131 = {1{`RANDOM}};
  r_lvl_output_ff_102 = _RAND_131[31:0];
  _RAND_132 = {1{`RANDOM}};
  r_lvl_output_ff_103 = _RAND_132[31:0];
  _RAND_133 = {1{`RANDOM}};
  r_lvl_output_ff_104 = _RAND_133[31:0];
  _RAND_134 = {1{`RANDOM}};
  r_lvl_output_ff_105 = _RAND_134[31:0];
  _RAND_135 = {1{`RANDOM}};
  r_lvl_output_ff_106 = _RAND_135[31:0];
  _RAND_136 = {1{`RANDOM}};
  r_lvl_output_ff_107 = _RAND_136[31:0];
  _RAND_137 = {1{`RANDOM}};
  r_lvl_output_ff_108 = _RAND_137[31:0];
  _RAND_138 = {1{`RANDOM}};
  r_lvl_output_ff_109 = _RAND_138[31:0];
  _RAND_139 = {1{`RANDOM}};
  r_lvl_output_ff_110 = _RAND_139[31:0];
  _RAND_140 = {1{`RANDOM}};
  r_lvl_output_ff_112 = _RAND_140[31:0];
  _RAND_141 = {1{`RANDOM}};
  r_lvl_output_ff_113 = _RAND_141[31:0];
  _RAND_142 = {1{`RANDOM}};
  r_lvl_output_ff_114 = _RAND_142[31:0];
  _RAND_143 = {1{`RANDOM}};
  r_lvl_output_ff_115 = _RAND_143[31:0];
  _RAND_144 = {1{`RANDOM}};
  r_lvl_output_ff_116 = _RAND_144[31:0];
  _RAND_145 = {1{`RANDOM}};
  r_lvl_output_ff_117 = _RAND_145[31:0];
  _RAND_146 = {1{`RANDOM}};
  r_lvl_output_ff_118 = _RAND_146[31:0];
  _RAND_147 = {1{`RANDOM}};
  r_lvl_output_ff_119 = _RAND_147[31:0];
  _RAND_148 = {1{`RANDOM}};
  r_lvl_output_ff_120 = _RAND_148[31:0];
  _RAND_149 = {1{`RANDOM}};
  r_lvl_output_ff_121 = _RAND_149[31:0];
  _RAND_150 = {1{`RANDOM}};
  r_lvl_output_ff_122 = _RAND_150[31:0];
  _RAND_151 = {1{`RANDOM}};
  r_lvl_output_ff_123 = _RAND_151[31:0];
  _RAND_152 = {1{`RANDOM}};
  r_lvl_output_ff_124 = _RAND_152[31:0];
  _RAND_153 = {1{`RANDOM}};
  r_lvl_output_ff_125 = _RAND_153[31:0];
  _RAND_154 = {1{`RANDOM}};
  r_lvl_output_ff_126 = _RAND_154[31:0];
  _RAND_155 = {1{`RANDOM}};
  r_lvl_output_ff_127 = _RAND_155[31:0];
  _RAND_156 = {1{`RANDOM}};
  r_lvl_output_ff_128 = _RAND_156[31:0];
  _RAND_157 = {1{`RANDOM}};
  r_lvl_output_ff_129 = _RAND_157[31:0];
  _RAND_158 = {1{`RANDOM}};
  r_lvl_output_ff_130 = _RAND_158[31:0];
  _RAND_159 = {1{`RANDOM}};
  r_lvl_output_ff_131 = _RAND_159[31:0];
  _RAND_160 = {1{`RANDOM}};
  r_lvl_output_ff_132 = _RAND_160[31:0];
  _RAND_161 = {1{`RANDOM}};
  r_lvl_output_ff_133 = _RAND_161[31:0];
  _RAND_162 = {1{`RANDOM}};
  r_lvl_output_ff_134 = _RAND_162[31:0];
  _RAND_163 = {1{`RANDOM}};
  r_lvl_output_ff_135 = _RAND_163[31:0];
  _RAND_164 = {1{`RANDOM}};
  r_lvl_output_ff_136 = _RAND_164[31:0];
  _RAND_165 = {1{`RANDOM}};
  r_lvl_output_ff_137 = _RAND_165[31:0];
  _RAND_166 = {1{`RANDOM}};
  r_lvl_output_ff_138 = _RAND_166[31:0];
  _RAND_167 = {1{`RANDOM}};
  r_lvl_output_ff_139 = _RAND_167[31:0];
  _RAND_168 = {1{`RANDOM}};
  r_lvl_output_ff_140 = _RAND_168[31:0];
  _RAND_169 = {1{`RANDOM}};
  r_lvl_output_ff_141 = _RAND_169[31:0];
  _RAND_170 = {1{`RANDOM}};
  r_lvl_output_ff_142 = _RAND_170[31:0];
  _RAND_171 = {1{`RANDOM}};
  r_lvl_output_ff_143 = _RAND_171[31:0];
  _RAND_172 = {1{`RANDOM}};
  r_lvl_output_ff_144 = _RAND_172[31:0];
  _RAND_173 = {1{`RANDOM}};
  r_lvl_output_ff_145 = _RAND_173[31:0];
  _RAND_174 = {1{`RANDOM}};
  r_lvl_output_ff_146 = _RAND_174[31:0];
  _RAND_175 = {1{`RANDOM}};
  r_lvl_output_ff_147 = _RAND_175[31:0];
  _RAND_176 = {1{`RANDOM}};
  r_lvl_output_ff_148 = _RAND_176[31:0];
  _RAND_177 = {1{`RANDOM}};
  r_lvl_output_ff_149 = _RAND_177[31:0];
  _RAND_178 = {1{`RANDOM}};
  r_lvl_output_ff_150 = _RAND_178[31:0];
  _RAND_179 = {1{`RANDOM}};
  r_lvl_output_ff_151 = _RAND_179[31:0];
  _RAND_180 = {1{`RANDOM}};
  r_lvl_output_ff_152 = _RAND_180[31:0];
  _RAND_181 = {1{`RANDOM}};
  r_lvl_output_ff_153 = _RAND_181[31:0];
  _RAND_182 = {1{`RANDOM}};
  r_lvl_output_ff_154 = _RAND_182[31:0];
  _RAND_183 = {1{`RANDOM}};
  r_lvl_output_ff_155 = _RAND_183[31:0];
  _RAND_184 = {1{`RANDOM}};
  r_lvl_output_ff_156 = _RAND_184[31:0];
  _RAND_185 = {1{`RANDOM}};
  r_lvl_output_ff_157 = _RAND_185[31:0];
  _RAND_186 = {1{`RANDOM}};
  r_lvl_output_ff_158 = _RAND_186[31:0];
  _RAND_187 = {1{`RANDOM}};
  r_lvl_output_ff_159 = _RAND_187[31:0];
  _RAND_188 = {1{`RANDOM}};
  r_lvl_output_ff_valid_0 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  r_lvl_output_ff_valid_1 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  r_lvl_output_ff_valid_2 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  r_lvl_output_ff_valid_3 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  r_lvl_output_ff_valid_4 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  r_lvl_output_ff_valid_5 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  r_lvl_output_ff_valid_6 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  r_lvl_output_ff_valid_7 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  r_lvl_output_ff_valid_8 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  r_lvl_output_ff_valid_9 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  r_lvl_output_ff_valid_10 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  r_lvl_output_ff_valid_11 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  r_lvl_output_ff_valid_12 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  r_lvl_output_ff_valid_13 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  r_lvl_output_ff_valid_14 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  r_lvl_output_ff_valid_15 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  r_lvl_output_ff_valid_16 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  r_lvl_output_ff_valid_17 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  r_lvl_output_ff_valid_18 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  r_lvl_output_ff_valid_19 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  r_lvl_output_ff_valid_20 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  r_lvl_output_ff_valid_21 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  r_lvl_output_ff_valid_22 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  r_lvl_output_ff_valid_23 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  r_lvl_output_ff_valid_24 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  r_lvl_output_ff_valid_25 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  r_lvl_output_ff_valid_26 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  r_lvl_output_ff_valid_27 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  r_lvl_output_ff_valid_28 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  r_lvl_output_ff_valid_29 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  r_lvl_output_ff_valid_30 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  r_lvl_output_ff_valid_31 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  r_lvl_output_ff_valid_32 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  r_lvl_output_ff_valid_33 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  r_lvl_output_ff_valid_34 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  r_lvl_output_ff_valid_35 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  r_lvl_output_ff_valid_36 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  r_lvl_output_ff_valid_37 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  r_lvl_output_ff_valid_38 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  r_lvl_output_ff_valid_39 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  r_lvl_output_ff_valid_40 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  r_lvl_output_ff_valid_41 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  r_lvl_output_ff_valid_42 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  r_lvl_output_ff_valid_43 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  r_lvl_output_ff_valid_44 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  r_lvl_output_ff_valid_45 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  r_lvl_output_ff_valid_46 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  r_lvl_output_ff_valid_47 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  r_lvl_output_ff_valid_48 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  r_lvl_output_ff_valid_49 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  r_lvl_output_ff_valid_50 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  r_lvl_output_ff_valid_51 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  r_lvl_output_ff_valid_52 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  r_lvl_output_ff_valid_53 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  r_lvl_output_ff_valid_54 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  r_lvl_output_ff_valid_55 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  r_lvl_output_ff_valid_56 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  r_lvl_output_ff_valid_57 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  r_lvl_output_ff_valid_58 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  r_lvl_output_ff_valid_59 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  r_lvl_output_ff_valid_60 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  r_lvl_output_ff_valid_61 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  r_lvl_output_ff_valid_62 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  r_lvl_output_ff_valid_63 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  r_lvl_output_ff_valid_64 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  r_lvl_output_ff_valid_65 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  r_lvl_output_ff_valid_66 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  r_lvl_output_ff_valid_67 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  r_lvl_output_ff_valid_68 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  r_lvl_output_ff_valid_69 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  r_lvl_output_ff_valid_70 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  r_lvl_output_ff_valid_71 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  r_lvl_output_ff_valid_72 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  r_lvl_output_ff_valid_73 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  r_lvl_output_ff_valid_74 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  r_lvl_output_ff_valid_75 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  r_lvl_output_ff_valid_76 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  r_lvl_output_ff_valid_77 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  r_lvl_output_ff_valid_78 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  r_lvl_output_ff_valid_79 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  r_lvl_output_ff_valid_80 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  r_lvl_output_ff_valid_81 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  r_lvl_output_ff_valid_82 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  r_lvl_output_ff_valid_83 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  r_lvl_output_ff_valid_84 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  r_lvl_output_ff_valid_85 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  r_lvl_output_ff_valid_86 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  r_lvl_output_ff_valid_87 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  r_lvl_output_ff_valid_88 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  r_lvl_output_ff_valid_89 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  r_lvl_output_ff_valid_90 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  r_lvl_output_ff_valid_91 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  r_lvl_output_ff_valid_92 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  r_lvl_output_ff_valid_93 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  r_lvl_output_ff_valid_94 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  r_lvl_output_ff_valid_95 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  r_lvl_output_ff_valid_96 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  r_lvl_output_ff_valid_97 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  r_lvl_output_ff_valid_98 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  r_lvl_output_ff_valid_99 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  r_lvl_output_ff_valid_100 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  r_lvl_output_ff_valid_101 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  r_lvl_output_ff_valid_102 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  r_lvl_output_ff_valid_103 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  r_lvl_output_ff_valid_104 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  r_lvl_output_ff_valid_105 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  r_lvl_output_ff_valid_106 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  r_lvl_output_ff_valid_107 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  r_lvl_output_ff_valid_108 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  r_lvl_output_ff_valid_109 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  r_lvl_output_ff_valid_110 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  r_lvl_output_ff_valid_111 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  r_lvl_output_ff_valid_112 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  r_lvl_output_ff_valid_113 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  r_lvl_output_ff_valid_114 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  r_lvl_output_ff_valid_115 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  r_lvl_output_ff_valid_116 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  r_lvl_output_ff_valid_117 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  r_lvl_output_ff_valid_118 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  r_lvl_output_ff_valid_119 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  r_lvl_output_ff_valid_120 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  r_lvl_output_ff_valid_121 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  r_lvl_output_ff_valid_122 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  r_lvl_output_ff_valid_123 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  r_lvl_output_ff_valid_124 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  r_lvl_output_ff_valid_125 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  r_lvl_output_ff_valid_126 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  r_lvl_output_ff_valid_127 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  r_lvl_output_ff_valid_128 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  r_lvl_output_ff_valid_129 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  r_lvl_output_ff_valid_130 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  r_lvl_output_ff_valid_131 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  r_lvl_output_ff_valid_132 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  r_lvl_output_ff_valid_133 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  r_lvl_output_ff_valid_134 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  r_lvl_output_ff_valid_135 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  r_lvl_output_ff_valid_136 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  r_lvl_output_ff_valid_137 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  r_lvl_output_ff_valid_138 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  r_lvl_output_ff_valid_139 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  r_lvl_output_ff_valid_140 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  r_lvl_output_ff_valid_141 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  r_lvl_output_ff_valid_142 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  r_lvl_output_ff_valid_143 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  r_lvl_output_ff_valid_144 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  r_lvl_output_ff_valid_145 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  r_lvl_output_ff_valid_146 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  r_lvl_output_ff_valid_147 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  r_lvl_output_ff_valid_148 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  r_lvl_output_ff_valid_149 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  r_lvl_output_ff_valid_150 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  r_lvl_output_ff_valid_151 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  r_lvl_output_ff_valid_152 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  r_lvl_output_ff_valid_153 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  r_lvl_output_ff_valid_154 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  r_lvl_output_ff_valid_155 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  r_lvl_output_ff_valid_156 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  r_lvl_output_ff_valid_157 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  r_lvl_output_ff_valid_158 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  r_lvl_output_ff_valid_159 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  r_valid_0 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  r_valid_1 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  r_valid_2 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  r_valid_3 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  r_valid_4 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  r_final_sum = _RAND_353[31:0];
  _RAND_354 = {1{`RANDOM}};
  r_final_add = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  r_final_add2 = _RAND_355[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
