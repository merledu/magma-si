module Muxes(
  input         clock,
  input         reset,
  input  [15:0] io_mat1_0_0,
  input  [15:0] io_mat1_0_1,
  input  [15:0] io_mat1_0_2,
  input  [15:0] io_mat1_0_3,
  input  [15:0] io_mat1_0_4,
  input  [15:0] io_mat1_0_5,
  input  [15:0] io_mat1_0_6,
  input  [15:0] io_mat1_0_7,
  input  [15:0] io_mat1_1_0,
  input  [15:0] io_mat1_1_1,
  input  [15:0] io_mat1_1_2,
  input  [15:0] io_mat1_1_3,
  input  [15:0] io_mat1_1_4,
  input  [15:0] io_mat1_1_5,
  input  [15:0] io_mat1_1_6,
  input  [15:0] io_mat1_1_7,
  input  [15:0] io_mat1_2_0,
  input  [15:0] io_mat1_2_1,
  input  [15:0] io_mat1_2_2,
  input  [15:0] io_mat1_2_3,
  input  [15:0] io_mat1_2_4,
  input  [15:0] io_mat1_2_5,
  input  [15:0] io_mat1_2_6,
  input  [15:0] io_mat1_2_7,
  input  [15:0] io_mat1_3_0,
  input  [15:0] io_mat1_3_1,
  input  [15:0] io_mat1_3_2,
  input  [15:0] io_mat1_3_3,
  input  [15:0] io_mat1_3_4,
  input  [15:0] io_mat1_3_5,
  input  [15:0] io_mat1_3_6,
  input  [15:0] io_mat1_3_7,
  input  [15:0] io_mat1_4_0,
  input  [15:0] io_mat1_4_1,
  input  [15:0] io_mat1_4_2,
  input  [15:0] io_mat1_4_3,
  input  [15:0] io_mat1_4_4,
  input  [15:0] io_mat1_4_5,
  input  [15:0] io_mat1_4_6,
  input  [15:0] io_mat1_4_7,
  input  [15:0] io_mat1_5_0,
  input  [15:0] io_mat1_5_1,
  input  [15:0] io_mat1_5_2,
  input  [15:0] io_mat1_5_3,
  input  [15:0] io_mat1_5_4,
  input  [15:0] io_mat1_5_5,
  input  [15:0] io_mat1_5_6,
  input  [15:0] io_mat1_5_7,
  input  [15:0] io_mat1_6_0,
  input  [15:0] io_mat1_6_1,
  input  [15:0] io_mat1_6_2,
  input  [15:0] io_mat1_6_3,
  input  [15:0] io_mat1_6_4,
  input  [15:0] io_mat1_6_5,
  input  [15:0] io_mat1_6_6,
  input  [15:0] io_mat1_6_7,
  input  [15:0] io_mat1_7_0,
  input  [15:0] io_mat1_7_1,
  input  [15:0] io_mat1_7_2,
  input  [15:0] io_mat1_7_3,
  input  [15:0] io_mat1_7_4,
  input  [15:0] io_mat1_7_5,
  input  [15:0] io_mat1_7_6,
  input  [15:0] io_mat1_7_7,
  input  [15:0] io_mat2_0,
  input  [15:0] io_mat2_1,
  input  [15:0] io_mat2_2,
  input  [15:0] io_mat2_3,
  input  [15:0] io_mat2_4,
  input  [15:0] io_mat2_5,
  input  [15:0] io_mat2_6,
  input  [15:0] io_mat2_7,
  input  [15:0] io_counterMatrix1_0_0,
  input  [15:0] io_counterMatrix1_0_1,
  input  [15:0] io_counterMatrix1_0_2,
  input  [15:0] io_counterMatrix1_0_3,
  input  [15:0] io_counterMatrix1_0_4,
  input  [15:0] io_counterMatrix1_0_5,
  input  [15:0] io_counterMatrix1_0_6,
  input  [15:0] io_counterMatrix1_0_7,
  input  [15:0] io_counterMatrix1_1_0,
  input  [15:0] io_counterMatrix1_1_1,
  input  [15:0] io_counterMatrix1_1_2,
  input  [15:0] io_counterMatrix1_1_3,
  input  [15:0] io_counterMatrix1_1_4,
  input  [15:0] io_counterMatrix1_1_5,
  input  [15:0] io_counterMatrix1_1_6,
  input  [15:0] io_counterMatrix1_1_7,
  input  [15:0] io_counterMatrix1_2_0,
  input  [15:0] io_counterMatrix1_2_1,
  input  [15:0] io_counterMatrix1_2_2,
  input  [15:0] io_counterMatrix1_2_3,
  input  [15:0] io_counterMatrix1_2_4,
  input  [15:0] io_counterMatrix1_2_5,
  input  [15:0] io_counterMatrix1_2_6,
  input  [15:0] io_counterMatrix1_2_7,
  input  [15:0] io_counterMatrix1_3_0,
  input  [15:0] io_counterMatrix1_3_1,
  input  [15:0] io_counterMatrix1_3_2,
  input  [15:0] io_counterMatrix1_3_3,
  input  [15:0] io_counterMatrix1_3_4,
  input  [15:0] io_counterMatrix1_3_5,
  input  [15:0] io_counterMatrix1_3_6,
  input  [15:0] io_counterMatrix1_3_7,
  input  [15:0] io_counterMatrix1_4_0,
  input  [15:0] io_counterMatrix1_4_1,
  input  [15:0] io_counterMatrix1_4_2,
  input  [15:0] io_counterMatrix1_4_3,
  input  [15:0] io_counterMatrix1_4_4,
  input  [15:0] io_counterMatrix1_4_5,
  input  [15:0] io_counterMatrix1_4_6,
  input  [15:0] io_counterMatrix1_4_7,
  input  [15:0] io_counterMatrix1_5_0,
  input  [15:0] io_counterMatrix1_5_1,
  input  [15:0] io_counterMatrix1_5_2,
  input  [15:0] io_counterMatrix1_5_3,
  input  [15:0] io_counterMatrix1_5_4,
  input  [15:0] io_counterMatrix1_5_5,
  input  [15:0] io_counterMatrix1_5_6,
  input  [15:0] io_counterMatrix1_5_7,
  input  [15:0] io_counterMatrix1_6_0,
  input  [15:0] io_counterMatrix1_6_1,
  input  [15:0] io_counterMatrix1_6_2,
  input  [15:0] io_counterMatrix1_6_3,
  input  [15:0] io_counterMatrix1_6_4,
  input  [15:0] io_counterMatrix1_6_5,
  input  [15:0] io_counterMatrix1_6_6,
  input  [15:0] io_counterMatrix1_6_7,
  input  [15:0] io_counterMatrix1_7_0,
  input  [15:0] io_counterMatrix1_7_1,
  input  [15:0] io_counterMatrix1_7_2,
  input  [15:0] io_counterMatrix1_7_3,
  input  [15:0] io_counterMatrix1_7_4,
  input  [15:0] io_counterMatrix1_7_5,
  input  [15:0] io_counterMatrix1_7_6,
  input  [15:0] io_counterMatrix1_7_7,
  input  [15:0] io_counterMatrix2_0,
  input  [15:0] io_counterMatrix2_1,
  input  [15:0] io_counterMatrix2_2,
  input  [15:0] io_counterMatrix2_3,
  input  [15:0] io_counterMatrix2_4,
  input  [15:0] io_counterMatrix2_5,
  input  [15:0] io_counterMatrix2_6,
  input  [15:0] io_counterMatrix2_7,
  output [3:0]  io_i_mux_bus_0,
  output [3:0]  io_i_mux_bus_1,
  output [3:0]  io_i_mux_bus_2,
  output [3:0]  io_i_mux_bus_3,
  output [15:0] io_Source_0,
  output [15:0] io_Source_1,
  output [15:0] io_Source_2,
  output [15:0] io_Source_3,
  output [15:0] io_destination_0,
  output [15:0] io_destination_1,
  output [15:0] io_destination_2,
  output [15:0] io_destination_3,
  output        io_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
`endif // RANDOMIZE_REG_INIT
  reg [15:0] prevStationary_matrix_0_0; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_0_1; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_0_2; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_0_3; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_0_4; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_0_5; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_0_6; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_0_7; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_1_0; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_1_1; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_1_2; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_1_3; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_1_4; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_1_5; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_1_6; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_1_7; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_2_0; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_2_1; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_2_2; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_2_3; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_2_4; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_2_5; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_2_6; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_2_7; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_3_0; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_3_1; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_3_2; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_3_3; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_3_4; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_3_5; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_3_6; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_3_7; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_4_0; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_4_1; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_4_2; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_4_3; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_4_4; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_4_5; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_4_6; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_4_7; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_5_0; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_5_1; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_5_2; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_5_3; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_5_4; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_5_5; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_5_6; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_5_7; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_6_0; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_6_1; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_6_2; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_6_3; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_6_4; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_6_5; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_6_6; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_6_7; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_7_0; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_7_1; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_7_2; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_7_3; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_7_4; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_7_5; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_7_6; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_7_7; // @[Muxes.scala 19:40]
  reg [15:0] prevStreaming_matrix_0; // @[Muxes.scala 20:39]
  reg [15:0] prevStreaming_matrix_1; // @[Muxes.scala 20:39]
  reg [15:0] prevStreaming_matrix_2; // @[Muxes.scala 20:39]
  reg [15:0] prevStreaming_matrix_3; // @[Muxes.scala 20:39]
  reg [15:0] prevStreaming_matrix_4; // @[Muxes.scala 20:39]
  reg [15:0] prevStreaming_matrix_5; // @[Muxes.scala 20:39]
  reg [15:0] prevStreaming_matrix_6; // @[Muxes.scala 20:39]
  reg [15:0] prevStreaming_matrix_7; // @[Muxes.scala 20:39]
  reg  matricesAreEqual; // @[Muxes.scala 21:31]
  reg  jValid; // @[Muxes.scala 27:25]
  reg [31:0] i; // @[Muxes.scala 28:20]
  reg [31:0] j; // @[Muxes.scala 29:20]
  reg [31:0] k; // @[Muxes.scala 30:20]
  reg [31:0] counter; // @[Muxes.scala 31:26]
  reg [3:0] mux_0; // @[Muxes.scala 32:22]
  reg [3:0] mux_1; // @[Muxes.scala 32:22]
  reg [3:0] mux_2; // @[Muxes.scala 32:22]
  reg [3:0] mux_3; // @[Muxes.scala 32:22]
  reg [3:0] mux_4; // @[Muxes.scala 32:22]
  reg [3:0] mux_5; // @[Muxes.scala 32:22]
  reg [3:0] mux_6; // @[Muxes.scala 32:22]
  reg [3:0] mux_7; // @[Muxes.scala 32:22]
  reg [3:0] mux_8; // @[Muxes.scala 32:22]
  reg [3:0] mux_9; // @[Muxes.scala 32:22]
  reg [3:0] mux_10; // @[Muxes.scala 32:22]
  reg [3:0] mux_11; // @[Muxes.scala 32:22]
  reg [3:0] mux_12; // @[Muxes.scala 32:22]
  reg [3:0] mux_13; // @[Muxes.scala 32:22]
  reg [3:0] mux_14; // @[Muxes.scala 32:22]
  reg [3:0] mux_15; // @[Muxes.scala 32:22]
  reg [3:0] mux_16; // @[Muxes.scala 32:22]
  reg [3:0] mux_17; // @[Muxes.scala 32:22]
  reg [3:0] mux_18; // @[Muxes.scala 32:22]
  reg [3:0] mux_19; // @[Muxes.scala 32:22]
  reg [3:0] mux_20; // @[Muxes.scala 32:22]
  reg [3:0] mux_21; // @[Muxes.scala 32:22]
  reg [3:0] mux_22; // @[Muxes.scala 32:22]
  reg [3:0] mux_23; // @[Muxes.scala 32:22]
  reg [3:0] mux_24; // @[Muxes.scala 32:22]
  reg [3:0] mux_25; // @[Muxes.scala 32:22]
  reg [3:0] mux_26; // @[Muxes.scala 32:22]
  reg [3:0] mux_27; // @[Muxes.scala 32:22]
  reg [3:0] mux_28; // @[Muxes.scala 32:22]
  reg [3:0] mux_29; // @[Muxes.scala 32:22]
  reg [3:0] mux_30; // @[Muxes.scala 32:22]
  reg [3:0] mux_31; // @[Muxes.scala 32:22]
  reg [3:0] mux_32; // @[Muxes.scala 32:22]
  reg [3:0] mux_33; // @[Muxes.scala 32:22]
  reg [3:0] mux_34; // @[Muxes.scala 32:22]
  reg [3:0] mux_35; // @[Muxes.scala 32:22]
  reg [3:0] mux_36; // @[Muxes.scala 32:22]
  reg [3:0] mux_37; // @[Muxes.scala 32:22]
  reg [3:0] mux_38; // @[Muxes.scala 32:22]
  reg [3:0] mux_39; // @[Muxes.scala 32:22]
  reg [3:0] mux_40; // @[Muxes.scala 32:22]
  reg [3:0] mux_41; // @[Muxes.scala 32:22]
  reg [3:0] mux_42; // @[Muxes.scala 32:22]
  reg [3:0] mux_43; // @[Muxes.scala 32:22]
  reg [3:0] mux_44; // @[Muxes.scala 32:22]
  reg [3:0] mux_45; // @[Muxes.scala 32:22]
  reg [3:0] mux_46; // @[Muxes.scala 32:22]
  reg [3:0] mux_47; // @[Muxes.scala 32:22]
  reg [3:0] mux_48; // @[Muxes.scala 32:22]
  reg [3:0] mux_49; // @[Muxes.scala 32:22]
  reg [3:0] mux_50; // @[Muxes.scala 32:22]
  reg [3:0] mux_51; // @[Muxes.scala 32:22]
  reg [3:0] mux_52; // @[Muxes.scala 32:22]
  reg [3:0] mux_53; // @[Muxes.scala 32:22]
  reg [3:0] mux_54; // @[Muxes.scala 32:22]
  reg [3:0] mux_55; // @[Muxes.scala 32:22]
  reg [3:0] mux_56; // @[Muxes.scala 32:22]
  reg [3:0] mux_57; // @[Muxes.scala 32:22]
  reg [3:0] mux_58; // @[Muxes.scala 32:22]
  reg [3:0] mux_59; // @[Muxes.scala 32:22]
  reg [3:0] mux_60; // @[Muxes.scala 32:22]
  reg [3:0] mux_61; // @[Muxes.scala 32:22]
  reg [3:0] mux_62; // @[Muxes.scala 32:22]
  reg [3:0] mux_63; // @[Muxes.scala 32:22]
  reg [15:0] src_0; // @[Muxes.scala 33:22]
  reg [15:0] src_1; // @[Muxes.scala 33:22]
  reg [15:0] src_2; // @[Muxes.scala 33:22]
  reg [15:0] src_3; // @[Muxes.scala 33:22]
  reg [15:0] src_4; // @[Muxes.scala 33:22]
  reg [15:0] src_5; // @[Muxes.scala 33:22]
  reg [15:0] src_6; // @[Muxes.scala 33:22]
  reg [15:0] src_7; // @[Muxes.scala 33:22]
  reg [15:0] src_8; // @[Muxes.scala 33:22]
  reg [15:0] src_9; // @[Muxes.scala 33:22]
  reg [15:0] src_10; // @[Muxes.scala 33:22]
  reg [15:0] src_11; // @[Muxes.scala 33:22]
  reg [15:0] src_12; // @[Muxes.scala 33:22]
  reg [15:0] src_13; // @[Muxes.scala 33:22]
  reg [15:0] src_14; // @[Muxes.scala 33:22]
  reg [15:0] src_15; // @[Muxes.scala 33:22]
  reg [15:0] src_16; // @[Muxes.scala 33:22]
  reg [15:0] src_17; // @[Muxes.scala 33:22]
  reg [15:0] src_18; // @[Muxes.scala 33:22]
  reg [15:0] src_19; // @[Muxes.scala 33:22]
  reg [15:0] src_20; // @[Muxes.scala 33:22]
  reg [15:0] src_21; // @[Muxes.scala 33:22]
  reg [15:0] src_22; // @[Muxes.scala 33:22]
  reg [15:0] src_23; // @[Muxes.scala 33:22]
  reg [15:0] src_24; // @[Muxes.scala 33:22]
  reg [15:0] src_25; // @[Muxes.scala 33:22]
  reg [15:0] src_26; // @[Muxes.scala 33:22]
  reg [15:0] src_27; // @[Muxes.scala 33:22]
  reg [15:0] src_28; // @[Muxes.scala 33:22]
  reg [15:0] src_29; // @[Muxes.scala 33:22]
  reg [15:0] src_30; // @[Muxes.scala 33:22]
  reg [15:0] src_31; // @[Muxes.scala 33:22]
  reg [15:0] src_32; // @[Muxes.scala 33:22]
  reg [15:0] src_33; // @[Muxes.scala 33:22]
  reg [15:0] src_34; // @[Muxes.scala 33:22]
  reg [15:0] src_35; // @[Muxes.scala 33:22]
  reg [15:0] src_36; // @[Muxes.scala 33:22]
  reg [15:0] src_37; // @[Muxes.scala 33:22]
  reg [15:0] src_38; // @[Muxes.scala 33:22]
  reg [15:0] src_39; // @[Muxes.scala 33:22]
  reg [15:0] src_40; // @[Muxes.scala 33:22]
  reg [15:0] src_41; // @[Muxes.scala 33:22]
  reg [15:0] src_42; // @[Muxes.scala 33:22]
  reg [15:0] src_43; // @[Muxes.scala 33:22]
  reg [15:0] src_44; // @[Muxes.scala 33:22]
  reg [15:0] src_45; // @[Muxes.scala 33:22]
  reg [15:0] src_46; // @[Muxes.scala 33:22]
  reg [15:0] src_47; // @[Muxes.scala 33:22]
  reg [15:0] src_48; // @[Muxes.scala 33:22]
  reg [15:0] src_49; // @[Muxes.scala 33:22]
  reg [15:0] src_50; // @[Muxes.scala 33:22]
  reg [15:0] src_51; // @[Muxes.scala 33:22]
  reg [15:0] src_52; // @[Muxes.scala 33:22]
  reg [15:0] src_53; // @[Muxes.scala 33:22]
  reg [15:0] src_54; // @[Muxes.scala 33:22]
  reg [15:0] src_55; // @[Muxes.scala 33:22]
  reg [15:0] src_56; // @[Muxes.scala 33:22]
  reg [15:0] src_57; // @[Muxes.scala 33:22]
  reg [15:0] src_58; // @[Muxes.scala 33:22]
  reg [15:0] src_59; // @[Muxes.scala 33:22]
  reg [15:0] src_60; // @[Muxes.scala 33:22]
  reg [15:0] src_61; // @[Muxes.scala 33:22]
  reg [15:0] src_62; // @[Muxes.scala 33:22]
  reg [15:0] src_63; // @[Muxes.scala 33:22]
  reg [15:0] dest_0; // @[Muxes.scala 34:23]
  reg [15:0] dest_1; // @[Muxes.scala 34:23]
  reg [15:0] dest_2; // @[Muxes.scala 34:23]
  reg [15:0] dest_3; // @[Muxes.scala 34:23]
  reg [15:0] dest_4; // @[Muxes.scala 34:23]
  reg [15:0] dest_5; // @[Muxes.scala 34:23]
  reg [15:0] dest_6; // @[Muxes.scala 34:23]
  reg [15:0] dest_7; // @[Muxes.scala 34:23]
  reg [15:0] dest_8; // @[Muxes.scala 34:23]
  reg [15:0] dest_9; // @[Muxes.scala 34:23]
  reg [15:0] dest_10; // @[Muxes.scala 34:23]
  reg [15:0] dest_11; // @[Muxes.scala 34:23]
  reg [15:0] dest_12; // @[Muxes.scala 34:23]
  reg [15:0] dest_13; // @[Muxes.scala 34:23]
  reg [15:0] dest_14; // @[Muxes.scala 34:23]
  reg [15:0] dest_15; // @[Muxes.scala 34:23]
  reg [15:0] dest_16; // @[Muxes.scala 34:23]
  reg [15:0] dest_17; // @[Muxes.scala 34:23]
  reg [15:0] dest_18; // @[Muxes.scala 34:23]
  reg [15:0] dest_19; // @[Muxes.scala 34:23]
  reg [15:0] dest_20; // @[Muxes.scala 34:23]
  reg [15:0] dest_21; // @[Muxes.scala 34:23]
  reg [15:0] dest_22; // @[Muxes.scala 34:23]
  reg [15:0] dest_23; // @[Muxes.scala 34:23]
  reg [15:0] dest_24; // @[Muxes.scala 34:23]
  reg [15:0] dest_25; // @[Muxes.scala 34:23]
  reg [15:0] dest_26; // @[Muxes.scala 34:23]
  reg [15:0] dest_27; // @[Muxes.scala 34:23]
  reg [15:0] dest_28; // @[Muxes.scala 34:23]
  reg [15:0] dest_29; // @[Muxes.scala 34:23]
  reg [15:0] dest_30; // @[Muxes.scala 34:23]
  reg [15:0] dest_31; // @[Muxes.scala 34:23]
  reg [15:0] dest_32; // @[Muxes.scala 34:23]
  reg [15:0] dest_33; // @[Muxes.scala 34:23]
  reg [15:0] dest_34; // @[Muxes.scala 34:23]
  reg [15:0] dest_35; // @[Muxes.scala 34:23]
  reg [15:0] dest_36; // @[Muxes.scala 34:23]
  reg [15:0] dest_37; // @[Muxes.scala 34:23]
  reg [15:0] dest_38; // @[Muxes.scala 34:23]
  reg [15:0] dest_39; // @[Muxes.scala 34:23]
  reg [15:0] dest_40; // @[Muxes.scala 34:23]
  reg [15:0] dest_41; // @[Muxes.scala 34:23]
  reg [15:0] dest_42; // @[Muxes.scala 34:23]
  reg [15:0] dest_43; // @[Muxes.scala 34:23]
  reg [15:0] dest_44; // @[Muxes.scala 34:23]
  reg [15:0] dest_45; // @[Muxes.scala 34:23]
  reg [15:0] dest_46; // @[Muxes.scala 34:23]
  reg [15:0] dest_47; // @[Muxes.scala 34:23]
  reg [15:0] dest_48; // @[Muxes.scala 34:23]
  reg [15:0] dest_49; // @[Muxes.scala 34:23]
  reg [15:0] dest_50; // @[Muxes.scala 34:23]
  reg [15:0] dest_51; // @[Muxes.scala 34:23]
  reg [15:0] dest_52; // @[Muxes.scala 34:23]
  reg [15:0] dest_53; // @[Muxes.scala 34:23]
  reg [15:0] dest_54; // @[Muxes.scala 34:23]
  reg [15:0] dest_55; // @[Muxes.scala 34:23]
  reg [15:0] dest_56; // @[Muxes.scala 34:23]
  reg [15:0] dest_57; // @[Muxes.scala 34:23]
  reg [15:0] dest_58; // @[Muxes.scala 34:23]
  reg [15:0] dest_59; // @[Muxes.scala 34:23]
  reg [15:0] dest_60; // @[Muxes.scala 34:23]
  reg [15:0] dest_61; // @[Muxes.scala 34:23]
  reg [15:0] dest_62; // @[Muxes.scala 34:23]
  reg [15:0] dest_63; // @[Muxes.scala 34:23]
  wire  _GEN_0 = io_mat1_0_0 != prevStationary_matrix_0_0 ? 1'h0 : 1'h1; // @[Muxes.scala 22:22 45:61 46:28]
  wire  _GEN_1 = io_mat1_0_1 != prevStationary_matrix_0_1 ? 1'h0 : _GEN_0; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_2 = io_mat1_0_2 != prevStationary_matrix_0_2 ? 1'h0 : _GEN_1; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_3 = io_mat1_0_3 != prevStationary_matrix_0_3 ? 1'h0 : _GEN_2; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_4 = io_mat1_0_4 != prevStationary_matrix_0_4 ? 1'h0 : _GEN_3; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_5 = io_mat1_0_5 != prevStationary_matrix_0_5 ? 1'h0 : _GEN_4; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_6 = io_mat1_0_6 != prevStationary_matrix_0_6 ? 1'h0 : _GEN_5; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_7 = io_mat1_0_7 != prevStationary_matrix_0_7 ? 1'h0 : _GEN_6; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_8 = io_mat2_0 != prevStreaming_matrix_0 ? 1'h0 : _GEN_7; // @[Muxes.scala 49:51 50:26]
  wire  _GEN_9 = io_mat1_1_0 != prevStationary_matrix_1_0 ? 1'h0 : _GEN_8; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_10 = io_mat1_1_1 != prevStationary_matrix_1_1 ? 1'h0 : _GEN_9; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_11 = io_mat1_1_2 != prevStationary_matrix_1_2 ? 1'h0 : _GEN_10; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_12 = io_mat1_1_3 != prevStationary_matrix_1_3 ? 1'h0 : _GEN_11; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_13 = io_mat1_1_4 != prevStationary_matrix_1_4 ? 1'h0 : _GEN_12; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_14 = io_mat1_1_5 != prevStationary_matrix_1_5 ? 1'h0 : _GEN_13; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_15 = io_mat1_1_6 != prevStationary_matrix_1_6 ? 1'h0 : _GEN_14; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_16 = io_mat1_1_7 != prevStationary_matrix_1_7 ? 1'h0 : _GEN_15; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_17 = io_mat2_1 != prevStreaming_matrix_1 ? 1'h0 : _GEN_16; // @[Muxes.scala 49:51 50:26]
  wire  _GEN_18 = io_mat1_2_0 != prevStationary_matrix_2_0 ? 1'h0 : _GEN_17; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_19 = io_mat1_2_1 != prevStationary_matrix_2_1 ? 1'h0 : _GEN_18; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_20 = io_mat1_2_2 != prevStationary_matrix_2_2 ? 1'h0 : _GEN_19; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_21 = io_mat1_2_3 != prevStationary_matrix_2_3 ? 1'h0 : _GEN_20; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_22 = io_mat1_2_4 != prevStationary_matrix_2_4 ? 1'h0 : _GEN_21; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_23 = io_mat1_2_5 != prevStationary_matrix_2_5 ? 1'h0 : _GEN_22; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_24 = io_mat1_2_6 != prevStationary_matrix_2_6 ? 1'h0 : _GEN_23; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_25 = io_mat1_2_7 != prevStationary_matrix_2_7 ? 1'h0 : _GEN_24; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_26 = io_mat2_2 != prevStreaming_matrix_2 ? 1'h0 : _GEN_25; // @[Muxes.scala 49:51 50:26]
  wire  _GEN_27 = io_mat1_3_0 != prevStationary_matrix_3_0 ? 1'h0 : _GEN_26; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_28 = io_mat1_3_1 != prevStationary_matrix_3_1 ? 1'h0 : _GEN_27; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_29 = io_mat1_3_2 != prevStationary_matrix_3_2 ? 1'h0 : _GEN_28; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_30 = io_mat1_3_3 != prevStationary_matrix_3_3 ? 1'h0 : _GEN_29; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_31 = io_mat1_3_4 != prevStationary_matrix_3_4 ? 1'h0 : _GEN_30; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_32 = io_mat1_3_5 != prevStationary_matrix_3_5 ? 1'h0 : _GEN_31; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_33 = io_mat1_3_6 != prevStationary_matrix_3_6 ? 1'h0 : _GEN_32; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_34 = io_mat1_3_7 != prevStationary_matrix_3_7 ? 1'h0 : _GEN_33; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_35 = io_mat2_3 != prevStreaming_matrix_3 ? 1'h0 : _GEN_34; // @[Muxes.scala 49:51 50:26]
  wire  _GEN_36 = io_mat1_4_0 != prevStationary_matrix_4_0 ? 1'h0 : _GEN_35; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_37 = io_mat1_4_1 != prevStationary_matrix_4_1 ? 1'h0 : _GEN_36; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_38 = io_mat1_4_2 != prevStationary_matrix_4_2 ? 1'h0 : _GEN_37; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_39 = io_mat1_4_3 != prevStationary_matrix_4_3 ? 1'h0 : _GEN_38; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_40 = io_mat1_4_4 != prevStationary_matrix_4_4 ? 1'h0 : _GEN_39; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_41 = io_mat1_4_5 != prevStationary_matrix_4_5 ? 1'h0 : _GEN_40; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_42 = io_mat1_4_6 != prevStationary_matrix_4_6 ? 1'h0 : _GEN_41; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_43 = io_mat1_4_7 != prevStationary_matrix_4_7 ? 1'h0 : _GEN_42; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_44 = io_mat2_4 != prevStreaming_matrix_4 ? 1'h0 : _GEN_43; // @[Muxes.scala 49:51 50:26]
  wire  _GEN_45 = io_mat1_5_0 != prevStationary_matrix_5_0 ? 1'h0 : _GEN_44; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_46 = io_mat1_5_1 != prevStationary_matrix_5_1 ? 1'h0 : _GEN_45; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_47 = io_mat1_5_2 != prevStationary_matrix_5_2 ? 1'h0 : _GEN_46; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_48 = io_mat1_5_3 != prevStationary_matrix_5_3 ? 1'h0 : _GEN_47; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_49 = io_mat1_5_4 != prevStationary_matrix_5_4 ? 1'h0 : _GEN_48; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_50 = io_mat1_5_5 != prevStationary_matrix_5_5 ? 1'h0 : _GEN_49; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_51 = io_mat1_5_6 != prevStationary_matrix_5_6 ? 1'h0 : _GEN_50; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_52 = io_mat1_5_7 != prevStationary_matrix_5_7 ? 1'h0 : _GEN_51; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_53 = io_mat2_5 != prevStreaming_matrix_5 ? 1'h0 : _GEN_52; // @[Muxes.scala 49:51 50:26]
  wire  _GEN_54 = io_mat1_6_0 != prevStationary_matrix_6_0 ? 1'h0 : _GEN_53; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_55 = io_mat1_6_1 != prevStationary_matrix_6_1 ? 1'h0 : _GEN_54; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_56 = io_mat1_6_2 != prevStationary_matrix_6_2 ? 1'h0 : _GEN_55; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_57 = io_mat1_6_3 != prevStationary_matrix_6_3 ? 1'h0 : _GEN_56; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_58 = io_mat1_6_4 != prevStationary_matrix_6_4 ? 1'h0 : _GEN_57; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_59 = io_mat1_6_5 != prevStationary_matrix_6_5 ? 1'h0 : _GEN_58; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_60 = io_mat1_6_6 != prevStationary_matrix_6_6 ? 1'h0 : _GEN_59; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_61 = io_mat1_6_7 != prevStationary_matrix_6_7 ? 1'h0 : _GEN_60; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_62 = io_mat2_6 != prevStreaming_matrix_6 ? 1'h0 : _GEN_61; // @[Muxes.scala 49:51 50:26]
  wire  _GEN_63 = io_mat1_7_0 != prevStationary_matrix_7_0 ? 1'h0 : _GEN_62; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_64 = io_mat1_7_1 != prevStationary_matrix_7_1 ? 1'h0 : _GEN_63; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_65 = io_mat1_7_2 != prevStationary_matrix_7_2 ? 1'h0 : _GEN_64; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_66 = io_mat1_7_3 != prevStationary_matrix_7_3 ? 1'h0 : _GEN_65; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_67 = io_mat1_7_4 != prevStationary_matrix_7_4 ? 1'h0 : _GEN_66; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_1676 = 3'h0 == j[2:0]; // @[Muxes.scala 54:{36,36}]
  wire  _GEN_1677 = 3'h1 == i[2:0]; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_73 = 3'h0 == j[2:0] & 3'h1 == i[2:0] ? io_counterMatrix1_0_1 : io_counterMatrix1_0_0; // @[Muxes.scala 54:{36,36}]
  wire  _GEN_1679 = 3'h2 == i[2:0]; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_74 = 3'h0 == j[2:0] & 3'h2 == i[2:0] ? io_counterMatrix1_0_2 : _GEN_73; // @[Muxes.scala 54:{36,36}]
  wire  _GEN_1681 = 3'h3 == i[2:0]; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_75 = 3'h0 == j[2:0] & 3'h3 == i[2:0] ? io_counterMatrix1_0_3 : _GEN_74; // @[Muxes.scala 54:{36,36}]
  wire  _GEN_1683 = 3'h4 == i[2:0]; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_76 = 3'h0 == j[2:0] & 3'h4 == i[2:0] ? io_counterMatrix1_0_4 : _GEN_75; // @[Muxes.scala 54:{36,36}]
  wire  _GEN_1685 = 3'h5 == i[2:0]; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_77 = 3'h0 == j[2:0] & 3'h5 == i[2:0] ? io_counterMatrix1_0_5 : _GEN_76; // @[Muxes.scala 54:{36,36}]
  wire  _GEN_1687 = 3'h6 == i[2:0]; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_78 = 3'h0 == j[2:0] & 3'h6 == i[2:0] ? io_counterMatrix1_0_6 : _GEN_77; // @[Muxes.scala 54:{36,36}]
  wire  _GEN_1689 = 3'h7 == i[2:0]; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_79 = 3'h0 == j[2:0] & 3'h7 == i[2:0] ? io_counterMatrix1_0_7 : _GEN_78; // @[Muxes.scala 54:{36,36}]
  wire  _GEN_1690 = 3'h1 == j[2:0]; // @[Muxes.scala 54:{36,36}]
  wire  _GEN_1691 = 3'h0 == i[2:0]; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_80 = 3'h1 == j[2:0] & 3'h0 == i[2:0] ? io_counterMatrix1_1_0 : _GEN_79; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_81 = 3'h1 == j[2:0] & 3'h1 == i[2:0] ? io_counterMatrix1_1_1 : _GEN_80; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_82 = 3'h1 == j[2:0] & 3'h2 == i[2:0] ? io_counterMatrix1_1_2 : _GEN_81; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_83 = 3'h1 == j[2:0] & 3'h3 == i[2:0] ? io_counterMatrix1_1_3 : _GEN_82; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_84 = 3'h1 == j[2:0] & 3'h4 == i[2:0] ? io_counterMatrix1_1_4 : _GEN_83; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_85 = 3'h1 == j[2:0] & 3'h5 == i[2:0] ? io_counterMatrix1_1_5 : _GEN_84; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_86 = 3'h1 == j[2:0] & 3'h6 == i[2:0] ? io_counterMatrix1_1_6 : _GEN_85; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_87 = 3'h1 == j[2:0] & 3'h7 == i[2:0] ? io_counterMatrix1_1_7 : _GEN_86; // @[Muxes.scala 54:{36,36}]
  wire  _GEN_1706 = 3'h2 == j[2:0]; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_88 = 3'h2 == j[2:0] & 3'h0 == i[2:0] ? io_counterMatrix1_2_0 : _GEN_87; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_89 = 3'h2 == j[2:0] & 3'h1 == i[2:0] ? io_counterMatrix1_2_1 : _GEN_88; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_90 = 3'h2 == j[2:0] & 3'h2 == i[2:0] ? io_counterMatrix1_2_2 : _GEN_89; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_91 = 3'h2 == j[2:0] & 3'h3 == i[2:0] ? io_counterMatrix1_2_3 : _GEN_90; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_92 = 3'h2 == j[2:0] & 3'h4 == i[2:0] ? io_counterMatrix1_2_4 : _GEN_91; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_93 = 3'h2 == j[2:0] & 3'h5 == i[2:0] ? io_counterMatrix1_2_5 : _GEN_92; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_94 = 3'h2 == j[2:0] & 3'h6 == i[2:0] ? io_counterMatrix1_2_6 : _GEN_93; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_95 = 3'h2 == j[2:0] & 3'h7 == i[2:0] ? io_counterMatrix1_2_7 : _GEN_94; // @[Muxes.scala 54:{36,36}]
  wire  _GEN_1722 = 3'h3 == j[2:0]; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_96 = 3'h3 == j[2:0] & 3'h0 == i[2:0] ? io_counterMatrix1_3_0 : _GEN_95; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_97 = 3'h3 == j[2:0] & 3'h1 == i[2:0] ? io_counterMatrix1_3_1 : _GEN_96; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_98 = 3'h3 == j[2:0] & 3'h2 == i[2:0] ? io_counterMatrix1_3_2 : _GEN_97; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_99 = 3'h3 == j[2:0] & 3'h3 == i[2:0] ? io_counterMatrix1_3_3 : _GEN_98; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_100 = 3'h3 == j[2:0] & 3'h4 == i[2:0] ? io_counterMatrix1_3_4 : _GEN_99; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_101 = 3'h3 == j[2:0] & 3'h5 == i[2:0] ? io_counterMatrix1_3_5 : _GEN_100; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_102 = 3'h3 == j[2:0] & 3'h6 == i[2:0] ? io_counterMatrix1_3_6 : _GEN_101; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_103 = 3'h3 == j[2:0] & 3'h7 == i[2:0] ? io_counterMatrix1_3_7 : _GEN_102; // @[Muxes.scala 54:{36,36}]
  wire  _GEN_1738 = 3'h4 == j[2:0]; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_104 = 3'h4 == j[2:0] & 3'h0 == i[2:0] ? io_counterMatrix1_4_0 : _GEN_103; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_105 = 3'h4 == j[2:0] & 3'h1 == i[2:0] ? io_counterMatrix1_4_1 : _GEN_104; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_106 = 3'h4 == j[2:0] & 3'h2 == i[2:0] ? io_counterMatrix1_4_2 : _GEN_105; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_107 = 3'h4 == j[2:0] & 3'h3 == i[2:0] ? io_counterMatrix1_4_3 : _GEN_106; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_108 = 3'h4 == j[2:0] & 3'h4 == i[2:0] ? io_counterMatrix1_4_4 : _GEN_107; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_109 = 3'h4 == j[2:0] & 3'h5 == i[2:0] ? io_counterMatrix1_4_5 : _GEN_108; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_110 = 3'h4 == j[2:0] & 3'h6 == i[2:0] ? io_counterMatrix1_4_6 : _GEN_109; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_111 = 3'h4 == j[2:0] & 3'h7 == i[2:0] ? io_counterMatrix1_4_7 : _GEN_110; // @[Muxes.scala 54:{36,36}]
  wire  _GEN_1754 = 3'h5 == j[2:0]; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_112 = 3'h5 == j[2:0] & 3'h0 == i[2:0] ? io_counterMatrix1_5_0 : _GEN_111; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_113 = 3'h5 == j[2:0] & 3'h1 == i[2:0] ? io_counterMatrix1_5_1 : _GEN_112; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_114 = 3'h5 == j[2:0] & 3'h2 == i[2:0] ? io_counterMatrix1_5_2 : _GEN_113; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_115 = 3'h5 == j[2:0] & 3'h3 == i[2:0] ? io_counterMatrix1_5_3 : _GEN_114; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_116 = 3'h5 == j[2:0] & 3'h4 == i[2:0] ? io_counterMatrix1_5_4 : _GEN_115; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_117 = 3'h5 == j[2:0] & 3'h5 == i[2:0] ? io_counterMatrix1_5_5 : _GEN_116; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_118 = 3'h5 == j[2:0] & 3'h6 == i[2:0] ? io_counterMatrix1_5_6 : _GEN_117; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_119 = 3'h5 == j[2:0] & 3'h7 == i[2:0] ? io_counterMatrix1_5_7 : _GEN_118; // @[Muxes.scala 54:{36,36}]
  wire  _GEN_1770 = 3'h6 == j[2:0]; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_120 = 3'h6 == j[2:0] & 3'h0 == i[2:0] ? io_counterMatrix1_6_0 : _GEN_119; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_121 = 3'h6 == j[2:0] & 3'h1 == i[2:0] ? io_counterMatrix1_6_1 : _GEN_120; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_122 = 3'h6 == j[2:0] & 3'h2 == i[2:0] ? io_counterMatrix1_6_2 : _GEN_121; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_123 = 3'h6 == j[2:0] & 3'h3 == i[2:0] ? io_counterMatrix1_6_3 : _GEN_122; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_124 = 3'h6 == j[2:0] & 3'h4 == i[2:0] ? io_counterMatrix1_6_4 : _GEN_123; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_125 = 3'h6 == j[2:0] & 3'h5 == i[2:0] ? io_counterMatrix1_6_5 : _GEN_124; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_126 = 3'h6 == j[2:0] & 3'h6 == i[2:0] ? io_counterMatrix1_6_6 : _GEN_125; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_127 = 3'h6 == j[2:0] & 3'h7 == i[2:0] ? io_counterMatrix1_6_7 : _GEN_126; // @[Muxes.scala 54:{36,36}]
  wire  _GEN_1786 = 3'h7 == j[2:0]; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_128 = 3'h7 == j[2:0] & 3'h0 == i[2:0] ? io_counterMatrix1_7_0 : _GEN_127; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_129 = 3'h7 == j[2:0] & 3'h1 == i[2:0] ? io_counterMatrix1_7_1 : _GEN_128; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_130 = 3'h7 == j[2:0] & 3'h2 == i[2:0] ? io_counterMatrix1_7_2 : _GEN_129; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_131 = 3'h7 == j[2:0] & 3'h3 == i[2:0] ? io_counterMatrix1_7_3 : _GEN_130; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_132 = 3'h7 == j[2:0] & 3'h4 == i[2:0] ? io_counterMatrix1_7_4 : _GEN_131; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_133 = 3'h7 == j[2:0] & 3'h5 == i[2:0] ? io_counterMatrix1_7_5 : _GEN_132; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_134 = 3'h7 == j[2:0] & 3'h6 == i[2:0] ? io_counterMatrix1_7_6 : _GEN_133; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_135 = 3'h7 == j[2:0] & 3'h7 == i[2:0] ? io_counterMatrix1_7_7 : _GEN_134; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_137 = 3'h1 == i[2:0] ? io_mat2_1 : io_mat2_0; // @[Muxes.scala 54:{60,60}]
  wire [15:0] _GEN_138 = 3'h2 == i[2:0] ? io_mat2_2 : _GEN_137; // @[Muxes.scala 54:{60,60}]
  wire [15:0] _GEN_139 = 3'h3 == i[2:0] ? io_mat2_3 : _GEN_138; // @[Muxes.scala 54:{60,60}]
  wire [15:0] _GEN_140 = 3'h4 == i[2:0] ? io_mat2_4 : _GEN_139; // @[Muxes.scala 54:{60,60}]
  wire [15:0] _GEN_141 = 3'h5 == i[2:0] ? io_mat2_5 : _GEN_140; // @[Muxes.scala 54:{60,60}]
  wire [15:0] _GEN_142 = 3'h6 == i[2:0] ? io_mat2_6 : _GEN_141; // @[Muxes.scala 54:{60,60}]
  wire [15:0] _GEN_143 = 3'h7 == i[2:0] ? io_mat2_7 : _GEN_142; // @[Muxes.scala 54:{60,60}]
  wire [15:0] _GEN_209 = 3'h1 == i[2:0] ? io_counterMatrix2_1 : io_counterMatrix2_0; // @[Muxes.scala 56:{38,38}]
  wire [15:0] _GEN_210 = 3'h2 == i[2:0] ? io_counterMatrix2_2 : _GEN_209; // @[Muxes.scala 56:{38,38}]
  wire [15:0] _GEN_211 = 3'h3 == i[2:0] ? io_counterMatrix2_3 : _GEN_210; // @[Muxes.scala 56:{38,38}]
  wire [15:0] _GEN_212 = 3'h4 == i[2:0] ? io_counterMatrix2_4 : _GEN_211; // @[Muxes.scala 56:{38,38}]
  wire [15:0] _GEN_213 = 3'h5 == i[2:0] ? io_counterMatrix2_5 : _GEN_212; // @[Muxes.scala 56:{38,38}]
  wire [15:0] _GEN_214 = 3'h6 == i[2:0] ? io_counterMatrix2_6 : _GEN_213; // @[Muxes.scala 56:{38,38}]
  wire [15:0] _GEN_215 = 3'h7 == i[2:0] ? io_counterMatrix2_7 : _GEN_214; // @[Muxes.scala 56:{38,38}]
  wire [15:0] _mux_T_2 = _GEN_215 - 16'h1; // @[Muxes.scala 57:51]
  wire [15:0] _mux_T_6 = _GEN_135 - 16'h1; // @[Muxes.scala 57:85]
  wire [15:0] _mux_T_8 = _mux_T_2 - _mux_T_6; // @[Muxes.scala 57:58]
  wire [3:0] _GEN_288 = 6'h0 == counter[5:0] ? _mux_T_8[3:0] : mux_0; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_289 = 6'h1 == counter[5:0] ? _mux_T_8[3:0] : mux_1; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_290 = 6'h2 == counter[5:0] ? _mux_T_8[3:0] : mux_2; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_291 = 6'h3 == counter[5:0] ? _mux_T_8[3:0] : mux_3; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_292 = 6'h4 == counter[5:0] ? _mux_T_8[3:0] : mux_4; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_293 = 6'h5 == counter[5:0] ? _mux_T_8[3:0] : mux_5; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_294 = 6'h6 == counter[5:0] ? _mux_T_8[3:0] : mux_6; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_295 = 6'h7 == counter[5:0] ? _mux_T_8[3:0] : mux_7; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_296 = 6'h8 == counter[5:0] ? _mux_T_8[3:0] : mux_8; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_297 = 6'h9 == counter[5:0] ? _mux_T_8[3:0] : mux_9; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_298 = 6'ha == counter[5:0] ? _mux_T_8[3:0] : mux_10; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_299 = 6'hb == counter[5:0] ? _mux_T_8[3:0] : mux_11; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_300 = 6'hc == counter[5:0] ? _mux_T_8[3:0] : mux_12; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_301 = 6'hd == counter[5:0] ? _mux_T_8[3:0] : mux_13; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_302 = 6'he == counter[5:0] ? _mux_T_8[3:0] : mux_14; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_303 = 6'hf == counter[5:0] ? _mux_T_8[3:0] : mux_15; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_304 = 6'h10 == counter[5:0] ? _mux_T_8[3:0] : mux_16; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_305 = 6'h11 == counter[5:0] ? _mux_T_8[3:0] : mux_17; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_306 = 6'h12 == counter[5:0] ? _mux_T_8[3:0] : mux_18; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_307 = 6'h13 == counter[5:0] ? _mux_T_8[3:0] : mux_19; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_308 = 6'h14 == counter[5:0] ? _mux_T_8[3:0] : mux_20; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_309 = 6'h15 == counter[5:0] ? _mux_T_8[3:0] : mux_21; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_310 = 6'h16 == counter[5:0] ? _mux_T_8[3:0] : mux_22; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_311 = 6'h17 == counter[5:0] ? _mux_T_8[3:0] : mux_23; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_312 = 6'h18 == counter[5:0] ? _mux_T_8[3:0] : mux_24; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_313 = 6'h19 == counter[5:0] ? _mux_T_8[3:0] : mux_25; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_314 = 6'h1a == counter[5:0] ? _mux_T_8[3:0] : mux_26; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_315 = 6'h1b == counter[5:0] ? _mux_T_8[3:0] : mux_27; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_316 = 6'h1c == counter[5:0] ? _mux_T_8[3:0] : mux_28; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_317 = 6'h1d == counter[5:0] ? _mux_T_8[3:0] : mux_29; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_318 = 6'h1e == counter[5:0] ? _mux_T_8[3:0] : mux_30; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_319 = 6'h1f == counter[5:0] ? _mux_T_8[3:0] : mux_31; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_320 = 6'h20 == counter[5:0] ? _mux_T_8[3:0] : mux_32; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_321 = 6'h21 == counter[5:0] ? _mux_T_8[3:0] : mux_33; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_322 = 6'h22 == counter[5:0] ? _mux_T_8[3:0] : mux_34; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_323 = 6'h23 == counter[5:0] ? _mux_T_8[3:0] : mux_35; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_324 = 6'h24 == counter[5:0] ? _mux_T_8[3:0] : mux_36; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_325 = 6'h25 == counter[5:0] ? _mux_T_8[3:0] : mux_37; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_326 = 6'h26 == counter[5:0] ? _mux_T_8[3:0] : mux_38; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_327 = 6'h27 == counter[5:0] ? _mux_T_8[3:0] : mux_39; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_328 = 6'h28 == counter[5:0] ? _mux_T_8[3:0] : mux_40; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_329 = 6'h29 == counter[5:0] ? _mux_T_8[3:0] : mux_41; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_330 = 6'h2a == counter[5:0] ? _mux_T_8[3:0] : mux_42; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_331 = 6'h2b == counter[5:0] ? _mux_T_8[3:0] : mux_43; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_332 = 6'h2c == counter[5:0] ? _mux_T_8[3:0] : mux_44; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_333 = 6'h2d == counter[5:0] ? _mux_T_8[3:0] : mux_45; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_334 = 6'h2e == counter[5:0] ? _mux_T_8[3:0] : mux_46; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_335 = 6'h2f == counter[5:0] ? _mux_T_8[3:0] : mux_47; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_336 = 6'h30 == counter[5:0] ? _mux_T_8[3:0] : mux_48; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_337 = 6'h31 == counter[5:0] ? _mux_T_8[3:0] : mux_49; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_338 = 6'h32 == counter[5:0] ? _mux_T_8[3:0] : mux_50; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_339 = 6'h33 == counter[5:0] ? _mux_T_8[3:0] : mux_51; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_340 = 6'h34 == counter[5:0] ? _mux_T_8[3:0] : mux_52; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_341 = 6'h35 == counter[5:0] ? _mux_T_8[3:0] : mux_53; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_342 = 6'h36 == counter[5:0] ? _mux_T_8[3:0] : mux_54; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_343 = 6'h37 == counter[5:0] ? _mux_T_8[3:0] : mux_55; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_344 = 6'h38 == counter[5:0] ? _mux_T_8[3:0] : mux_56; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_345 = 6'h39 == counter[5:0] ? _mux_T_8[3:0] : mux_57; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_346 = 6'h3a == counter[5:0] ? _mux_T_8[3:0] : mux_58; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_347 = 6'h3b == counter[5:0] ? _mux_T_8[3:0] : mux_59; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_348 = 6'h3c == counter[5:0] ? _mux_T_8[3:0] : mux_60; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_349 = 6'h3d == counter[5:0] ? _mux_T_8[3:0] : mux_61; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_350 = 6'h3e == counter[5:0] ? _mux_T_8[3:0] : mux_62; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_351 = 6'h3f == counter[5:0] ? _mux_T_8[3:0] : mux_63; // @[Muxes.scala 32:22 57:{24,24}]
  wire [15:0] _GEN_352 = 6'h0 == counter[5:0] ? _GEN_143 : src_0; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_353 = 6'h1 == counter[5:0] ? _GEN_143 : src_1; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_354 = 6'h2 == counter[5:0] ? _GEN_143 : src_2; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_355 = 6'h3 == counter[5:0] ? _GEN_143 : src_3; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_356 = 6'h4 == counter[5:0] ? _GEN_143 : src_4; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_357 = 6'h5 == counter[5:0] ? _GEN_143 : src_5; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_358 = 6'h6 == counter[5:0] ? _GEN_143 : src_6; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_359 = 6'h7 == counter[5:0] ? _GEN_143 : src_7; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_360 = 6'h8 == counter[5:0] ? _GEN_143 : src_8; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_361 = 6'h9 == counter[5:0] ? _GEN_143 : src_9; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_362 = 6'ha == counter[5:0] ? _GEN_143 : src_10; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_363 = 6'hb == counter[5:0] ? _GEN_143 : src_11; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_364 = 6'hc == counter[5:0] ? _GEN_143 : src_12; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_365 = 6'hd == counter[5:0] ? _GEN_143 : src_13; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_366 = 6'he == counter[5:0] ? _GEN_143 : src_14; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_367 = 6'hf == counter[5:0] ? _GEN_143 : src_15; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_368 = 6'h10 == counter[5:0] ? _GEN_143 : src_16; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_369 = 6'h11 == counter[5:0] ? _GEN_143 : src_17; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_370 = 6'h12 == counter[5:0] ? _GEN_143 : src_18; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_371 = 6'h13 == counter[5:0] ? _GEN_143 : src_19; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_372 = 6'h14 == counter[5:0] ? _GEN_143 : src_20; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_373 = 6'h15 == counter[5:0] ? _GEN_143 : src_21; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_374 = 6'h16 == counter[5:0] ? _GEN_143 : src_22; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_375 = 6'h17 == counter[5:0] ? _GEN_143 : src_23; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_376 = 6'h18 == counter[5:0] ? _GEN_143 : src_24; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_377 = 6'h19 == counter[5:0] ? _GEN_143 : src_25; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_378 = 6'h1a == counter[5:0] ? _GEN_143 : src_26; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_379 = 6'h1b == counter[5:0] ? _GEN_143 : src_27; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_380 = 6'h1c == counter[5:0] ? _GEN_143 : src_28; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_381 = 6'h1d == counter[5:0] ? _GEN_143 : src_29; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_382 = 6'h1e == counter[5:0] ? _GEN_143 : src_30; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_383 = 6'h1f == counter[5:0] ? _GEN_143 : src_31; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_384 = 6'h20 == counter[5:0] ? _GEN_143 : src_32; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_385 = 6'h21 == counter[5:0] ? _GEN_143 : src_33; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_386 = 6'h22 == counter[5:0] ? _GEN_143 : src_34; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_387 = 6'h23 == counter[5:0] ? _GEN_143 : src_35; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_388 = 6'h24 == counter[5:0] ? _GEN_143 : src_36; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_389 = 6'h25 == counter[5:0] ? _GEN_143 : src_37; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_390 = 6'h26 == counter[5:0] ? _GEN_143 : src_38; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_391 = 6'h27 == counter[5:0] ? _GEN_143 : src_39; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_392 = 6'h28 == counter[5:0] ? _GEN_143 : src_40; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_393 = 6'h29 == counter[5:0] ? _GEN_143 : src_41; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_394 = 6'h2a == counter[5:0] ? _GEN_143 : src_42; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_395 = 6'h2b == counter[5:0] ? _GEN_143 : src_43; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_396 = 6'h2c == counter[5:0] ? _GEN_143 : src_44; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_397 = 6'h2d == counter[5:0] ? _GEN_143 : src_45; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_398 = 6'h2e == counter[5:0] ? _GEN_143 : src_46; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_399 = 6'h2f == counter[5:0] ? _GEN_143 : src_47; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_400 = 6'h30 == counter[5:0] ? _GEN_143 : src_48; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_401 = 6'h31 == counter[5:0] ? _GEN_143 : src_49; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_402 = 6'h32 == counter[5:0] ? _GEN_143 : src_50; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_403 = 6'h33 == counter[5:0] ? _GEN_143 : src_51; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_404 = 6'h34 == counter[5:0] ? _GEN_143 : src_52; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_405 = 6'h35 == counter[5:0] ? _GEN_143 : src_53; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_406 = 6'h36 == counter[5:0] ? _GEN_143 : src_54; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_407 = 6'h37 == counter[5:0] ? _GEN_143 : src_55; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_408 = 6'h38 == counter[5:0] ? _GEN_143 : src_56; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_409 = 6'h39 == counter[5:0] ? _GEN_143 : src_57; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_410 = 6'h3a == counter[5:0] ? _GEN_143 : src_58; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_411 = 6'h3b == counter[5:0] ? _GEN_143 : src_59; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_412 = 6'h3c == counter[5:0] ? _GEN_143 : src_60; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_413 = 6'h3d == counter[5:0] ? _GEN_143 : src_61; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_414 = 6'h3e == counter[5:0] ? _GEN_143 : src_62; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_415 = 6'h3f == counter[5:0] ? _GEN_143 : src_63; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_489 = _GEN_1676 & _GEN_1677 ? io_mat1_0_1 : io_mat1_0_0; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_490 = _GEN_1676 & _GEN_1679 ? io_mat1_0_2 : _GEN_489; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_491 = _GEN_1676 & _GEN_1681 ? io_mat1_0_3 : _GEN_490; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_492 = _GEN_1676 & _GEN_1683 ? io_mat1_0_4 : _GEN_491; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_493 = _GEN_1676 & _GEN_1685 ? io_mat1_0_5 : _GEN_492; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_494 = _GEN_1676 & _GEN_1687 ? io_mat1_0_6 : _GEN_493; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_495 = _GEN_1676 & _GEN_1689 ? io_mat1_0_7 : _GEN_494; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_496 = _GEN_1690 & _GEN_1691 ? io_mat1_1_0 : _GEN_495; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_497 = _GEN_1690 & _GEN_1677 ? io_mat1_1_1 : _GEN_496; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_498 = _GEN_1690 & _GEN_1679 ? io_mat1_1_2 : _GEN_497; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_499 = _GEN_1690 & _GEN_1681 ? io_mat1_1_3 : _GEN_498; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_500 = _GEN_1690 & _GEN_1683 ? io_mat1_1_4 : _GEN_499; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_501 = _GEN_1690 & _GEN_1685 ? io_mat1_1_5 : _GEN_500; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_502 = _GEN_1690 & _GEN_1687 ? io_mat1_1_6 : _GEN_501; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_503 = _GEN_1690 & _GEN_1689 ? io_mat1_1_7 : _GEN_502; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_504 = _GEN_1706 & _GEN_1691 ? io_mat1_2_0 : _GEN_503; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_505 = _GEN_1706 & _GEN_1677 ? io_mat1_2_1 : _GEN_504; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_506 = _GEN_1706 & _GEN_1679 ? io_mat1_2_2 : _GEN_505; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_507 = _GEN_1706 & _GEN_1681 ? io_mat1_2_3 : _GEN_506; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_508 = _GEN_1706 & _GEN_1683 ? io_mat1_2_4 : _GEN_507; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_509 = _GEN_1706 & _GEN_1685 ? io_mat1_2_5 : _GEN_508; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_510 = _GEN_1706 & _GEN_1687 ? io_mat1_2_6 : _GEN_509; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_511 = _GEN_1706 & _GEN_1689 ? io_mat1_2_7 : _GEN_510; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_512 = _GEN_1722 & _GEN_1691 ? io_mat1_3_0 : _GEN_511; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_513 = _GEN_1722 & _GEN_1677 ? io_mat1_3_1 : _GEN_512; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_514 = _GEN_1722 & _GEN_1679 ? io_mat1_3_2 : _GEN_513; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_515 = _GEN_1722 & _GEN_1681 ? io_mat1_3_3 : _GEN_514; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_516 = _GEN_1722 & _GEN_1683 ? io_mat1_3_4 : _GEN_515; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_517 = _GEN_1722 & _GEN_1685 ? io_mat1_3_5 : _GEN_516; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_518 = _GEN_1722 & _GEN_1687 ? io_mat1_3_6 : _GEN_517; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_519 = _GEN_1722 & _GEN_1689 ? io_mat1_3_7 : _GEN_518; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_520 = _GEN_1738 & _GEN_1691 ? io_mat1_4_0 : _GEN_519; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_521 = _GEN_1738 & _GEN_1677 ? io_mat1_4_1 : _GEN_520; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_522 = _GEN_1738 & _GEN_1679 ? io_mat1_4_2 : _GEN_521; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_523 = _GEN_1738 & _GEN_1681 ? io_mat1_4_3 : _GEN_522; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_524 = _GEN_1738 & _GEN_1683 ? io_mat1_4_4 : _GEN_523; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_525 = _GEN_1738 & _GEN_1685 ? io_mat1_4_5 : _GEN_524; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_526 = _GEN_1738 & _GEN_1687 ? io_mat1_4_6 : _GEN_525; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_527 = _GEN_1738 & _GEN_1689 ? io_mat1_4_7 : _GEN_526; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_528 = _GEN_1754 & _GEN_1691 ? io_mat1_5_0 : _GEN_527; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_529 = _GEN_1754 & _GEN_1677 ? io_mat1_5_1 : _GEN_528; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_530 = _GEN_1754 & _GEN_1679 ? io_mat1_5_2 : _GEN_529; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_531 = _GEN_1754 & _GEN_1681 ? io_mat1_5_3 : _GEN_530; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_532 = _GEN_1754 & _GEN_1683 ? io_mat1_5_4 : _GEN_531; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_533 = _GEN_1754 & _GEN_1685 ? io_mat1_5_5 : _GEN_532; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_534 = _GEN_1754 & _GEN_1687 ? io_mat1_5_6 : _GEN_533; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_535 = _GEN_1754 & _GEN_1689 ? io_mat1_5_7 : _GEN_534; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_536 = _GEN_1770 & _GEN_1691 ? io_mat1_6_0 : _GEN_535; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_537 = _GEN_1770 & _GEN_1677 ? io_mat1_6_1 : _GEN_536; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_538 = _GEN_1770 & _GEN_1679 ? io_mat1_6_2 : _GEN_537; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_539 = _GEN_1770 & _GEN_1681 ? io_mat1_6_3 : _GEN_538; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_540 = _GEN_1770 & _GEN_1683 ? io_mat1_6_4 : _GEN_539; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_541 = _GEN_1770 & _GEN_1685 ? io_mat1_6_5 : _GEN_540; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_542 = _GEN_1770 & _GEN_1687 ? io_mat1_6_6 : _GEN_541; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_543 = _GEN_1770 & _GEN_1689 ? io_mat1_6_7 : _GEN_542; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_544 = _GEN_1786 & _GEN_1691 ? io_mat1_7_0 : _GEN_543; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_545 = _GEN_1786 & _GEN_1677 ? io_mat1_7_1 : _GEN_544; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_546 = _GEN_1786 & _GEN_1679 ? io_mat1_7_2 : _GEN_545; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_547 = _GEN_1786 & _GEN_1681 ? io_mat1_7_3 : _GEN_546; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_548 = _GEN_1786 & _GEN_1683 ? io_mat1_7_4 : _GEN_547; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_549 = _GEN_1786 & _GEN_1685 ? io_mat1_7_5 : _GEN_548; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_550 = _GEN_1786 & _GEN_1687 ? io_mat1_7_6 : _GEN_549; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_551 = _GEN_1786 & _GEN_1689 ? io_mat1_7_7 : _GEN_550; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_424 = 6'h0 == counter[5:0] ? _GEN_551 : dest_0; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_425 = 6'h1 == counter[5:0] ? _GEN_551 : dest_1; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_426 = 6'h2 == counter[5:0] ? _GEN_551 : dest_2; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_427 = 6'h3 == counter[5:0] ? _GEN_551 : dest_3; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_428 = 6'h4 == counter[5:0] ? _GEN_551 : dest_4; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_429 = 6'h5 == counter[5:0] ? _GEN_551 : dest_5; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_430 = 6'h6 == counter[5:0] ? _GEN_551 : dest_6; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_431 = 6'h7 == counter[5:0] ? _GEN_551 : dest_7; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_432 = 6'h8 == counter[5:0] ? _GEN_551 : dest_8; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_433 = 6'h9 == counter[5:0] ? _GEN_551 : dest_9; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_434 = 6'ha == counter[5:0] ? _GEN_551 : dest_10; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_435 = 6'hb == counter[5:0] ? _GEN_551 : dest_11; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_436 = 6'hc == counter[5:0] ? _GEN_551 : dest_12; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_437 = 6'hd == counter[5:0] ? _GEN_551 : dest_13; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_438 = 6'he == counter[5:0] ? _GEN_551 : dest_14; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_439 = 6'hf == counter[5:0] ? _GEN_551 : dest_15; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_440 = 6'h10 == counter[5:0] ? _GEN_551 : dest_16; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_441 = 6'h11 == counter[5:0] ? _GEN_551 : dest_17; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_442 = 6'h12 == counter[5:0] ? _GEN_551 : dest_18; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_443 = 6'h13 == counter[5:0] ? _GEN_551 : dest_19; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_444 = 6'h14 == counter[5:0] ? _GEN_551 : dest_20; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_445 = 6'h15 == counter[5:0] ? _GEN_551 : dest_21; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_446 = 6'h16 == counter[5:0] ? _GEN_551 : dest_22; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_447 = 6'h17 == counter[5:0] ? _GEN_551 : dest_23; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_448 = 6'h18 == counter[5:0] ? _GEN_551 : dest_24; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_449 = 6'h19 == counter[5:0] ? _GEN_551 : dest_25; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_450 = 6'h1a == counter[5:0] ? _GEN_551 : dest_26; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_451 = 6'h1b == counter[5:0] ? _GEN_551 : dest_27; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_452 = 6'h1c == counter[5:0] ? _GEN_551 : dest_28; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_453 = 6'h1d == counter[5:0] ? _GEN_551 : dest_29; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_454 = 6'h1e == counter[5:0] ? _GEN_551 : dest_30; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_455 = 6'h1f == counter[5:0] ? _GEN_551 : dest_31; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_456 = 6'h20 == counter[5:0] ? _GEN_551 : dest_32; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_457 = 6'h21 == counter[5:0] ? _GEN_551 : dest_33; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_458 = 6'h22 == counter[5:0] ? _GEN_551 : dest_34; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_459 = 6'h23 == counter[5:0] ? _GEN_551 : dest_35; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_460 = 6'h24 == counter[5:0] ? _GEN_551 : dest_36; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_461 = 6'h25 == counter[5:0] ? _GEN_551 : dest_37; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_462 = 6'h26 == counter[5:0] ? _GEN_551 : dest_38; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_463 = 6'h27 == counter[5:0] ? _GEN_551 : dest_39; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_464 = 6'h28 == counter[5:0] ? _GEN_551 : dest_40; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_465 = 6'h29 == counter[5:0] ? _GEN_551 : dest_41; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_466 = 6'h2a == counter[5:0] ? _GEN_551 : dest_42; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_467 = 6'h2b == counter[5:0] ? _GEN_551 : dest_43; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_468 = 6'h2c == counter[5:0] ? _GEN_551 : dest_44; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_469 = 6'h2d == counter[5:0] ? _GEN_551 : dest_45; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_470 = 6'h2e == counter[5:0] ? _GEN_551 : dest_46; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_471 = 6'h2f == counter[5:0] ? _GEN_551 : dest_47; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_472 = 6'h30 == counter[5:0] ? _GEN_551 : dest_48; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_473 = 6'h31 == counter[5:0] ? _GEN_551 : dest_49; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_474 = 6'h32 == counter[5:0] ? _GEN_551 : dest_50; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_475 = 6'h33 == counter[5:0] ? _GEN_551 : dest_51; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_476 = 6'h34 == counter[5:0] ? _GEN_551 : dest_52; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_477 = 6'h35 == counter[5:0] ? _GEN_551 : dest_53; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_478 = 6'h36 == counter[5:0] ? _GEN_551 : dest_54; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_479 = 6'h37 == counter[5:0] ? _GEN_551 : dest_55; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_480 = 6'h38 == counter[5:0] ? _GEN_551 : dest_56; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_481 = 6'h39 == counter[5:0] ? _GEN_551 : dest_57; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_482 = 6'h3a == counter[5:0] ? _GEN_551 : dest_58; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_483 = 6'h3b == counter[5:0] ? _GEN_551 : dest_59; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_484 = 6'h3c == counter[5:0] ? _GEN_551 : dest_60; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_485 = 6'h3d == counter[5:0] ? _GEN_551 : dest_61; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_486 = 6'h3e == counter[5:0] ? _GEN_551 : dest_62; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_487 = 6'h3f == counter[5:0] ? _GEN_551 : dest_63; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _mux_T_17 = _mux_T_6 - _mux_T_2; // @[Muxes.scala 61:61]
  wire [3:0] _GEN_624 = 6'h0 == counter[5:0] ? _mux_T_17[3:0] : mux_0; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_625 = 6'h1 == counter[5:0] ? _mux_T_17[3:0] : mux_1; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_626 = 6'h2 == counter[5:0] ? _mux_T_17[3:0] : mux_2; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_627 = 6'h3 == counter[5:0] ? _mux_T_17[3:0] : mux_3; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_628 = 6'h4 == counter[5:0] ? _mux_T_17[3:0] : mux_4; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_629 = 6'h5 == counter[5:0] ? _mux_T_17[3:0] : mux_5; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_630 = 6'h6 == counter[5:0] ? _mux_T_17[3:0] : mux_6; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_631 = 6'h7 == counter[5:0] ? _mux_T_17[3:0] : mux_7; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_632 = 6'h8 == counter[5:0] ? _mux_T_17[3:0] : mux_8; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_633 = 6'h9 == counter[5:0] ? _mux_T_17[3:0] : mux_9; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_634 = 6'ha == counter[5:0] ? _mux_T_17[3:0] : mux_10; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_635 = 6'hb == counter[5:0] ? _mux_T_17[3:0] : mux_11; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_636 = 6'hc == counter[5:0] ? _mux_T_17[3:0] : mux_12; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_637 = 6'hd == counter[5:0] ? _mux_T_17[3:0] : mux_13; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_638 = 6'he == counter[5:0] ? _mux_T_17[3:0] : mux_14; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_639 = 6'hf == counter[5:0] ? _mux_T_17[3:0] : mux_15; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_640 = 6'h10 == counter[5:0] ? _mux_T_17[3:0] : mux_16; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_641 = 6'h11 == counter[5:0] ? _mux_T_17[3:0] : mux_17; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_642 = 6'h12 == counter[5:0] ? _mux_T_17[3:0] : mux_18; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_643 = 6'h13 == counter[5:0] ? _mux_T_17[3:0] : mux_19; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_644 = 6'h14 == counter[5:0] ? _mux_T_17[3:0] : mux_20; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_645 = 6'h15 == counter[5:0] ? _mux_T_17[3:0] : mux_21; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_646 = 6'h16 == counter[5:0] ? _mux_T_17[3:0] : mux_22; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_647 = 6'h17 == counter[5:0] ? _mux_T_17[3:0] : mux_23; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_648 = 6'h18 == counter[5:0] ? _mux_T_17[3:0] : mux_24; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_649 = 6'h19 == counter[5:0] ? _mux_T_17[3:0] : mux_25; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_650 = 6'h1a == counter[5:0] ? _mux_T_17[3:0] : mux_26; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_651 = 6'h1b == counter[5:0] ? _mux_T_17[3:0] : mux_27; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_652 = 6'h1c == counter[5:0] ? _mux_T_17[3:0] : mux_28; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_653 = 6'h1d == counter[5:0] ? _mux_T_17[3:0] : mux_29; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_654 = 6'h1e == counter[5:0] ? _mux_T_17[3:0] : mux_30; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_655 = 6'h1f == counter[5:0] ? _mux_T_17[3:0] : mux_31; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_656 = 6'h20 == counter[5:0] ? _mux_T_17[3:0] : mux_32; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_657 = 6'h21 == counter[5:0] ? _mux_T_17[3:0] : mux_33; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_658 = 6'h22 == counter[5:0] ? _mux_T_17[3:0] : mux_34; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_659 = 6'h23 == counter[5:0] ? _mux_T_17[3:0] : mux_35; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_660 = 6'h24 == counter[5:0] ? _mux_T_17[3:0] : mux_36; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_661 = 6'h25 == counter[5:0] ? _mux_T_17[3:0] : mux_37; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_662 = 6'h26 == counter[5:0] ? _mux_T_17[3:0] : mux_38; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_663 = 6'h27 == counter[5:0] ? _mux_T_17[3:0] : mux_39; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_664 = 6'h28 == counter[5:0] ? _mux_T_17[3:0] : mux_40; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_665 = 6'h29 == counter[5:0] ? _mux_T_17[3:0] : mux_41; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_666 = 6'h2a == counter[5:0] ? _mux_T_17[3:0] : mux_42; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_667 = 6'h2b == counter[5:0] ? _mux_T_17[3:0] : mux_43; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_668 = 6'h2c == counter[5:0] ? _mux_T_17[3:0] : mux_44; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_669 = 6'h2d == counter[5:0] ? _mux_T_17[3:0] : mux_45; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_670 = 6'h2e == counter[5:0] ? _mux_T_17[3:0] : mux_46; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_671 = 6'h2f == counter[5:0] ? _mux_T_17[3:0] : mux_47; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_672 = 6'h30 == counter[5:0] ? _mux_T_17[3:0] : mux_48; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_673 = 6'h31 == counter[5:0] ? _mux_T_17[3:0] : mux_49; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_674 = 6'h32 == counter[5:0] ? _mux_T_17[3:0] : mux_50; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_675 = 6'h33 == counter[5:0] ? _mux_T_17[3:0] : mux_51; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_676 = 6'h34 == counter[5:0] ? _mux_T_17[3:0] : mux_52; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_677 = 6'h35 == counter[5:0] ? _mux_T_17[3:0] : mux_53; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_678 = 6'h36 == counter[5:0] ? _mux_T_17[3:0] : mux_54; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_679 = 6'h37 == counter[5:0] ? _mux_T_17[3:0] : mux_55; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_680 = 6'h38 == counter[5:0] ? _mux_T_17[3:0] : mux_56; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_681 = 6'h39 == counter[5:0] ? _mux_T_17[3:0] : mux_57; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_682 = 6'h3a == counter[5:0] ? _mux_T_17[3:0] : mux_58; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_683 = 6'h3b == counter[5:0] ? _mux_T_17[3:0] : mux_59; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_684 = 6'h3c == counter[5:0] ? _mux_T_17[3:0] : mux_60; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_685 = 6'h3d == counter[5:0] ? _mux_T_17[3:0] : mux_61; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_686 = 6'h3e == counter[5:0] ? _mux_T_17[3:0] : mux_62; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_687 = 6'h3f == counter[5:0] ? _mux_T_17[3:0] : mux_63; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_888 = _GEN_135 <= _GEN_215 ? _GEN_288 : _GEN_624; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_889 = _GEN_135 <= _GEN_215 ? _GEN_289 : _GEN_625; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_890 = _GEN_135 <= _GEN_215 ? _GEN_290 : _GEN_626; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_891 = _GEN_135 <= _GEN_215 ? _GEN_291 : _GEN_627; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_892 = _GEN_135 <= _GEN_215 ? _GEN_292 : _GEN_628; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_893 = _GEN_135 <= _GEN_215 ? _GEN_293 : _GEN_629; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_894 = _GEN_135 <= _GEN_215 ? _GEN_294 : _GEN_630; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_895 = _GEN_135 <= _GEN_215 ? _GEN_295 : _GEN_631; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_896 = _GEN_135 <= _GEN_215 ? _GEN_296 : _GEN_632; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_897 = _GEN_135 <= _GEN_215 ? _GEN_297 : _GEN_633; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_898 = _GEN_135 <= _GEN_215 ? _GEN_298 : _GEN_634; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_899 = _GEN_135 <= _GEN_215 ? _GEN_299 : _GEN_635; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_900 = _GEN_135 <= _GEN_215 ? _GEN_300 : _GEN_636; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_901 = _GEN_135 <= _GEN_215 ? _GEN_301 : _GEN_637; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_902 = _GEN_135 <= _GEN_215 ? _GEN_302 : _GEN_638; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_903 = _GEN_135 <= _GEN_215 ? _GEN_303 : _GEN_639; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_904 = _GEN_135 <= _GEN_215 ? _GEN_304 : _GEN_640; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_905 = _GEN_135 <= _GEN_215 ? _GEN_305 : _GEN_641; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_906 = _GEN_135 <= _GEN_215 ? _GEN_306 : _GEN_642; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_907 = _GEN_135 <= _GEN_215 ? _GEN_307 : _GEN_643; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_908 = _GEN_135 <= _GEN_215 ? _GEN_308 : _GEN_644; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_909 = _GEN_135 <= _GEN_215 ? _GEN_309 : _GEN_645; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_910 = _GEN_135 <= _GEN_215 ? _GEN_310 : _GEN_646; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_911 = _GEN_135 <= _GEN_215 ? _GEN_311 : _GEN_647; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_912 = _GEN_135 <= _GEN_215 ? _GEN_312 : _GEN_648; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_913 = _GEN_135 <= _GEN_215 ? _GEN_313 : _GEN_649; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_914 = _GEN_135 <= _GEN_215 ? _GEN_314 : _GEN_650; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_915 = _GEN_135 <= _GEN_215 ? _GEN_315 : _GEN_651; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_916 = _GEN_135 <= _GEN_215 ? _GEN_316 : _GEN_652; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_917 = _GEN_135 <= _GEN_215 ? _GEN_317 : _GEN_653; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_918 = _GEN_135 <= _GEN_215 ? _GEN_318 : _GEN_654; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_919 = _GEN_135 <= _GEN_215 ? _GEN_319 : _GEN_655; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_920 = _GEN_135 <= _GEN_215 ? _GEN_320 : _GEN_656; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_921 = _GEN_135 <= _GEN_215 ? _GEN_321 : _GEN_657; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_922 = _GEN_135 <= _GEN_215 ? _GEN_322 : _GEN_658; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_923 = _GEN_135 <= _GEN_215 ? _GEN_323 : _GEN_659; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_924 = _GEN_135 <= _GEN_215 ? _GEN_324 : _GEN_660; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_925 = _GEN_135 <= _GEN_215 ? _GEN_325 : _GEN_661; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_926 = _GEN_135 <= _GEN_215 ? _GEN_326 : _GEN_662; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_927 = _GEN_135 <= _GEN_215 ? _GEN_327 : _GEN_663; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_928 = _GEN_135 <= _GEN_215 ? _GEN_328 : _GEN_664; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_929 = _GEN_135 <= _GEN_215 ? _GEN_329 : _GEN_665; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_930 = _GEN_135 <= _GEN_215 ? _GEN_330 : _GEN_666; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_931 = _GEN_135 <= _GEN_215 ? _GEN_331 : _GEN_667; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_932 = _GEN_135 <= _GEN_215 ? _GEN_332 : _GEN_668; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_933 = _GEN_135 <= _GEN_215 ? _GEN_333 : _GEN_669; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_934 = _GEN_135 <= _GEN_215 ? _GEN_334 : _GEN_670; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_935 = _GEN_135 <= _GEN_215 ? _GEN_335 : _GEN_671; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_936 = _GEN_135 <= _GEN_215 ? _GEN_336 : _GEN_672; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_937 = _GEN_135 <= _GEN_215 ? _GEN_337 : _GEN_673; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_938 = _GEN_135 <= _GEN_215 ? _GEN_338 : _GEN_674; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_939 = _GEN_135 <= _GEN_215 ? _GEN_339 : _GEN_675; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_940 = _GEN_135 <= _GEN_215 ? _GEN_340 : _GEN_676; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_941 = _GEN_135 <= _GEN_215 ? _GEN_341 : _GEN_677; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_942 = _GEN_135 <= _GEN_215 ? _GEN_342 : _GEN_678; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_943 = _GEN_135 <= _GEN_215 ? _GEN_343 : _GEN_679; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_944 = _GEN_135 <= _GEN_215 ? _GEN_344 : _GEN_680; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_945 = _GEN_135 <= _GEN_215 ? _GEN_345 : _GEN_681; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_946 = _GEN_135 <= _GEN_215 ? _GEN_346 : _GEN_682; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_947 = _GEN_135 <= _GEN_215 ? _GEN_347 : _GEN_683; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_948 = _GEN_135 <= _GEN_215 ? _GEN_348 : _GEN_684; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_949 = _GEN_135 <= _GEN_215 ? _GEN_349 : _GEN_685; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_950 = _GEN_135 <= _GEN_215 ? _GEN_350 : _GEN_686; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_951 = _GEN_135 <= _GEN_215 ? _GEN_351 : _GEN_687; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_952 = _GEN_135 <= _GEN_215 ? _GEN_352 : _GEN_352; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_953 = _GEN_135 <= _GEN_215 ? _GEN_353 : _GEN_353; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_954 = _GEN_135 <= _GEN_215 ? _GEN_354 : _GEN_354; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_955 = _GEN_135 <= _GEN_215 ? _GEN_355 : _GEN_355; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_956 = _GEN_135 <= _GEN_215 ? _GEN_356 : _GEN_356; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_957 = _GEN_135 <= _GEN_215 ? _GEN_357 : _GEN_357; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_958 = _GEN_135 <= _GEN_215 ? _GEN_358 : _GEN_358; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_959 = _GEN_135 <= _GEN_215 ? _GEN_359 : _GEN_359; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_960 = _GEN_135 <= _GEN_215 ? _GEN_360 : _GEN_360; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_961 = _GEN_135 <= _GEN_215 ? _GEN_361 : _GEN_361; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_962 = _GEN_135 <= _GEN_215 ? _GEN_362 : _GEN_362; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_963 = _GEN_135 <= _GEN_215 ? _GEN_363 : _GEN_363; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_964 = _GEN_135 <= _GEN_215 ? _GEN_364 : _GEN_364; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_965 = _GEN_135 <= _GEN_215 ? _GEN_365 : _GEN_365; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_966 = _GEN_135 <= _GEN_215 ? _GEN_366 : _GEN_366; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_967 = _GEN_135 <= _GEN_215 ? _GEN_367 : _GEN_367; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_968 = _GEN_135 <= _GEN_215 ? _GEN_368 : _GEN_368; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_969 = _GEN_135 <= _GEN_215 ? _GEN_369 : _GEN_369; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_970 = _GEN_135 <= _GEN_215 ? _GEN_370 : _GEN_370; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_971 = _GEN_135 <= _GEN_215 ? _GEN_371 : _GEN_371; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_972 = _GEN_135 <= _GEN_215 ? _GEN_372 : _GEN_372; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_973 = _GEN_135 <= _GEN_215 ? _GEN_373 : _GEN_373; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_974 = _GEN_135 <= _GEN_215 ? _GEN_374 : _GEN_374; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_975 = _GEN_135 <= _GEN_215 ? _GEN_375 : _GEN_375; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_976 = _GEN_135 <= _GEN_215 ? _GEN_376 : _GEN_376; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_977 = _GEN_135 <= _GEN_215 ? _GEN_377 : _GEN_377; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_978 = _GEN_135 <= _GEN_215 ? _GEN_378 : _GEN_378; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_979 = _GEN_135 <= _GEN_215 ? _GEN_379 : _GEN_379; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_980 = _GEN_135 <= _GEN_215 ? _GEN_380 : _GEN_380; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_981 = _GEN_135 <= _GEN_215 ? _GEN_381 : _GEN_381; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_982 = _GEN_135 <= _GEN_215 ? _GEN_382 : _GEN_382; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_983 = _GEN_135 <= _GEN_215 ? _GEN_383 : _GEN_383; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_984 = _GEN_135 <= _GEN_215 ? _GEN_384 : _GEN_384; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_985 = _GEN_135 <= _GEN_215 ? _GEN_385 : _GEN_385; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_986 = _GEN_135 <= _GEN_215 ? _GEN_386 : _GEN_386; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_987 = _GEN_135 <= _GEN_215 ? _GEN_387 : _GEN_387; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_988 = _GEN_135 <= _GEN_215 ? _GEN_388 : _GEN_388; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_989 = _GEN_135 <= _GEN_215 ? _GEN_389 : _GEN_389; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_990 = _GEN_135 <= _GEN_215 ? _GEN_390 : _GEN_390; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_991 = _GEN_135 <= _GEN_215 ? _GEN_391 : _GEN_391; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_992 = _GEN_135 <= _GEN_215 ? _GEN_392 : _GEN_392; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_993 = _GEN_135 <= _GEN_215 ? _GEN_393 : _GEN_393; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_994 = _GEN_135 <= _GEN_215 ? _GEN_394 : _GEN_394; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_995 = _GEN_135 <= _GEN_215 ? _GEN_395 : _GEN_395; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_996 = _GEN_135 <= _GEN_215 ? _GEN_396 : _GEN_396; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_997 = _GEN_135 <= _GEN_215 ? _GEN_397 : _GEN_397; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_998 = _GEN_135 <= _GEN_215 ? _GEN_398 : _GEN_398; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_999 = _GEN_135 <= _GEN_215 ? _GEN_399 : _GEN_399; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1000 = _GEN_135 <= _GEN_215 ? _GEN_400 : _GEN_400; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1001 = _GEN_135 <= _GEN_215 ? _GEN_401 : _GEN_401; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1002 = _GEN_135 <= _GEN_215 ? _GEN_402 : _GEN_402; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1003 = _GEN_135 <= _GEN_215 ? _GEN_403 : _GEN_403; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1004 = _GEN_135 <= _GEN_215 ? _GEN_404 : _GEN_404; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1005 = _GEN_135 <= _GEN_215 ? _GEN_405 : _GEN_405; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1006 = _GEN_135 <= _GEN_215 ? _GEN_406 : _GEN_406; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1007 = _GEN_135 <= _GEN_215 ? _GEN_407 : _GEN_407; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1008 = _GEN_135 <= _GEN_215 ? _GEN_408 : _GEN_408; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1009 = _GEN_135 <= _GEN_215 ? _GEN_409 : _GEN_409; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1010 = _GEN_135 <= _GEN_215 ? _GEN_410 : _GEN_410; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1011 = _GEN_135 <= _GEN_215 ? _GEN_411 : _GEN_411; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1012 = _GEN_135 <= _GEN_215 ? _GEN_412 : _GEN_412; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1013 = _GEN_135 <= _GEN_215 ? _GEN_413 : _GEN_413; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1014 = _GEN_135 <= _GEN_215 ? _GEN_414 : _GEN_414; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1015 = _GEN_135 <= _GEN_215 ? _GEN_415 : _GEN_415; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1016 = _GEN_135 <= _GEN_215 ? _GEN_424 : _GEN_424; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1017 = _GEN_135 <= _GEN_215 ? _GEN_425 : _GEN_425; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1018 = _GEN_135 <= _GEN_215 ? _GEN_426 : _GEN_426; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1019 = _GEN_135 <= _GEN_215 ? _GEN_427 : _GEN_427; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1020 = _GEN_135 <= _GEN_215 ? _GEN_428 : _GEN_428; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1021 = _GEN_135 <= _GEN_215 ? _GEN_429 : _GEN_429; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1022 = _GEN_135 <= _GEN_215 ? _GEN_430 : _GEN_430; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1023 = _GEN_135 <= _GEN_215 ? _GEN_431 : _GEN_431; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1024 = _GEN_135 <= _GEN_215 ? _GEN_432 : _GEN_432; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1025 = _GEN_135 <= _GEN_215 ? _GEN_433 : _GEN_433; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1026 = _GEN_135 <= _GEN_215 ? _GEN_434 : _GEN_434; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1027 = _GEN_135 <= _GEN_215 ? _GEN_435 : _GEN_435; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1028 = _GEN_135 <= _GEN_215 ? _GEN_436 : _GEN_436; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1029 = _GEN_135 <= _GEN_215 ? _GEN_437 : _GEN_437; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1030 = _GEN_135 <= _GEN_215 ? _GEN_438 : _GEN_438; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1031 = _GEN_135 <= _GEN_215 ? _GEN_439 : _GEN_439; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1032 = _GEN_135 <= _GEN_215 ? _GEN_440 : _GEN_440; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1033 = _GEN_135 <= _GEN_215 ? _GEN_441 : _GEN_441; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1034 = _GEN_135 <= _GEN_215 ? _GEN_442 : _GEN_442; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1035 = _GEN_135 <= _GEN_215 ? _GEN_443 : _GEN_443; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1036 = _GEN_135 <= _GEN_215 ? _GEN_444 : _GEN_444; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1037 = _GEN_135 <= _GEN_215 ? _GEN_445 : _GEN_445; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1038 = _GEN_135 <= _GEN_215 ? _GEN_446 : _GEN_446; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1039 = _GEN_135 <= _GEN_215 ? _GEN_447 : _GEN_447; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1040 = _GEN_135 <= _GEN_215 ? _GEN_448 : _GEN_448; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1041 = _GEN_135 <= _GEN_215 ? _GEN_449 : _GEN_449; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1042 = _GEN_135 <= _GEN_215 ? _GEN_450 : _GEN_450; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1043 = _GEN_135 <= _GEN_215 ? _GEN_451 : _GEN_451; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1044 = _GEN_135 <= _GEN_215 ? _GEN_452 : _GEN_452; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1045 = _GEN_135 <= _GEN_215 ? _GEN_453 : _GEN_453; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1046 = _GEN_135 <= _GEN_215 ? _GEN_454 : _GEN_454; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1047 = _GEN_135 <= _GEN_215 ? _GEN_455 : _GEN_455; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1048 = _GEN_135 <= _GEN_215 ? _GEN_456 : _GEN_456; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1049 = _GEN_135 <= _GEN_215 ? _GEN_457 : _GEN_457; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1050 = _GEN_135 <= _GEN_215 ? _GEN_458 : _GEN_458; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1051 = _GEN_135 <= _GEN_215 ? _GEN_459 : _GEN_459; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1052 = _GEN_135 <= _GEN_215 ? _GEN_460 : _GEN_460; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1053 = _GEN_135 <= _GEN_215 ? _GEN_461 : _GEN_461; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1054 = _GEN_135 <= _GEN_215 ? _GEN_462 : _GEN_462; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1055 = _GEN_135 <= _GEN_215 ? _GEN_463 : _GEN_463; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1056 = _GEN_135 <= _GEN_215 ? _GEN_464 : _GEN_464; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1057 = _GEN_135 <= _GEN_215 ? _GEN_465 : _GEN_465; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1058 = _GEN_135 <= _GEN_215 ? _GEN_466 : _GEN_466; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1059 = _GEN_135 <= _GEN_215 ? _GEN_467 : _GEN_467; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1060 = _GEN_135 <= _GEN_215 ? _GEN_468 : _GEN_468; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1061 = _GEN_135 <= _GEN_215 ? _GEN_469 : _GEN_469; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1062 = _GEN_135 <= _GEN_215 ? _GEN_470 : _GEN_470; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1063 = _GEN_135 <= _GEN_215 ? _GEN_471 : _GEN_471; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1064 = _GEN_135 <= _GEN_215 ? _GEN_472 : _GEN_472; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1065 = _GEN_135 <= _GEN_215 ? _GEN_473 : _GEN_473; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1066 = _GEN_135 <= _GEN_215 ? _GEN_474 : _GEN_474; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1067 = _GEN_135 <= _GEN_215 ? _GEN_475 : _GEN_475; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1068 = _GEN_135 <= _GEN_215 ? _GEN_476 : _GEN_476; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1069 = _GEN_135 <= _GEN_215 ? _GEN_477 : _GEN_477; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1070 = _GEN_135 <= _GEN_215 ? _GEN_478 : _GEN_478; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1071 = _GEN_135 <= _GEN_215 ? _GEN_479 : _GEN_479; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1072 = _GEN_135 <= _GEN_215 ? _GEN_480 : _GEN_480; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1073 = _GEN_135 <= _GEN_215 ? _GEN_481 : _GEN_481; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1074 = _GEN_135 <= _GEN_215 ? _GEN_482 : _GEN_482; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1075 = _GEN_135 <= _GEN_215 ? _GEN_483 : _GEN_483; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1076 = _GEN_135 <= _GEN_215 ? _GEN_484 : _GEN_484; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1077 = _GEN_135 <= _GEN_215 ? _GEN_485 : _GEN_485; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1078 = _GEN_135 <= _GEN_215 ? _GEN_486 : _GEN_486; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_1079 = _GEN_135 <= _GEN_215 ? _GEN_487 : _GEN_487; // @[Muxes.scala 56:62]
  wire  _T_88 = ~jValid; // @[Muxes.scala 66:15]
  wire  _T_89 = j == 32'h7; // @[Muxes.scala 68:22]
  wire  _T_90 = i == 32'h7; // @[Muxes.scala 68:56]
  wire  _T_91 = j == 32'h7 & i == 32'h7; // @[Muxes.scala 68:50]
  wire [31:0] _counter_T_1 = counter + 32'h1; // @[Muxes.scala 69:30]
  wire [31:0] _GEN_1080 = ~(j == 32'h7 & i == 32'h7) ? _counter_T_1 : counter; // @[Muxes.scala 68:85 69:19 31:26]
  wire [31:0] _GEN_1081 = ~jValid ? _GEN_1080 : counter; // @[Muxes.scala 66:24 31:26]
  wire [3:0] _GEN_1082 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_888 : mux_0; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1083 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_889 : mux_1; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1084 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_890 : mux_2; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1085 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_891 : mux_3; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1086 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_892 : mux_4; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1087 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_893 : mux_5; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1088 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_894 : mux_6; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1089 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_895 : mux_7; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1090 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_896 : mux_8; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1091 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_897 : mux_9; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1092 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_898 : mux_10; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1093 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_899 : mux_11; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1094 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_900 : mux_12; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1095 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_901 : mux_13; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1096 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_902 : mux_14; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1097 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_903 : mux_15; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1098 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_904 : mux_16; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1099 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_905 : mux_17; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1100 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_906 : mux_18; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1101 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_907 : mux_19; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1102 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_908 : mux_20; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1103 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_909 : mux_21; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1104 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_910 : mux_22; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1105 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_911 : mux_23; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1106 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_912 : mux_24; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1107 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_913 : mux_25; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1108 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_914 : mux_26; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1109 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_915 : mux_27; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1110 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_916 : mux_28; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1111 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_917 : mux_29; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1112 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_918 : mux_30; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1113 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_919 : mux_31; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1114 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_920 : mux_32; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1115 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_921 : mux_33; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1116 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_922 : mux_34; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1117 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_923 : mux_35; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1118 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_924 : mux_36; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1119 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_925 : mux_37; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1120 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_926 : mux_38; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1121 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_927 : mux_39; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1122 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_928 : mux_40; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1123 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_929 : mux_41; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1124 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_930 : mux_42; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1125 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_931 : mux_43; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1126 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_932 : mux_44; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1127 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_933 : mux_45; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1128 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_934 : mux_46; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1129 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_935 : mux_47; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1130 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_936 : mux_48; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1131 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_937 : mux_49; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1132 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_938 : mux_50; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1133 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_939 : mux_51; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1134 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_940 : mux_52; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1135 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_941 : mux_53; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1136 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_942 : mux_54; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1137 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_943 : mux_55; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1138 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_944 : mux_56; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1139 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_945 : mux_57; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1140 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_946 : mux_58; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1141 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_947 : mux_59; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1142 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_948 : mux_60; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1143 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_949 : mux_61; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1144 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_950 : mux_62; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_1145 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_951 : mux_63; // @[Muxes.scala 32:22 54:70]
  wire [15:0] _GEN_1146 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_952 : src_0; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1147 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_953 : src_1; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1148 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_954 : src_2; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1149 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_955 : src_3; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1150 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_956 : src_4; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1151 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_957 : src_5; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1152 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_958 : src_6; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1153 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_959 : src_7; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1154 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_960 : src_8; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1155 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_961 : src_9; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1156 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_962 : src_10; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1157 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_963 : src_11; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1158 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_964 : src_12; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1159 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_965 : src_13; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1160 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_966 : src_14; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1161 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_967 : src_15; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1162 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_968 : src_16; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1163 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_969 : src_17; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1164 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_970 : src_18; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1165 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_971 : src_19; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1166 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_972 : src_20; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1167 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_973 : src_21; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1168 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_974 : src_22; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1169 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_975 : src_23; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1170 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_976 : src_24; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1171 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_977 : src_25; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1172 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_978 : src_26; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1173 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_979 : src_27; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1174 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_980 : src_28; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1175 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_981 : src_29; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1176 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_982 : src_30; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1177 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_983 : src_31; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1178 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_984 : src_32; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1179 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_985 : src_33; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1180 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_986 : src_34; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1181 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_987 : src_35; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1182 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_988 : src_36; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1183 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_989 : src_37; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1184 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_990 : src_38; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1185 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_991 : src_39; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1186 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_992 : src_40; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1187 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_993 : src_41; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1188 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_994 : src_42; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1189 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_995 : src_43; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1190 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_996 : src_44; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1191 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_997 : src_45; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1192 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_998 : src_46; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1193 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_999 : src_47; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1194 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1000 : src_48; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1195 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1001 : src_49; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1196 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1002 : src_50; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1197 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1003 : src_51; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1198 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1004 : src_52; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1199 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1005 : src_53; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1200 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1006 : src_54; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1201 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1007 : src_55; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1202 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1008 : src_56; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1203 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1009 : src_57; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1204 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1010 : src_58; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1205 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1011 : src_59; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1206 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1012 : src_60; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1207 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1013 : src_61; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1208 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1014 : src_62; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1209 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1015 : src_63; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_1210 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1016 : dest_0; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1211 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1017 : dest_1; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1212 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1018 : dest_2; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1213 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1019 : dest_3; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1214 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1020 : dest_4; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1215 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1021 : dest_5; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1216 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1022 : dest_6; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1217 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1023 : dest_7; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1218 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1024 : dest_8; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1219 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1025 : dest_9; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1220 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1026 : dest_10; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1221 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1027 : dest_11; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1222 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1028 : dest_12; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1223 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1029 : dest_13; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1224 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1030 : dest_14; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1225 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1031 : dest_15; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1226 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1032 : dest_16; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1227 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1033 : dest_17; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1228 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1034 : dest_18; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1229 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1035 : dest_19; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1230 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1036 : dest_20; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1231 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1037 : dest_21; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1232 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1038 : dest_22; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1233 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1039 : dest_23; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1234 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1040 : dest_24; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1235 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1041 : dest_25; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1236 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1042 : dest_26; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1237 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1043 : dest_27; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1238 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1044 : dest_28; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1239 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1045 : dest_29; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1240 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1046 : dest_30; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1241 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1047 : dest_31; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1242 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1048 : dest_32; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1243 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1049 : dest_33; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1244 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1050 : dest_34; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1245 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1051 : dest_35; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1246 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1052 : dest_36; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1247 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1053 : dest_37; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1248 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1054 : dest_38; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1249 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1055 : dest_39; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1250 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1056 : dest_40; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1251 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1057 : dest_41; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1252 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1058 : dest_42; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1253 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1059 : dest_43; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1254 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1060 : dest_44; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1255 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1061 : dest_45; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1256 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1062 : dest_46; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1257 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1063 : dest_47; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1258 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1064 : dest_48; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1259 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1065 : dest_49; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1260 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1066 : dest_50; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1261 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1067 : dest_51; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1262 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1068 : dest_52; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1263 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1069 : dest_53; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1264 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1070 : dest_54; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1265 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1071 : dest_55; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1266 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1072 : dest_56; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1267 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1073 : dest_57; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1268 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1074 : dest_58; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1269 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1075 : dest_59; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1270 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1076 : dest_60; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1271 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1077 : dest_61; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1272 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1078 : dest_62; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_1273 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1079 : dest_63; // @[Muxes.scala 34:23 54:70]
  wire [31:0] _GEN_1274 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_1081 : counter; // @[Muxes.scala 31:26 54:70]
  wire [31:0] _j_T_1 = j + 32'h1; // @[Muxes.scala 79:16]
  wire [31:0] _i_T_1 = i + 32'h1; // @[Muxes.scala 85:18]
  wire [31:0] _GEN_1275 = i < 32'h7 ? _i_T_1 : i; // @[Muxes.scala 84:42 85:13 28:20]
  wire  _GEN_1276 = _T_91 | jValid; // @[Muxes.scala 80:83 81:16 27:25]
  reg [31:0] jNext; // @[Muxes.scala 105:24]
  wire [31:0] _k_T_1 = k + 32'h1; // @[Muxes.scala 114:14]
  assign io_i_mux_bus_0 = mux_0; // @[Muxes.scala 35:18]
  assign io_i_mux_bus_1 = mux_1; // @[Muxes.scala 35:18]
  assign io_i_mux_bus_2 = mux_2; // @[Muxes.scala 35:18]
  assign io_i_mux_bus_3 = mux_3; // @[Muxes.scala 35:18]
  assign io_Source_0 = src_0; // @[Muxes.scala 36:15]
  assign io_Source_1 = src_1; // @[Muxes.scala 36:15]
  assign io_Source_2 = src_2; // @[Muxes.scala 36:15]
  assign io_Source_3 = src_3; // @[Muxes.scala 36:15]
  assign io_destination_0 = dest_0; // @[Muxes.scala 37:20]
  assign io_destination_1 = dest_1; // @[Muxes.scala 37:20]
  assign io_destination_2 = dest_2; // @[Muxes.scala 37:20]
  assign io_destination_3 = dest_3; // @[Muxes.scala 37:20]
  assign io_valid = k != 32'h0 & _T_89 & _T_90 & jNext == 32'h6; // @[Muxes.scala 108:86]
  always @(posedge clock) begin
    prevStationary_matrix_0_0 <= io_mat1_0_0; // @[Muxes.scala 19:40]
    prevStationary_matrix_0_1 <= io_mat1_0_1; // @[Muxes.scala 19:40]
    prevStationary_matrix_0_2 <= io_mat1_0_2; // @[Muxes.scala 19:40]
    prevStationary_matrix_0_3 <= io_mat1_0_3; // @[Muxes.scala 19:40]
    prevStationary_matrix_0_4 <= io_mat1_0_4; // @[Muxes.scala 19:40]
    prevStationary_matrix_0_5 <= io_mat1_0_5; // @[Muxes.scala 19:40]
    prevStationary_matrix_0_6 <= io_mat1_0_6; // @[Muxes.scala 19:40]
    prevStationary_matrix_0_7 <= io_mat1_0_7; // @[Muxes.scala 19:40]
    prevStationary_matrix_1_0 <= io_mat1_1_0; // @[Muxes.scala 19:40]
    prevStationary_matrix_1_1 <= io_mat1_1_1; // @[Muxes.scala 19:40]
    prevStationary_matrix_1_2 <= io_mat1_1_2; // @[Muxes.scala 19:40]
    prevStationary_matrix_1_3 <= io_mat1_1_3; // @[Muxes.scala 19:40]
    prevStationary_matrix_1_4 <= io_mat1_1_4; // @[Muxes.scala 19:40]
    prevStationary_matrix_1_5 <= io_mat1_1_5; // @[Muxes.scala 19:40]
    prevStationary_matrix_1_6 <= io_mat1_1_6; // @[Muxes.scala 19:40]
    prevStationary_matrix_1_7 <= io_mat1_1_7; // @[Muxes.scala 19:40]
    prevStationary_matrix_2_0 <= io_mat1_2_0; // @[Muxes.scala 19:40]
    prevStationary_matrix_2_1 <= io_mat1_2_1; // @[Muxes.scala 19:40]
    prevStationary_matrix_2_2 <= io_mat1_2_2; // @[Muxes.scala 19:40]
    prevStationary_matrix_2_3 <= io_mat1_2_3; // @[Muxes.scala 19:40]
    prevStationary_matrix_2_4 <= io_mat1_2_4; // @[Muxes.scala 19:40]
    prevStationary_matrix_2_5 <= io_mat1_2_5; // @[Muxes.scala 19:40]
    prevStationary_matrix_2_6 <= io_mat1_2_6; // @[Muxes.scala 19:40]
    prevStationary_matrix_2_7 <= io_mat1_2_7; // @[Muxes.scala 19:40]
    prevStationary_matrix_3_0 <= io_mat1_3_0; // @[Muxes.scala 19:40]
    prevStationary_matrix_3_1 <= io_mat1_3_1; // @[Muxes.scala 19:40]
    prevStationary_matrix_3_2 <= io_mat1_3_2; // @[Muxes.scala 19:40]
    prevStationary_matrix_3_3 <= io_mat1_3_3; // @[Muxes.scala 19:40]
    prevStationary_matrix_3_4 <= io_mat1_3_4; // @[Muxes.scala 19:40]
    prevStationary_matrix_3_5 <= io_mat1_3_5; // @[Muxes.scala 19:40]
    prevStationary_matrix_3_6 <= io_mat1_3_6; // @[Muxes.scala 19:40]
    prevStationary_matrix_3_7 <= io_mat1_3_7; // @[Muxes.scala 19:40]
    prevStationary_matrix_4_0 <= io_mat1_4_0; // @[Muxes.scala 19:40]
    prevStationary_matrix_4_1 <= io_mat1_4_1; // @[Muxes.scala 19:40]
    prevStationary_matrix_4_2 <= io_mat1_4_2; // @[Muxes.scala 19:40]
    prevStationary_matrix_4_3 <= io_mat1_4_3; // @[Muxes.scala 19:40]
    prevStationary_matrix_4_4 <= io_mat1_4_4; // @[Muxes.scala 19:40]
    prevStationary_matrix_4_5 <= io_mat1_4_5; // @[Muxes.scala 19:40]
    prevStationary_matrix_4_6 <= io_mat1_4_6; // @[Muxes.scala 19:40]
    prevStationary_matrix_4_7 <= io_mat1_4_7; // @[Muxes.scala 19:40]
    prevStationary_matrix_5_0 <= io_mat1_5_0; // @[Muxes.scala 19:40]
    prevStationary_matrix_5_1 <= io_mat1_5_1; // @[Muxes.scala 19:40]
    prevStationary_matrix_5_2 <= io_mat1_5_2; // @[Muxes.scala 19:40]
    prevStationary_matrix_5_3 <= io_mat1_5_3; // @[Muxes.scala 19:40]
    prevStationary_matrix_5_4 <= io_mat1_5_4; // @[Muxes.scala 19:40]
    prevStationary_matrix_5_5 <= io_mat1_5_5; // @[Muxes.scala 19:40]
    prevStationary_matrix_5_6 <= io_mat1_5_6; // @[Muxes.scala 19:40]
    prevStationary_matrix_5_7 <= io_mat1_5_7; // @[Muxes.scala 19:40]
    prevStationary_matrix_6_0 <= io_mat1_6_0; // @[Muxes.scala 19:40]
    prevStationary_matrix_6_1 <= io_mat1_6_1; // @[Muxes.scala 19:40]
    prevStationary_matrix_6_2 <= io_mat1_6_2; // @[Muxes.scala 19:40]
    prevStationary_matrix_6_3 <= io_mat1_6_3; // @[Muxes.scala 19:40]
    prevStationary_matrix_6_4 <= io_mat1_6_4; // @[Muxes.scala 19:40]
    prevStationary_matrix_6_5 <= io_mat1_6_5; // @[Muxes.scala 19:40]
    prevStationary_matrix_6_6 <= io_mat1_6_6; // @[Muxes.scala 19:40]
    prevStationary_matrix_6_7 <= io_mat1_6_7; // @[Muxes.scala 19:40]
    prevStationary_matrix_7_0 <= io_mat1_7_0; // @[Muxes.scala 19:40]
    prevStationary_matrix_7_1 <= io_mat1_7_1; // @[Muxes.scala 19:40]
    prevStationary_matrix_7_2 <= io_mat1_7_2; // @[Muxes.scala 19:40]
    prevStationary_matrix_7_3 <= io_mat1_7_3; // @[Muxes.scala 19:40]
    prevStationary_matrix_7_4 <= io_mat1_7_4; // @[Muxes.scala 19:40]
    prevStationary_matrix_7_5 <= io_mat1_7_5; // @[Muxes.scala 19:40]
    prevStationary_matrix_7_6 <= io_mat1_7_6; // @[Muxes.scala 19:40]
    prevStationary_matrix_7_7 <= io_mat1_7_7; // @[Muxes.scala 19:40]
    prevStreaming_matrix_0 <= io_mat2_0; // @[Muxes.scala 20:39]
    prevStreaming_matrix_1 <= io_mat2_1; // @[Muxes.scala 20:39]
    prevStreaming_matrix_2 <= io_mat2_2; // @[Muxes.scala 20:39]
    prevStreaming_matrix_3 <= io_mat2_3; // @[Muxes.scala 20:39]
    prevStreaming_matrix_4 <= io_mat2_4; // @[Muxes.scala 20:39]
    prevStreaming_matrix_5 <= io_mat2_5; // @[Muxes.scala 20:39]
    prevStreaming_matrix_6 <= io_mat2_6; // @[Muxes.scala 20:39]
    prevStreaming_matrix_7 <= io_mat2_7; // @[Muxes.scala 20:39]
    if (io_mat2_7 != prevStreaming_matrix_7) begin // @[Muxes.scala 49:51]
      matricesAreEqual <= 1'h0; // @[Muxes.scala 50:26]
    end else if (io_mat1_7_7 != prevStationary_matrix_7_7) begin // @[Muxes.scala 45:61]
      matricesAreEqual <= 1'h0; // @[Muxes.scala 46:28]
    end else if (io_mat1_7_6 != prevStationary_matrix_7_6) begin // @[Muxes.scala 45:61]
      matricesAreEqual <= 1'h0; // @[Muxes.scala 46:28]
    end else if (io_mat1_7_5 != prevStationary_matrix_7_5) begin // @[Muxes.scala 45:61]
      matricesAreEqual <= 1'h0; // @[Muxes.scala 46:28]
    end else begin
      matricesAreEqual <= _GEN_67;
    end
    if (reset) begin // @[Muxes.scala 27:25]
      jValid <= 1'h0; // @[Muxes.scala 27:25]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      if (!(j < 32'h7)) begin // @[Muxes.scala 78:40]
        jValid <= _GEN_1276;
      end
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      jValid <= 1'h0; // @[Muxes.scala 93:14]
    end
    if (reset) begin // @[Muxes.scala 28:20]
      i <= 32'h0; // @[Muxes.scala 28:20]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      if (!(j < 32'h7)) begin // @[Muxes.scala 78:40]
        if (!(_T_91)) begin // @[Muxes.scala 80:83]
          i <= _GEN_1275;
        end
      end
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      i <= 32'h0; // @[Muxes.scala 91:9]
    end
    if (reset) begin // @[Muxes.scala 29:20]
      j <= 32'h0; // @[Muxes.scala 29:20]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      if (j < 32'h7) begin // @[Muxes.scala 78:40]
        j <= _j_T_1; // @[Muxes.scala 79:11]
      end else if (!(_T_91)) begin // @[Muxes.scala 80:83]
        j <= 32'h0; // @[Muxes.scala 83:11]
      end
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      j <= 32'h0; // @[Muxes.scala 92:9]
    end
    if (reset) begin // @[Muxes.scala 30:20]
      k <= 32'h0; // @[Muxes.scala 30:20]
    end else if (_T_90 & _T_89) begin // @[Muxes.scala 113:76]
      k <= _k_T_1; // @[Muxes.scala 114:9]
    end
    if (reset) begin // @[Muxes.scala 31:26]
      counter <= 32'h0; // @[Muxes.scala 31:26]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      counter <= _GEN_1274;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      counter <= 32'h0; // @[Muxes.scala 94:15]
    end else begin
      counter <= _GEN_1274;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_0 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_0 <= _GEN_1082;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_0 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_0 <= _GEN_1082;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_1 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_1 <= _GEN_1083;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_1 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_1 <= _GEN_1083;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_2 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_2 <= _GEN_1084;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_2 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_2 <= _GEN_1084;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_3 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_3 <= _GEN_1085;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_3 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_3 <= _GEN_1085;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_4 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_4 <= _GEN_1086;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_4 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_4 <= _GEN_1086;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_5 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_5 <= _GEN_1087;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_5 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_5 <= _GEN_1087;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_6 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_6 <= _GEN_1088;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_6 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_6 <= _GEN_1088;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_7 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_7 <= _GEN_1089;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_7 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_7 <= _GEN_1089;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_8 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_8 <= _GEN_1090;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_8 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_8 <= _GEN_1090;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_9 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_9 <= _GEN_1091;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_9 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_9 <= _GEN_1091;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_10 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_10 <= _GEN_1092;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_10 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_10 <= _GEN_1092;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_11 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_11 <= _GEN_1093;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_11 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_11 <= _GEN_1093;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_12 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_12 <= _GEN_1094;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_12 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_12 <= _GEN_1094;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_13 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_13 <= _GEN_1095;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_13 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_13 <= _GEN_1095;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_14 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_14 <= _GEN_1096;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_14 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_14 <= _GEN_1096;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_15 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_15 <= _GEN_1097;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_15 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_15 <= _GEN_1097;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_16 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_16 <= _GEN_1098;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_16 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_16 <= _GEN_1098;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_17 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_17 <= _GEN_1099;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_17 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_17 <= _GEN_1099;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_18 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_18 <= _GEN_1100;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_18 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_18 <= _GEN_1100;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_19 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_19 <= _GEN_1101;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_19 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_19 <= _GEN_1101;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_20 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_20 <= _GEN_1102;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_20 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_20 <= _GEN_1102;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_21 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_21 <= _GEN_1103;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_21 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_21 <= _GEN_1103;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_22 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_22 <= _GEN_1104;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_22 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_22 <= _GEN_1104;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_23 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_23 <= _GEN_1105;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_23 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_23 <= _GEN_1105;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_24 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_24 <= _GEN_1106;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_24 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_24 <= _GEN_1106;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_25 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_25 <= _GEN_1107;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_25 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_25 <= _GEN_1107;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_26 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_26 <= _GEN_1108;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_26 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_26 <= _GEN_1108;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_27 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_27 <= _GEN_1109;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_27 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_27 <= _GEN_1109;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_28 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_28 <= _GEN_1110;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_28 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_28 <= _GEN_1110;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_29 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_29 <= _GEN_1111;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_29 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_29 <= _GEN_1111;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_30 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_30 <= _GEN_1112;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_30 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_30 <= _GEN_1112;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_31 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_31 <= _GEN_1113;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_31 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_31 <= _GEN_1113;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_32 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_32 <= _GEN_1114;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_32 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_32 <= _GEN_1114;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_33 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_33 <= _GEN_1115;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_33 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_33 <= _GEN_1115;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_34 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_34 <= _GEN_1116;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_34 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_34 <= _GEN_1116;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_35 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_35 <= _GEN_1117;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_35 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_35 <= _GEN_1117;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_36 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_36 <= _GEN_1118;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_36 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_36 <= _GEN_1118;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_37 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_37 <= _GEN_1119;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_37 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_37 <= _GEN_1119;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_38 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_38 <= _GEN_1120;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_38 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_38 <= _GEN_1120;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_39 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_39 <= _GEN_1121;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_39 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_39 <= _GEN_1121;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_40 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_40 <= _GEN_1122;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_40 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_40 <= _GEN_1122;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_41 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_41 <= _GEN_1123;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_41 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_41 <= _GEN_1123;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_42 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_42 <= _GEN_1124;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_42 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_42 <= _GEN_1124;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_43 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_43 <= _GEN_1125;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_43 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_43 <= _GEN_1125;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_44 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_44 <= _GEN_1126;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_44 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_44 <= _GEN_1126;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_45 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_45 <= _GEN_1127;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_45 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_45 <= _GEN_1127;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_46 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_46 <= _GEN_1128;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_46 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_46 <= _GEN_1128;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_47 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_47 <= _GEN_1129;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_47 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_47 <= _GEN_1129;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_48 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_48 <= _GEN_1130;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_48 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_48 <= _GEN_1130;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_49 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_49 <= _GEN_1131;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_49 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_49 <= _GEN_1131;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_50 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_50 <= _GEN_1132;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_50 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_50 <= _GEN_1132;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_51 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_51 <= _GEN_1133;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_51 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_51 <= _GEN_1133;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_52 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_52 <= _GEN_1134;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_52 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_52 <= _GEN_1134;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_53 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_53 <= _GEN_1135;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_53 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_53 <= _GEN_1135;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_54 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_54 <= _GEN_1136;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_54 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_54 <= _GEN_1136;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_55 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_55 <= _GEN_1137;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_55 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_55 <= _GEN_1137;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_56 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_56 <= _GEN_1138;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_56 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_56 <= _GEN_1138;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_57 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_57 <= _GEN_1139;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_57 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_57 <= _GEN_1139;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_58 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_58 <= _GEN_1140;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_58 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_58 <= _GEN_1140;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_59 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_59 <= _GEN_1141;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_59 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_59 <= _GEN_1141;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_60 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_60 <= _GEN_1142;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_60 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_60 <= _GEN_1142;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_61 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_61 <= _GEN_1143;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_61 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_61 <= _GEN_1143;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_62 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_62 <= _GEN_1144;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_62 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_62 <= _GEN_1144;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_63 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_63 <= _GEN_1145;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_63 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_63 <= _GEN_1145;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_0 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_0 <= _GEN_1146;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_0 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_0 <= _GEN_1146;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_1 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_1 <= _GEN_1147;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_1 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_1 <= _GEN_1147;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_2 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_2 <= _GEN_1148;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_2 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_2 <= _GEN_1148;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_3 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_3 <= _GEN_1149;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_3 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_3 <= _GEN_1149;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_4 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_4 <= _GEN_1150;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_4 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_4 <= _GEN_1150;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_5 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_5 <= _GEN_1151;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_5 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_5 <= _GEN_1151;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_6 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_6 <= _GEN_1152;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_6 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_6 <= _GEN_1152;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_7 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_7 <= _GEN_1153;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_7 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_7 <= _GEN_1153;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_8 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_8 <= _GEN_1154;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_8 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_8 <= _GEN_1154;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_9 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_9 <= _GEN_1155;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_9 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_9 <= _GEN_1155;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_10 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_10 <= _GEN_1156;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_10 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_10 <= _GEN_1156;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_11 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_11 <= _GEN_1157;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_11 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_11 <= _GEN_1157;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_12 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_12 <= _GEN_1158;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_12 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_12 <= _GEN_1158;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_13 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_13 <= _GEN_1159;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_13 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_13 <= _GEN_1159;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_14 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_14 <= _GEN_1160;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_14 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_14 <= _GEN_1160;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_15 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_15 <= _GEN_1161;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_15 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_15 <= _GEN_1161;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_16 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_16 <= _GEN_1162;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_16 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_16 <= _GEN_1162;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_17 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_17 <= _GEN_1163;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_17 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_17 <= _GEN_1163;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_18 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_18 <= _GEN_1164;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_18 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_18 <= _GEN_1164;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_19 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_19 <= _GEN_1165;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_19 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_19 <= _GEN_1165;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_20 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_20 <= _GEN_1166;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_20 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_20 <= _GEN_1166;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_21 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_21 <= _GEN_1167;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_21 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_21 <= _GEN_1167;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_22 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_22 <= _GEN_1168;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_22 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_22 <= _GEN_1168;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_23 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_23 <= _GEN_1169;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_23 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_23 <= _GEN_1169;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_24 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_24 <= _GEN_1170;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_24 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_24 <= _GEN_1170;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_25 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_25 <= _GEN_1171;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_25 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_25 <= _GEN_1171;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_26 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_26 <= _GEN_1172;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_26 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_26 <= _GEN_1172;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_27 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_27 <= _GEN_1173;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_27 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_27 <= _GEN_1173;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_28 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_28 <= _GEN_1174;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_28 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_28 <= _GEN_1174;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_29 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_29 <= _GEN_1175;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_29 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_29 <= _GEN_1175;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_30 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_30 <= _GEN_1176;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_30 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_30 <= _GEN_1176;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_31 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_31 <= _GEN_1177;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_31 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_31 <= _GEN_1177;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_32 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_32 <= _GEN_1178;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_32 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_32 <= _GEN_1178;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_33 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_33 <= _GEN_1179;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_33 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_33 <= _GEN_1179;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_34 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_34 <= _GEN_1180;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_34 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_34 <= _GEN_1180;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_35 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_35 <= _GEN_1181;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_35 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_35 <= _GEN_1181;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_36 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_36 <= _GEN_1182;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_36 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_36 <= _GEN_1182;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_37 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_37 <= _GEN_1183;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_37 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_37 <= _GEN_1183;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_38 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_38 <= _GEN_1184;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_38 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_38 <= _GEN_1184;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_39 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_39 <= _GEN_1185;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_39 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_39 <= _GEN_1185;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_40 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_40 <= _GEN_1186;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_40 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_40 <= _GEN_1186;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_41 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_41 <= _GEN_1187;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_41 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_41 <= _GEN_1187;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_42 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_42 <= _GEN_1188;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_42 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_42 <= _GEN_1188;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_43 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_43 <= _GEN_1189;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_43 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_43 <= _GEN_1189;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_44 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_44 <= _GEN_1190;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_44 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_44 <= _GEN_1190;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_45 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_45 <= _GEN_1191;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_45 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_45 <= _GEN_1191;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_46 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_46 <= _GEN_1192;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_46 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_46 <= _GEN_1192;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_47 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_47 <= _GEN_1193;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_47 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_47 <= _GEN_1193;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_48 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_48 <= _GEN_1194;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_48 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_48 <= _GEN_1194;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_49 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_49 <= _GEN_1195;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_49 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_49 <= _GEN_1195;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_50 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_50 <= _GEN_1196;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_50 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_50 <= _GEN_1196;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_51 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_51 <= _GEN_1197;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_51 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_51 <= _GEN_1197;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_52 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_52 <= _GEN_1198;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_52 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_52 <= _GEN_1198;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_53 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_53 <= _GEN_1199;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_53 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_53 <= _GEN_1199;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_54 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_54 <= _GEN_1200;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_54 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_54 <= _GEN_1200;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_55 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_55 <= _GEN_1201;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_55 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_55 <= _GEN_1201;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_56 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_56 <= _GEN_1202;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_56 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_56 <= _GEN_1202;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_57 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_57 <= _GEN_1203;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_57 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_57 <= _GEN_1203;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_58 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_58 <= _GEN_1204;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_58 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_58 <= _GEN_1204;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_59 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_59 <= _GEN_1205;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_59 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_59 <= _GEN_1205;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_60 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_60 <= _GEN_1206;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_60 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_60 <= _GEN_1206;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_61 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_61 <= _GEN_1207;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_61 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_61 <= _GEN_1207;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_62 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_62 <= _GEN_1208;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_62 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_62 <= _GEN_1208;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_63 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_63 <= _GEN_1209;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_63 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_63 <= _GEN_1209;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_0 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_0 <= _GEN_1210;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_0 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_0 <= _GEN_1210;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_1 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_1 <= _GEN_1211;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_1 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_1 <= _GEN_1211;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_2 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_2 <= _GEN_1212;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_2 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_2 <= _GEN_1212;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_3 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_3 <= _GEN_1213;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_3 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_3 <= _GEN_1213;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_4 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_4 <= _GEN_1214;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_4 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_4 <= _GEN_1214;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_5 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_5 <= _GEN_1215;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_5 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_5 <= _GEN_1215;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_6 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_6 <= _GEN_1216;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_6 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_6 <= _GEN_1216;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_7 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_7 <= _GEN_1217;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_7 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_7 <= _GEN_1217;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_8 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_8 <= _GEN_1218;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_8 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_8 <= _GEN_1218;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_9 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_9 <= _GEN_1219;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_9 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_9 <= _GEN_1219;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_10 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_10 <= _GEN_1220;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_10 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_10 <= _GEN_1220;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_11 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_11 <= _GEN_1221;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_11 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_11 <= _GEN_1221;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_12 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_12 <= _GEN_1222;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_12 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_12 <= _GEN_1222;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_13 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_13 <= _GEN_1223;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_13 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_13 <= _GEN_1223;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_14 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_14 <= _GEN_1224;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_14 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_14 <= _GEN_1224;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_15 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_15 <= _GEN_1225;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_15 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_15 <= _GEN_1225;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_16 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_16 <= _GEN_1226;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_16 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_16 <= _GEN_1226;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_17 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_17 <= _GEN_1227;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_17 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_17 <= _GEN_1227;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_18 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_18 <= _GEN_1228;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_18 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_18 <= _GEN_1228;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_19 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_19 <= _GEN_1229;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_19 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_19 <= _GEN_1229;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_20 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_20 <= _GEN_1230;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_20 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_20 <= _GEN_1230;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_21 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_21 <= _GEN_1231;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_21 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_21 <= _GEN_1231;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_22 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_22 <= _GEN_1232;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_22 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_22 <= _GEN_1232;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_23 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_23 <= _GEN_1233;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_23 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_23 <= _GEN_1233;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_24 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_24 <= _GEN_1234;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_24 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_24 <= _GEN_1234;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_25 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_25 <= _GEN_1235;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_25 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_25 <= _GEN_1235;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_26 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_26 <= _GEN_1236;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_26 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_26 <= _GEN_1236;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_27 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_27 <= _GEN_1237;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_27 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_27 <= _GEN_1237;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_28 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_28 <= _GEN_1238;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_28 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_28 <= _GEN_1238;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_29 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_29 <= _GEN_1239;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_29 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_29 <= _GEN_1239;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_30 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_30 <= _GEN_1240;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_30 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_30 <= _GEN_1240;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_31 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_31 <= _GEN_1241;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_31 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_31 <= _GEN_1241;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_32 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_32 <= _GEN_1242;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_32 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_32 <= _GEN_1242;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_33 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_33 <= _GEN_1243;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_33 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_33 <= _GEN_1243;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_34 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_34 <= _GEN_1244;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_34 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_34 <= _GEN_1244;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_35 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_35 <= _GEN_1245;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_35 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_35 <= _GEN_1245;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_36 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_36 <= _GEN_1246;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_36 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_36 <= _GEN_1246;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_37 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_37 <= _GEN_1247;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_37 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_37 <= _GEN_1247;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_38 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_38 <= _GEN_1248;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_38 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_38 <= _GEN_1248;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_39 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_39 <= _GEN_1249;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_39 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_39 <= _GEN_1249;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_40 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_40 <= _GEN_1250;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_40 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_40 <= _GEN_1250;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_41 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_41 <= _GEN_1251;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_41 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_41 <= _GEN_1251;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_42 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_42 <= _GEN_1252;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_42 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_42 <= _GEN_1252;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_43 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_43 <= _GEN_1253;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_43 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_43 <= _GEN_1253;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_44 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_44 <= _GEN_1254;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_44 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_44 <= _GEN_1254;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_45 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_45 <= _GEN_1255;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_45 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_45 <= _GEN_1255;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_46 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_46 <= _GEN_1256;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_46 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_46 <= _GEN_1256;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_47 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_47 <= _GEN_1257;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_47 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_47 <= _GEN_1257;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_48 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_48 <= _GEN_1258;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_48 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_48 <= _GEN_1258;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_49 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_49 <= _GEN_1259;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_49 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_49 <= _GEN_1259;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_50 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_50 <= _GEN_1260;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_50 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_50 <= _GEN_1260;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_51 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_51 <= _GEN_1261;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_51 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_51 <= _GEN_1261;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_52 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_52 <= _GEN_1262;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_52 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_52 <= _GEN_1262;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_53 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_53 <= _GEN_1263;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_53 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_53 <= _GEN_1263;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_54 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_54 <= _GEN_1264;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_54 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_54 <= _GEN_1264;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_55 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_55 <= _GEN_1265;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_55 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_55 <= _GEN_1265;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_56 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_56 <= _GEN_1266;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_56 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_56 <= _GEN_1266;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_57 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_57 <= _GEN_1267;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_57 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_57 <= _GEN_1267;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_58 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_58 <= _GEN_1268;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_58 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_58 <= _GEN_1268;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_59 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_59 <= _GEN_1269;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_59 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_59 <= _GEN_1269;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_60 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_60 <= _GEN_1270;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_60 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_60 <= _GEN_1270;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_61 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_61 <= _GEN_1271;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_61 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_61 <= _GEN_1271;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_62 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_62 <= _GEN_1272;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_62 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_62 <= _GEN_1272;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_63 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_63 <= _GEN_1273;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_63 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_63 <= _GEN_1273;
    end
    if (reset) begin // @[Muxes.scala 105:24]
      jNext <= 32'h0; // @[Muxes.scala 105:24]
    end else begin
      jNext <= j; // @[Muxes.scala 106:11]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  prevStationary_matrix_0_0 = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  prevStationary_matrix_0_1 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  prevStationary_matrix_0_2 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  prevStationary_matrix_0_3 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  prevStationary_matrix_0_4 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  prevStationary_matrix_0_5 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  prevStationary_matrix_0_6 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  prevStationary_matrix_0_7 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  prevStationary_matrix_1_0 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  prevStationary_matrix_1_1 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  prevStationary_matrix_1_2 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  prevStationary_matrix_1_3 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  prevStationary_matrix_1_4 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  prevStationary_matrix_1_5 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  prevStationary_matrix_1_6 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  prevStationary_matrix_1_7 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  prevStationary_matrix_2_0 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  prevStationary_matrix_2_1 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  prevStationary_matrix_2_2 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  prevStationary_matrix_2_3 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  prevStationary_matrix_2_4 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  prevStationary_matrix_2_5 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  prevStationary_matrix_2_6 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  prevStationary_matrix_2_7 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  prevStationary_matrix_3_0 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  prevStationary_matrix_3_1 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  prevStationary_matrix_3_2 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  prevStationary_matrix_3_3 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  prevStationary_matrix_3_4 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  prevStationary_matrix_3_5 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  prevStationary_matrix_3_6 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  prevStationary_matrix_3_7 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  prevStationary_matrix_4_0 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  prevStationary_matrix_4_1 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  prevStationary_matrix_4_2 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  prevStationary_matrix_4_3 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  prevStationary_matrix_4_4 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  prevStationary_matrix_4_5 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  prevStationary_matrix_4_6 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  prevStationary_matrix_4_7 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  prevStationary_matrix_5_0 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  prevStationary_matrix_5_1 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  prevStationary_matrix_5_2 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  prevStationary_matrix_5_3 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  prevStationary_matrix_5_4 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  prevStationary_matrix_5_5 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  prevStationary_matrix_5_6 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  prevStationary_matrix_5_7 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  prevStationary_matrix_6_0 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  prevStationary_matrix_6_1 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  prevStationary_matrix_6_2 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  prevStationary_matrix_6_3 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  prevStationary_matrix_6_4 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  prevStationary_matrix_6_5 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  prevStationary_matrix_6_6 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  prevStationary_matrix_6_7 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  prevStationary_matrix_7_0 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  prevStationary_matrix_7_1 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  prevStationary_matrix_7_2 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  prevStationary_matrix_7_3 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  prevStationary_matrix_7_4 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  prevStationary_matrix_7_5 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  prevStationary_matrix_7_6 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  prevStationary_matrix_7_7 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  prevStreaming_matrix_0 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  prevStreaming_matrix_1 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  prevStreaming_matrix_2 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  prevStreaming_matrix_3 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  prevStreaming_matrix_4 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  prevStreaming_matrix_5 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  prevStreaming_matrix_6 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  prevStreaming_matrix_7 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  matricesAreEqual = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  jValid = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  i = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  j = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  k = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  counter = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  mux_0 = _RAND_78[3:0];
  _RAND_79 = {1{`RANDOM}};
  mux_1 = _RAND_79[3:0];
  _RAND_80 = {1{`RANDOM}};
  mux_2 = _RAND_80[3:0];
  _RAND_81 = {1{`RANDOM}};
  mux_3 = _RAND_81[3:0];
  _RAND_82 = {1{`RANDOM}};
  mux_4 = _RAND_82[3:0];
  _RAND_83 = {1{`RANDOM}};
  mux_5 = _RAND_83[3:0];
  _RAND_84 = {1{`RANDOM}};
  mux_6 = _RAND_84[3:0];
  _RAND_85 = {1{`RANDOM}};
  mux_7 = _RAND_85[3:0];
  _RAND_86 = {1{`RANDOM}};
  mux_8 = _RAND_86[3:0];
  _RAND_87 = {1{`RANDOM}};
  mux_9 = _RAND_87[3:0];
  _RAND_88 = {1{`RANDOM}};
  mux_10 = _RAND_88[3:0];
  _RAND_89 = {1{`RANDOM}};
  mux_11 = _RAND_89[3:0];
  _RAND_90 = {1{`RANDOM}};
  mux_12 = _RAND_90[3:0];
  _RAND_91 = {1{`RANDOM}};
  mux_13 = _RAND_91[3:0];
  _RAND_92 = {1{`RANDOM}};
  mux_14 = _RAND_92[3:0];
  _RAND_93 = {1{`RANDOM}};
  mux_15 = _RAND_93[3:0];
  _RAND_94 = {1{`RANDOM}};
  mux_16 = _RAND_94[3:0];
  _RAND_95 = {1{`RANDOM}};
  mux_17 = _RAND_95[3:0];
  _RAND_96 = {1{`RANDOM}};
  mux_18 = _RAND_96[3:0];
  _RAND_97 = {1{`RANDOM}};
  mux_19 = _RAND_97[3:0];
  _RAND_98 = {1{`RANDOM}};
  mux_20 = _RAND_98[3:0];
  _RAND_99 = {1{`RANDOM}};
  mux_21 = _RAND_99[3:0];
  _RAND_100 = {1{`RANDOM}};
  mux_22 = _RAND_100[3:0];
  _RAND_101 = {1{`RANDOM}};
  mux_23 = _RAND_101[3:0];
  _RAND_102 = {1{`RANDOM}};
  mux_24 = _RAND_102[3:0];
  _RAND_103 = {1{`RANDOM}};
  mux_25 = _RAND_103[3:0];
  _RAND_104 = {1{`RANDOM}};
  mux_26 = _RAND_104[3:0];
  _RAND_105 = {1{`RANDOM}};
  mux_27 = _RAND_105[3:0];
  _RAND_106 = {1{`RANDOM}};
  mux_28 = _RAND_106[3:0];
  _RAND_107 = {1{`RANDOM}};
  mux_29 = _RAND_107[3:0];
  _RAND_108 = {1{`RANDOM}};
  mux_30 = _RAND_108[3:0];
  _RAND_109 = {1{`RANDOM}};
  mux_31 = _RAND_109[3:0];
  _RAND_110 = {1{`RANDOM}};
  mux_32 = _RAND_110[3:0];
  _RAND_111 = {1{`RANDOM}};
  mux_33 = _RAND_111[3:0];
  _RAND_112 = {1{`RANDOM}};
  mux_34 = _RAND_112[3:0];
  _RAND_113 = {1{`RANDOM}};
  mux_35 = _RAND_113[3:0];
  _RAND_114 = {1{`RANDOM}};
  mux_36 = _RAND_114[3:0];
  _RAND_115 = {1{`RANDOM}};
  mux_37 = _RAND_115[3:0];
  _RAND_116 = {1{`RANDOM}};
  mux_38 = _RAND_116[3:0];
  _RAND_117 = {1{`RANDOM}};
  mux_39 = _RAND_117[3:0];
  _RAND_118 = {1{`RANDOM}};
  mux_40 = _RAND_118[3:0];
  _RAND_119 = {1{`RANDOM}};
  mux_41 = _RAND_119[3:0];
  _RAND_120 = {1{`RANDOM}};
  mux_42 = _RAND_120[3:0];
  _RAND_121 = {1{`RANDOM}};
  mux_43 = _RAND_121[3:0];
  _RAND_122 = {1{`RANDOM}};
  mux_44 = _RAND_122[3:0];
  _RAND_123 = {1{`RANDOM}};
  mux_45 = _RAND_123[3:0];
  _RAND_124 = {1{`RANDOM}};
  mux_46 = _RAND_124[3:0];
  _RAND_125 = {1{`RANDOM}};
  mux_47 = _RAND_125[3:0];
  _RAND_126 = {1{`RANDOM}};
  mux_48 = _RAND_126[3:0];
  _RAND_127 = {1{`RANDOM}};
  mux_49 = _RAND_127[3:0];
  _RAND_128 = {1{`RANDOM}};
  mux_50 = _RAND_128[3:0];
  _RAND_129 = {1{`RANDOM}};
  mux_51 = _RAND_129[3:0];
  _RAND_130 = {1{`RANDOM}};
  mux_52 = _RAND_130[3:0];
  _RAND_131 = {1{`RANDOM}};
  mux_53 = _RAND_131[3:0];
  _RAND_132 = {1{`RANDOM}};
  mux_54 = _RAND_132[3:0];
  _RAND_133 = {1{`RANDOM}};
  mux_55 = _RAND_133[3:0];
  _RAND_134 = {1{`RANDOM}};
  mux_56 = _RAND_134[3:0];
  _RAND_135 = {1{`RANDOM}};
  mux_57 = _RAND_135[3:0];
  _RAND_136 = {1{`RANDOM}};
  mux_58 = _RAND_136[3:0];
  _RAND_137 = {1{`RANDOM}};
  mux_59 = _RAND_137[3:0];
  _RAND_138 = {1{`RANDOM}};
  mux_60 = _RAND_138[3:0];
  _RAND_139 = {1{`RANDOM}};
  mux_61 = _RAND_139[3:0];
  _RAND_140 = {1{`RANDOM}};
  mux_62 = _RAND_140[3:0];
  _RAND_141 = {1{`RANDOM}};
  mux_63 = _RAND_141[3:0];
  _RAND_142 = {1{`RANDOM}};
  src_0 = _RAND_142[15:0];
  _RAND_143 = {1{`RANDOM}};
  src_1 = _RAND_143[15:0];
  _RAND_144 = {1{`RANDOM}};
  src_2 = _RAND_144[15:0];
  _RAND_145 = {1{`RANDOM}};
  src_3 = _RAND_145[15:0];
  _RAND_146 = {1{`RANDOM}};
  src_4 = _RAND_146[15:0];
  _RAND_147 = {1{`RANDOM}};
  src_5 = _RAND_147[15:0];
  _RAND_148 = {1{`RANDOM}};
  src_6 = _RAND_148[15:0];
  _RAND_149 = {1{`RANDOM}};
  src_7 = _RAND_149[15:0];
  _RAND_150 = {1{`RANDOM}};
  src_8 = _RAND_150[15:0];
  _RAND_151 = {1{`RANDOM}};
  src_9 = _RAND_151[15:0];
  _RAND_152 = {1{`RANDOM}};
  src_10 = _RAND_152[15:0];
  _RAND_153 = {1{`RANDOM}};
  src_11 = _RAND_153[15:0];
  _RAND_154 = {1{`RANDOM}};
  src_12 = _RAND_154[15:0];
  _RAND_155 = {1{`RANDOM}};
  src_13 = _RAND_155[15:0];
  _RAND_156 = {1{`RANDOM}};
  src_14 = _RAND_156[15:0];
  _RAND_157 = {1{`RANDOM}};
  src_15 = _RAND_157[15:0];
  _RAND_158 = {1{`RANDOM}};
  src_16 = _RAND_158[15:0];
  _RAND_159 = {1{`RANDOM}};
  src_17 = _RAND_159[15:0];
  _RAND_160 = {1{`RANDOM}};
  src_18 = _RAND_160[15:0];
  _RAND_161 = {1{`RANDOM}};
  src_19 = _RAND_161[15:0];
  _RAND_162 = {1{`RANDOM}};
  src_20 = _RAND_162[15:0];
  _RAND_163 = {1{`RANDOM}};
  src_21 = _RAND_163[15:0];
  _RAND_164 = {1{`RANDOM}};
  src_22 = _RAND_164[15:0];
  _RAND_165 = {1{`RANDOM}};
  src_23 = _RAND_165[15:0];
  _RAND_166 = {1{`RANDOM}};
  src_24 = _RAND_166[15:0];
  _RAND_167 = {1{`RANDOM}};
  src_25 = _RAND_167[15:0];
  _RAND_168 = {1{`RANDOM}};
  src_26 = _RAND_168[15:0];
  _RAND_169 = {1{`RANDOM}};
  src_27 = _RAND_169[15:0];
  _RAND_170 = {1{`RANDOM}};
  src_28 = _RAND_170[15:0];
  _RAND_171 = {1{`RANDOM}};
  src_29 = _RAND_171[15:0];
  _RAND_172 = {1{`RANDOM}};
  src_30 = _RAND_172[15:0];
  _RAND_173 = {1{`RANDOM}};
  src_31 = _RAND_173[15:0];
  _RAND_174 = {1{`RANDOM}};
  src_32 = _RAND_174[15:0];
  _RAND_175 = {1{`RANDOM}};
  src_33 = _RAND_175[15:0];
  _RAND_176 = {1{`RANDOM}};
  src_34 = _RAND_176[15:0];
  _RAND_177 = {1{`RANDOM}};
  src_35 = _RAND_177[15:0];
  _RAND_178 = {1{`RANDOM}};
  src_36 = _RAND_178[15:0];
  _RAND_179 = {1{`RANDOM}};
  src_37 = _RAND_179[15:0];
  _RAND_180 = {1{`RANDOM}};
  src_38 = _RAND_180[15:0];
  _RAND_181 = {1{`RANDOM}};
  src_39 = _RAND_181[15:0];
  _RAND_182 = {1{`RANDOM}};
  src_40 = _RAND_182[15:0];
  _RAND_183 = {1{`RANDOM}};
  src_41 = _RAND_183[15:0];
  _RAND_184 = {1{`RANDOM}};
  src_42 = _RAND_184[15:0];
  _RAND_185 = {1{`RANDOM}};
  src_43 = _RAND_185[15:0];
  _RAND_186 = {1{`RANDOM}};
  src_44 = _RAND_186[15:0];
  _RAND_187 = {1{`RANDOM}};
  src_45 = _RAND_187[15:0];
  _RAND_188 = {1{`RANDOM}};
  src_46 = _RAND_188[15:0];
  _RAND_189 = {1{`RANDOM}};
  src_47 = _RAND_189[15:0];
  _RAND_190 = {1{`RANDOM}};
  src_48 = _RAND_190[15:0];
  _RAND_191 = {1{`RANDOM}};
  src_49 = _RAND_191[15:0];
  _RAND_192 = {1{`RANDOM}};
  src_50 = _RAND_192[15:0];
  _RAND_193 = {1{`RANDOM}};
  src_51 = _RAND_193[15:0];
  _RAND_194 = {1{`RANDOM}};
  src_52 = _RAND_194[15:0];
  _RAND_195 = {1{`RANDOM}};
  src_53 = _RAND_195[15:0];
  _RAND_196 = {1{`RANDOM}};
  src_54 = _RAND_196[15:0];
  _RAND_197 = {1{`RANDOM}};
  src_55 = _RAND_197[15:0];
  _RAND_198 = {1{`RANDOM}};
  src_56 = _RAND_198[15:0];
  _RAND_199 = {1{`RANDOM}};
  src_57 = _RAND_199[15:0];
  _RAND_200 = {1{`RANDOM}};
  src_58 = _RAND_200[15:0];
  _RAND_201 = {1{`RANDOM}};
  src_59 = _RAND_201[15:0];
  _RAND_202 = {1{`RANDOM}};
  src_60 = _RAND_202[15:0];
  _RAND_203 = {1{`RANDOM}};
  src_61 = _RAND_203[15:0];
  _RAND_204 = {1{`RANDOM}};
  src_62 = _RAND_204[15:0];
  _RAND_205 = {1{`RANDOM}};
  src_63 = _RAND_205[15:0];
  _RAND_206 = {1{`RANDOM}};
  dest_0 = _RAND_206[15:0];
  _RAND_207 = {1{`RANDOM}};
  dest_1 = _RAND_207[15:0];
  _RAND_208 = {1{`RANDOM}};
  dest_2 = _RAND_208[15:0];
  _RAND_209 = {1{`RANDOM}};
  dest_3 = _RAND_209[15:0];
  _RAND_210 = {1{`RANDOM}};
  dest_4 = _RAND_210[15:0];
  _RAND_211 = {1{`RANDOM}};
  dest_5 = _RAND_211[15:0];
  _RAND_212 = {1{`RANDOM}};
  dest_6 = _RAND_212[15:0];
  _RAND_213 = {1{`RANDOM}};
  dest_7 = _RAND_213[15:0];
  _RAND_214 = {1{`RANDOM}};
  dest_8 = _RAND_214[15:0];
  _RAND_215 = {1{`RANDOM}};
  dest_9 = _RAND_215[15:0];
  _RAND_216 = {1{`RANDOM}};
  dest_10 = _RAND_216[15:0];
  _RAND_217 = {1{`RANDOM}};
  dest_11 = _RAND_217[15:0];
  _RAND_218 = {1{`RANDOM}};
  dest_12 = _RAND_218[15:0];
  _RAND_219 = {1{`RANDOM}};
  dest_13 = _RAND_219[15:0];
  _RAND_220 = {1{`RANDOM}};
  dest_14 = _RAND_220[15:0];
  _RAND_221 = {1{`RANDOM}};
  dest_15 = _RAND_221[15:0];
  _RAND_222 = {1{`RANDOM}};
  dest_16 = _RAND_222[15:0];
  _RAND_223 = {1{`RANDOM}};
  dest_17 = _RAND_223[15:0];
  _RAND_224 = {1{`RANDOM}};
  dest_18 = _RAND_224[15:0];
  _RAND_225 = {1{`RANDOM}};
  dest_19 = _RAND_225[15:0];
  _RAND_226 = {1{`RANDOM}};
  dest_20 = _RAND_226[15:0];
  _RAND_227 = {1{`RANDOM}};
  dest_21 = _RAND_227[15:0];
  _RAND_228 = {1{`RANDOM}};
  dest_22 = _RAND_228[15:0];
  _RAND_229 = {1{`RANDOM}};
  dest_23 = _RAND_229[15:0];
  _RAND_230 = {1{`RANDOM}};
  dest_24 = _RAND_230[15:0];
  _RAND_231 = {1{`RANDOM}};
  dest_25 = _RAND_231[15:0];
  _RAND_232 = {1{`RANDOM}};
  dest_26 = _RAND_232[15:0];
  _RAND_233 = {1{`RANDOM}};
  dest_27 = _RAND_233[15:0];
  _RAND_234 = {1{`RANDOM}};
  dest_28 = _RAND_234[15:0];
  _RAND_235 = {1{`RANDOM}};
  dest_29 = _RAND_235[15:0];
  _RAND_236 = {1{`RANDOM}};
  dest_30 = _RAND_236[15:0];
  _RAND_237 = {1{`RANDOM}};
  dest_31 = _RAND_237[15:0];
  _RAND_238 = {1{`RANDOM}};
  dest_32 = _RAND_238[15:0];
  _RAND_239 = {1{`RANDOM}};
  dest_33 = _RAND_239[15:0];
  _RAND_240 = {1{`RANDOM}};
  dest_34 = _RAND_240[15:0];
  _RAND_241 = {1{`RANDOM}};
  dest_35 = _RAND_241[15:0];
  _RAND_242 = {1{`RANDOM}};
  dest_36 = _RAND_242[15:0];
  _RAND_243 = {1{`RANDOM}};
  dest_37 = _RAND_243[15:0];
  _RAND_244 = {1{`RANDOM}};
  dest_38 = _RAND_244[15:0];
  _RAND_245 = {1{`RANDOM}};
  dest_39 = _RAND_245[15:0];
  _RAND_246 = {1{`RANDOM}};
  dest_40 = _RAND_246[15:0];
  _RAND_247 = {1{`RANDOM}};
  dest_41 = _RAND_247[15:0];
  _RAND_248 = {1{`RANDOM}};
  dest_42 = _RAND_248[15:0];
  _RAND_249 = {1{`RANDOM}};
  dest_43 = _RAND_249[15:0];
  _RAND_250 = {1{`RANDOM}};
  dest_44 = _RAND_250[15:0];
  _RAND_251 = {1{`RANDOM}};
  dest_45 = _RAND_251[15:0];
  _RAND_252 = {1{`RANDOM}};
  dest_46 = _RAND_252[15:0];
  _RAND_253 = {1{`RANDOM}};
  dest_47 = _RAND_253[15:0];
  _RAND_254 = {1{`RANDOM}};
  dest_48 = _RAND_254[15:0];
  _RAND_255 = {1{`RANDOM}};
  dest_49 = _RAND_255[15:0];
  _RAND_256 = {1{`RANDOM}};
  dest_50 = _RAND_256[15:0];
  _RAND_257 = {1{`RANDOM}};
  dest_51 = _RAND_257[15:0];
  _RAND_258 = {1{`RANDOM}};
  dest_52 = _RAND_258[15:0];
  _RAND_259 = {1{`RANDOM}};
  dest_53 = _RAND_259[15:0];
  _RAND_260 = {1{`RANDOM}};
  dest_54 = _RAND_260[15:0];
  _RAND_261 = {1{`RANDOM}};
  dest_55 = _RAND_261[15:0];
  _RAND_262 = {1{`RANDOM}};
  dest_56 = _RAND_262[15:0];
  _RAND_263 = {1{`RANDOM}};
  dest_57 = _RAND_263[15:0];
  _RAND_264 = {1{`RANDOM}};
  dest_58 = _RAND_264[15:0];
  _RAND_265 = {1{`RANDOM}};
  dest_59 = _RAND_265[15:0];
  _RAND_266 = {1{`RANDOM}};
  dest_60 = _RAND_266[15:0];
  _RAND_267 = {1{`RANDOM}};
  dest_61 = _RAND_267[15:0];
  _RAND_268 = {1{`RANDOM}};
  dest_62 = _RAND_268[15:0];
  _RAND_269 = {1{`RANDOM}};
  dest_63 = _RAND_269[15:0];
  _RAND_270 = {1{`RANDOM}};
  jNext = _RAND_270[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SourceDestination(
  input         clock,
  input         reset,
  input  [15:0] io_Stationary_matrix_0_0,
  input  [15:0] io_Stationary_matrix_0_1,
  input  [15:0] io_Stationary_matrix_0_2,
  input  [15:0] io_Stationary_matrix_0_3,
  input  [15:0] io_Stationary_matrix_0_4,
  input  [15:0] io_Stationary_matrix_0_5,
  input  [15:0] io_Stationary_matrix_0_6,
  input  [15:0] io_Stationary_matrix_0_7,
  input  [15:0] io_Stationary_matrix_1_0,
  input  [15:0] io_Stationary_matrix_1_1,
  input  [15:0] io_Stationary_matrix_1_2,
  input  [15:0] io_Stationary_matrix_1_3,
  input  [15:0] io_Stationary_matrix_1_4,
  input  [15:0] io_Stationary_matrix_1_5,
  input  [15:0] io_Stationary_matrix_1_6,
  input  [15:0] io_Stationary_matrix_1_7,
  input  [15:0] io_Stationary_matrix_2_0,
  input  [15:0] io_Stationary_matrix_2_1,
  input  [15:0] io_Stationary_matrix_2_2,
  input  [15:0] io_Stationary_matrix_2_3,
  input  [15:0] io_Stationary_matrix_2_4,
  input  [15:0] io_Stationary_matrix_2_5,
  input  [15:0] io_Stationary_matrix_2_6,
  input  [15:0] io_Stationary_matrix_2_7,
  input  [15:0] io_Stationary_matrix_3_0,
  input  [15:0] io_Stationary_matrix_3_1,
  input  [15:0] io_Stationary_matrix_3_2,
  input  [15:0] io_Stationary_matrix_3_3,
  input  [15:0] io_Stationary_matrix_3_4,
  input  [15:0] io_Stationary_matrix_3_5,
  input  [15:0] io_Stationary_matrix_3_6,
  input  [15:0] io_Stationary_matrix_3_7,
  input  [15:0] io_Stationary_matrix_4_0,
  input  [15:0] io_Stationary_matrix_4_1,
  input  [15:0] io_Stationary_matrix_4_2,
  input  [15:0] io_Stationary_matrix_4_3,
  input  [15:0] io_Stationary_matrix_4_4,
  input  [15:0] io_Stationary_matrix_4_5,
  input  [15:0] io_Stationary_matrix_4_6,
  input  [15:0] io_Stationary_matrix_4_7,
  input  [15:0] io_Stationary_matrix_5_0,
  input  [15:0] io_Stationary_matrix_5_1,
  input  [15:0] io_Stationary_matrix_5_2,
  input  [15:0] io_Stationary_matrix_5_3,
  input  [15:0] io_Stationary_matrix_5_4,
  input  [15:0] io_Stationary_matrix_5_5,
  input  [15:0] io_Stationary_matrix_5_6,
  input  [15:0] io_Stationary_matrix_5_7,
  input  [15:0] io_Stationary_matrix_6_0,
  input  [15:0] io_Stationary_matrix_6_1,
  input  [15:0] io_Stationary_matrix_6_2,
  input  [15:0] io_Stationary_matrix_6_3,
  input  [15:0] io_Stationary_matrix_6_4,
  input  [15:0] io_Stationary_matrix_6_5,
  input  [15:0] io_Stationary_matrix_6_6,
  input  [15:0] io_Stationary_matrix_6_7,
  input  [15:0] io_Stationary_matrix_7_0,
  input  [15:0] io_Stationary_matrix_7_1,
  input  [15:0] io_Stationary_matrix_7_2,
  input  [15:0] io_Stationary_matrix_7_3,
  input  [15:0] io_Stationary_matrix_7_4,
  input  [15:0] io_Stationary_matrix_7_5,
  input  [15:0] io_Stationary_matrix_7_6,
  input  [15:0] io_Stationary_matrix_7_7,
  input  [15:0] io_Streaming_matrix_0,
  input  [15:0] io_Streaming_matrix_1,
  input  [15:0] io_Streaming_matrix_2,
  input  [15:0] io_Streaming_matrix_3,
  input  [15:0] io_Streaming_matrix_4,
  input  [15:0] io_Streaming_matrix_5,
  input  [15:0] io_Streaming_matrix_6,
  input  [15:0] io_Streaming_matrix_7,
  output [15:0] io_counterMatrix1_bits_0_0,
  output [15:0] io_counterMatrix1_bits_0_1,
  output [15:0] io_counterMatrix1_bits_0_2,
  output [15:0] io_counterMatrix1_bits_0_3,
  output [15:0] io_counterMatrix1_bits_0_4,
  output [15:0] io_counterMatrix1_bits_0_5,
  output [15:0] io_counterMatrix1_bits_0_6,
  output [15:0] io_counterMatrix1_bits_0_7,
  output [15:0] io_counterMatrix1_bits_1_0,
  output [15:0] io_counterMatrix1_bits_1_1,
  output [15:0] io_counterMatrix1_bits_1_2,
  output [15:0] io_counterMatrix1_bits_1_3,
  output [15:0] io_counterMatrix1_bits_1_4,
  output [15:0] io_counterMatrix1_bits_1_5,
  output [15:0] io_counterMatrix1_bits_1_6,
  output [15:0] io_counterMatrix1_bits_1_7,
  output [15:0] io_counterMatrix1_bits_2_0,
  output [15:0] io_counterMatrix1_bits_2_1,
  output [15:0] io_counterMatrix1_bits_2_2,
  output [15:0] io_counterMatrix1_bits_2_3,
  output [15:0] io_counterMatrix1_bits_2_4,
  output [15:0] io_counterMatrix1_bits_2_5,
  output [15:0] io_counterMatrix1_bits_2_6,
  output [15:0] io_counterMatrix1_bits_2_7,
  output [15:0] io_counterMatrix1_bits_3_0,
  output [15:0] io_counterMatrix1_bits_3_1,
  output [15:0] io_counterMatrix1_bits_3_2,
  output [15:0] io_counterMatrix1_bits_3_3,
  output [15:0] io_counterMatrix1_bits_3_4,
  output [15:0] io_counterMatrix1_bits_3_5,
  output [15:0] io_counterMatrix1_bits_3_6,
  output [15:0] io_counterMatrix1_bits_3_7,
  output [15:0] io_counterMatrix1_bits_4_0,
  output [15:0] io_counterMatrix1_bits_4_1,
  output [15:0] io_counterMatrix1_bits_4_2,
  output [15:0] io_counterMatrix1_bits_4_3,
  output [15:0] io_counterMatrix1_bits_4_4,
  output [15:0] io_counterMatrix1_bits_4_5,
  output [15:0] io_counterMatrix1_bits_4_6,
  output [15:0] io_counterMatrix1_bits_4_7,
  output [15:0] io_counterMatrix1_bits_5_0,
  output [15:0] io_counterMatrix1_bits_5_1,
  output [15:0] io_counterMatrix1_bits_5_2,
  output [15:0] io_counterMatrix1_bits_5_3,
  output [15:0] io_counterMatrix1_bits_5_4,
  output [15:0] io_counterMatrix1_bits_5_5,
  output [15:0] io_counterMatrix1_bits_5_6,
  output [15:0] io_counterMatrix1_bits_5_7,
  output [15:0] io_counterMatrix1_bits_6_0,
  output [15:0] io_counterMatrix1_bits_6_1,
  output [15:0] io_counterMatrix1_bits_6_2,
  output [15:0] io_counterMatrix1_bits_6_3,
  output [15:0] io_counterMatrix1_bits_6_4,
  output [15:0] io_counterMatrix1_bits_6_5,
  output [15:0] io_counterMatrix1_bits_6_6,
  output [15:0] io_counterMatrix1_bits_6_7,
  output [15:0] io_counterMatrix1_bits_7_0,
  output [15:0] io_counterMatrix1_bits_7_1,
  output [15:0] io_counterMatrix1_bits_7_2,
  output [15:0] io_counterMatrix1_bits_7_3,
  output [15:0] io_counterMatrix1_bits_7_4,
  output [15:0] io_counterMatrix1_bits_7_5,
  output [15:0] io_counterMatrix1_bits_7_6,
  output [15:0] io_counterMatrix1_bits_7_7,
  output [15:0] io_counterMatrix2_bits_0,
  output [15:0] io_counterMatrix2_bits_1,
  output [15:0] io_counterMatrix2_bits_2,
  output [15:0] io_counterMatrix2_bits_3,
  output [15:0] io_counterMatrix2_bits_4,
  output [15:0] io_counterMatrix2_bits_5,
  output [15:0] io_counterMatrix2_bits_6,
  output [15:0] io_counterMatrix2_bits_7,
  output        io_valid,
  input         io_start
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
`endif // RANDOMIZE_REG_INIT
  reg [15:0] prevStationary_matrix_0_0; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_0_1; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_0_2; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_0_3; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_0_4; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_0_5; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_0_6; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_0_7; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_1_0; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_1_1; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_1_2; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_1_3; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_1_4; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_1_5; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_1_6; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_1_7; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_2_0; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_2_1; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_2_2; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_2_3; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_2_4; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_2_5; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_2_6; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_2_7; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_3_0; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_3_1; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_3_2; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_3_3; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_3_4; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_3_5; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_3_6; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_3_7; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_4_0; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_4_1; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_4_2; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_4_3; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_4_4; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_4_5; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_4_6; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_4_7; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_5_0; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_5_1; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_5_2; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_5_3; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_5_4; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_5_5; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_5_6; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_5_7; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_6_0; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_6_1; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_6_2; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_6_3; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_6_4; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_6_5; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_6_6; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_6_7; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_7_0; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_7_1; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_7_2; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_7_3; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_7_4; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_7_5; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_7_6; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_7_7; // @[SourceDestination.scala 15:40]
  reg  matricesAreEqual; // @[SourceDestination.scala 16:31]
  reg [15:0] counterRegs1_0_0; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_0_1; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_0_2; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_0_3; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_0_4; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_0_5; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_0_6; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_0_7; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_1_0; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_1_1; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_1_2; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_1_3; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_1_4; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_1_5; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_1_6; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_1_7; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_2_0; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_2_1; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_2_2; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_2_3; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_2_4; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_2_5; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_2_6; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_2_7; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_3_0; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_3_1; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_3_2; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_3_3; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_3_4; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_3_5; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_3_6; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_3_7; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_4_0; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_4_1; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_4_2; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_4_3; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_4_4; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_4_5; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_4_6; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_4_7; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_5_0; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_5_1; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_5_2; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_5_3; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_5_4; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_5_5; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_5_6; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_5_7; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_6_0; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_6_1; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_6_2; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_6_3; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_6_4; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_6_5; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_6_6; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_6_7; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_7_0; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_7_1; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_7_2; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_7_3; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_7_4; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_7_5; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_7_6; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_7_7; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs2_0; // @[SourceDestination.scala 18:31]
  reg [15:0] counterRegs2_1; // @[SourceDestination.scala 18:31]
  reg [15:0] counterRegs2_2; // @[SourceDestination.scala 18:31]
  reg [15:0] counterRegs2_3; // @[SourceDestination.scala 18:31]
  reg [15:0] counterRegs2_4; // @[SourceDestination.scala 18:31]
  reg [15:0] counterRegs2_5; // @[SourceDestination.scala 18:31]
  reg [15:0] counterRegs2_6; // @[SourceDestination.scala 18:31]
  reg [15:0] counterRegs2_7; // @[SourceDestination.scala 18:31]
  reg [31:0] i; // @[SourceDestination.scala 20:20]
  reg [31:0] j; // @[SourceDestination.scala 21:20]
  reg  jValid; // @[SourceDestination.scala 25:21]
  reg [31:0] k; // @[SourceDestination.scala 26:20]
  reg [31:0] counter1; // @[SourceDestination.scala 28:27]
  reg [31:0] counter2; // @[SourceDestination.scala 29:27]
  wire  _reg_i_T_2 = j == 32'h7 & i == 32'h7; // @[SourceDestination.scala 31:57]
  wire  _GEN_0 = io_Stationary_matrix_0_0 != prevStationary_matrix_0_0 ? 1'h0 : 1'h1; // @[SourceDestination.scala 36:22 40:74 41:28]
  wire  _GEN_1 = io_Stationary_matrix_0_1 != prevStationary_matrix_0_1 ? 1'h0 : _GEN_0; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_2 = io_Stationary_matrix_0_2 != prevStationary_matrix_0_2 ? 1'h0 : _GEN_1; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_3 = io_Stationary_matrix_0_3 != prevStationary_matrix_0_3 ? 1'h0 : _GEN_2; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_4 = io_Stationary_matrix_0_4 != prevStationary_matrix_0_4 ? 1'h0 : _GEN_3; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_5 = io_Stationary_matrix_0_5 != prevStationary_matrix_0_5 ? 1'h0 : _GEN_4; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_6 = io_Stationary_matrix_0_6 != prevStationary_matrix_0_6 ? 1'h0 : _GEN_5; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_7 = io_Stationary_matrix_0_7 != prevStationary_matrix_0_7 ? 1'h0 : _GEN_6; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_8 = io_Stationary_matrix_1_0 != prevStationary_matrix_1_0 ? 1'h0 : _GEN_7; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_9 = io_Stationary_matrix_1_1 != prevStationary_matrix_1_1 ? 1'h0 : _GEN_8; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_10 = io_Stationary_matrix_1_2 != prevStationary_matrix_1_2 ? 1'h0 : _GEN_9; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_11 = io_Stationary_matrix_1_3 != prevStationary_matrix_1_3 ? 1'h0 : _GEN_10; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_12 = io_Stationary_matrix_1_4 != prevStationary_matrix_1_4 ? 1'h0 : _GEN_11; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_13 = io_Stationary_matrix_1_5 != prevStationary_matrix_1_5 ? 1'h0 : _GEN_12; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_14 = io_Stationary_matrix_1_6 != prevStationary_matrix_1_6 ? 1'h0 : _GEN_13; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_15 = io_Stationary_matrix_1_7 != prevStationary_matrix_1_7 ? 1'h0 : _GEN_14; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_16 = io_Stationary_matrix_2_0 != prevStationary_matrix_2_0 ? 1'h0 : _GEN_15; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_17 = io_Stationary_matrix_2_1 != prevStationary_matrix_2_1 ? 1'h0 : _GEN_16; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_18 = io_Stationary_matrix_2_2 != prevStationary_matrix_2_2 ? 1'h0 : _GEN_17; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_19 = io_Stationary_matrix_2_3 != prevStationary_matrix_2_3 ? 1'h0 : _GEN_18; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_20 = io_Stationary_matrix_2_4 != prevStationary_matrix_2_4 ? 1'h0 : _GEN_19; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_21 = io_Stationary_matrix_2_5 != prevStationary_matrix_2_5 ? 1'h0 : _GEN_20; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_22 = io_Stationary_matrix_2_6 != prevStationary_matrix_2_6 ? 1'h0 : _GEN_21; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_23 = io_Stationary_matrix_2_7 != prevStationary_matrix_2_7 ? 1'h0 : _GEN_22; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_24 = io_Stationary_matrix_3_0 != prevStationary_matrix_3_0 ? 1'h0 : _GEN_23; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_25 = io_Stationary_matrix_3_1 != prevStationary_matrix_3_1 ? 1'h0 : _GEN_24; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_26 = io_Stationary_matrix_3_2 != prevStationary_matrix_3_2 ? 1'h0 : _GEN_25; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_27 = io_Stationary_matrix_3_3 != prevStationary_matrix_3_3 ? 1'h0 : _GEN_26; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_28 = io_Stationary_matrix_3_4 != prevStationary_matrix_3_4 ? 1'h0 : _GEN_27; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_29 = io_Stationary_matrix_3_5 != prevStationary_matrix_3_5 ? 1'h0 : _GEN_28; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_30 = io_Stationary_matrix_3_6 != prevStationary_matrix_3_6 ? 1'h0 : _GEN_29; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_31 = io_Stationary_matrix_3_7 != prevStationary_matrix_3_7 ? 1'h0 : _GEN_30; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_32 = io_Stationary_matrix_4_0 != prevStationary_matrix_4_0 ? 1'h0 : _GEN_31; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_33 = io_Stationary_matrix_4_1 != prevStationary_matrix_4_1 ? 1'h0 : _GEN_32; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_34 = io_Stationary_matrix_4_2 != prevStationary_matrix_4_2 ? 1'h0 : _GEN_33; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_35 = io_Stationary_matrix_4_3 != prevStationary_matrix_4_3 ? 1'h0 : _GEN_34; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_36 = io_Stationary_matrix_4_4 != prevStationary_matrix_4_4 ? 1'h0 : _GEN_35; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_37 = io_Stationary_matrix_4_5 != prevStationary_matrix_4_5 ? 1'h0 : _GEN_36; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_38 = io_Stationary_matrix_4_6 != prevStationary_matrix_4_6 ? 1'h0 : _GEN_37; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_39 = io_Stationary_matrix_4_7 != prevStationary_matrix_4_7 ? 1'h0 : _GEN_38; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_40 = io_Stationary_matrix_5_0 != prevStationary_matrix_5_0 ? 1'h0 : _GEN_39; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_41 = io_Stationary_matrix_5_1 != prevStationary_matrix_5_1 ? 1'h0 : _GEN_40; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_42 = io_Stationary_matrix_5_2 != prevStationary_matrix_5_2 ? 1'h0 : _GEN_41; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_43 = io_Stationary_matrix_5_3 != prevStationary_matrix_5_3 ? 1'h0 : _GEN_42; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_44 = io_Stationary_matrix_5_4 != prevStationary_matrix_5_4 ? 1'h0 : _GEN_43; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_45 = io_Stationary_matrix_5_5 != prevStationary_matrix_5_5 ? 1'h0 : _GEN_44; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_46 = io_Stationary_matrix_5_6 != prevStationary_matrix_5_6 ? 1'h0 : _GEN_45; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_47 = io_Stationary_matrix_5_7 != prevStationary_matrix_5_7 ? 1'h0 : _GEN_46; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_48 = io_Stationary_matrix_6_0 != prevStationary_matrix_6_0 ? 1'h0 : _GEN_47; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_49 = io_Stationary_matrix_6_1 != prevStationary_matrix_6_1 ? 1'h0 : _GEN_48; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_50 = io_Stationary_matrix_6_2 != prevStationary_matrix_6_2 ? 1'h0 : _GEN_49; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_51 = io_Stationary_matrix_6_3 != prevStationary_matrix_6_3 ? 1'h0 : _GEN_50; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_52 = io_Stationary_matrix_6_4 != prevStationary_matrix_6_4 ? 1'h0 : _GEN_51; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_53 = io_Stationary_matrix_6_5 != prevStationary_matrix_6_5 ? 1'h0 : _GEN_52; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_54 = io_Stationary_matrix_6_6 != prevStationary_matrix_6_6 ? 1'h0 : _GEN_53; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_55 = io_Stationary_matrix_6_7 != prevStationary_matrix_6_7 ? 1'h0 : _GEN_54; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_56 = io_Stationary_matrix_7_0 != prevStationary_matrix_7_0 ? 1'h0 : _GEN_55; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_57 = io_Stationary_matrix_7_1 != prevStationary_matrix_7_1 ? 1'h0 : _GEN_56; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_58 = io_Stationary_matrix_7_2 != prevStationary_matrix_7_2 ? 1'h0 : _GEN_57; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_59 = io_Stationary_matrix_7_3 != prevStationary_matrix_7_3 ? 1'h0 : _GEN_58; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_60 = io_Stationary_matrix_7_4 != prevStationary_matrix_7_4 ? 1'h0 : _GEN_59; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_796 = 3'h0 == i[2:0]; // @[SourceDestination.scala 53:{38,38}]
  wire  _GEN_797 = 3'h1 == j[2:0]; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_65 = 3'h0 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_0_1 : io_Stationary_matrix_0_0; // @[SourceDestination.scala 53:{38,38}]
  wire  _GEN_799 = 3'h2 == j[2:0]; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_66 = 3'h0 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_0_2 : _GEN_65; // @[SourceDestination.scala 53:{38,38}]
  wire  _GEN_801 = 3'h3 == j[2:0]; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_67 = 3'h0 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_0_3 : _GEN_66; // @[SourceDestination.scala 53:{38,38}]
  wire  _GEN_803 = 3'h4 == j[2:0]; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_68 = 3'h0 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_0_4 : _GEN_67; // @[SourceDestination.scala 53:{38,38}]
  wire  _GEN_805 = 3'h5 == j[2:0]; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_69 = 3'h0 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_0_5 : _GEN_68; // @[SourceDestination.scala 53:{38,38}]
  wire  _GEN_807 = 3'h6 == j[2:0]; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_70 = 3'h0 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_0_6 : _GEN_69; // @[SourceDestination.scala 53:{38,38}]
  wire  _GEN_809 = 3'h7 == j[2:0]; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_71 = 3'h0 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_0_7 : _GEN_70; // @[SourceDestination.scala 53:{38,38}]
  wire  _GEN_810 = 3'h1 == i[2:0]; // @[SourceDestination.scala 53:{38,38}]
  wire  _GEN_811 = 3'h0 == j[2:0]; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_72 = 3'h1 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_1_0 : _GEN_71; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_73 = 3'h1 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_1_1 : _GEN_72; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_74 = 3'h1 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_1_2 : _GEN_73; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_75 = 3'h1 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_1_3 : _GEN_74; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_76 = 3'h1 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_1_4 : _GEN_75; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_77 = 3'h1 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_1_5 : _GEN_76; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_78 = 3'h1 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_1_6 : _GEN_77; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_79 = 3'h1 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_1_7 : _GEN_78; // @[SourceDestination.scala 53:{38,38}]
  wire  _GEN_826 = 3'h2 == i[2:0]; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_80 = 3'h2 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_2_0 : _GEN_79; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_81 = 3'h2 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_2_1 : _GEN_80; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_82 = 3'h2 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_2_2 : _GEN_81; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_83 = 3'h2 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_2_3 : _GEN_82; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_84 = 3'h2 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_2_4 : _GEN_83; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_85 = 3'h2 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_2_5 : _GEN_84; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_86 = 3'h2 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_2_6 : _GEN_85; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_87 = 3'h2 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_2_7 : _GEN_86; // @[SourceDestination.scala 53:{38,38}]
  wire  _GEN_842 = 3'h3 == i[2:0]; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_88 = 3'h3 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_3_0 : _GEN_87; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_89 = 3'h3 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_3_1 : _GEN_88; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_90 = 3'h3 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_3_2 : _GEN_89; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_91 = 3'h3 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_3_3 : _GEN_90; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_92 = 3'h3 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_3_4 : _GEN_91; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_93 = 3'h3 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_3_5 : _GEN_92; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_94 = 3'h3 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_3_6 : _GEN_93; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_95 = 3'h3 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_3_7 : _GEN_94; // @[SourceDestination.scala 53:{38,38}]
  wire  _GEN_858 = 3'h4 == i[2:0]; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_96 = 3'h4 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_4_0 : _GEN_95; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_97 = 3'h4 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_4_1 : _GEN_96; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_98 = 3'h4 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_4_2 : _GEN_97; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_99 = 3'h4 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_4_3 : _GEN_98; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_100 = 3'h4 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_4_4 : _GEN_99; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_101 = 3'h4 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_4_5 : _GEN_100; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_102 = 3'h4 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_4_6 : _GEN_101; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_103 = 3'h4 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_4_7 : _GEN_102; // @[SourceDestination.scala 53:{38,38}]
  wire  _GEN_874 = 3'h5 == i[2:0]; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_104 = 3'h5 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_5_0 : _GEN_103; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_105 = 3'h5 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_5_1 : _GEN_104; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_106 = 3'h5 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_5_2 : _GEN_105; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_107 = 3'h5 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_5_3 : _GEN_106; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_108 = 3'h5 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_5_4 : _GEN_107; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_109 = 3'h5 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_5_5 : _GEN_108; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_110 = 3'h5 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_5_6 : _GEN_109; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_111 = 3'h5 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_5_7 : _GEN_110; // @[SourceDestination.scala 53:{38,38}]
  wire  _GEN_890 = 3'h6 == i[2:0]; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_112 = 3'h6 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_6_0 : _GEN_111; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_113 = 3'h6 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_6_1 : _GEN_112; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_114 = 3'h6 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_6_2 : _GEN_113; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_115 = 3'h6 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_6_3 : _GEN_114; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_116 = 3'h6 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_6_4 : _GEN_115; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_117 = 3'h6 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_6_5 : _GEN_116; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_118 = 3'h6 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_6_6 : _GEN_117; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_119 = 3'h6 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_6_7 : _GEN_118; // @[SourceDestination.scala 53:{38,38}]
  wire  _GEN_906 = 3'h7 == i[2:0]; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_120 = 3'h7 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_7_0 : _GEN_119; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_121 = 3'h7 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_7_1 : _GEN_120; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_122 = 3'h7 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_7_2 : _GEN_121; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_123 = 3'h7 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_7_3 : _GEN_122; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_124 = 3'h7 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_7_4 : _GEN_123; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_125 = 3'h7 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_7_5 : _GEN_124; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_126 = 3'h7 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_7_6 : _GEN_125; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_127 = 3'h7 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_7_7 : _GEN_126; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_128 = _GEN_796 & _GEN_811 ? counter1[15:0] : counterRegs1_0_0; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_129 = _GEN_796 & _GEN_797 ? counter1[15:0] : counterRegs1_0_1; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_130 = _GEN_796 & _GEN_799 ? counter1[15:0] : counterRegs1_0_2; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_131 = _GEN_796 & _GEN_801 ? counter1[15:0] : counterRegs1_0_3; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_132 = _GEN_796 & _GEN_803 ? counter1[15:0] : counterRegs1_0_4; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_133 = _GEN_796 & _GEN_805 ? counter1[15:0] : counterRegs1_0_5; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_134 = _GEN_796 & _GEN_807 ? counter1[15:0] : counterRegs1_0_6; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_135 = _GEN_796 & _GEN_809 ? counter1[15:0] : counterRegs1_0_7; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_136 = _GEN_810 & _GEN_811 ? counter1[15:0] : counterRegs1_1_0; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_137 = _GEN_810 & _GEN_797 ? counter1[15:0] : counterRegs1_1_1; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_138 = _GEN_810 & _GEN_799 ? counter1[15:0] : counterRegs1_1_2; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_139 = _GEN_810 & _GEN_801 ? counter1[15:0] : counterRegs1_1_3; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_140 = _GEN_810 & _GEN_803 ? counter1[15:0] : counterRegs1_1_4; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_141 = _GEN_810 & _GEN_805 ? counter1[15:0] : counterRegs1_1_5; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_142 = _GEN_810 & _GEN_807 ? counter1[15:0] : counterRegs1_1_6; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_143 = _GEN_810 & _GEN_809 ? counter1[15:0] : counterRegs1_1_7; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_144 = _GEN_826 & _GEN_811 ? counter1[15:0] : counterRegs1_2_0; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_145 = _GEN_826 & _GEN_797 ? counter1[15:0] : counterRegs1_2_1; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_146 = _GEN_826 & _GEN_799 ? counter1[15:0] : counterRegs1_2_2; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_147 = _GEN_826 & _GEN_801 ? counter1[15:0] : counterRegs1_2_3; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_148 = _GEN_826 & _GEN_803 ? counter1[15:0] : counterRegs1_2_4; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_149 = _GEN_826 & _GEN_805 ? counter1[15:0] : counterRegs1_2_5; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_150 = _GEN_826 & _GEN_807 ? counter1[15:0] : counterRegs1_2_6; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_151 = _GEN_826 & _GEN_809 ? counter1[15:0] : counterRegs1_2_7; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_152 = _GEN_842 & _GEN_811 ? counter1[15:0] : counterRegs1_3_0; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_153 = _GEN_842 & _GEN_797 ? counter1[15:0] : counterRegs1_3_1; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_154 = _GEN_842 & _GEN_799 ? counter1[15:0] : counterRegs1_3_2; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_155 = _GEN_842 & _GEN_801 ? counter1[15:0] : counterRegs1_3_3; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_156 = _GEN_842 & _GEN_803 ? counter1[15:0] : counterRegs1_3_4; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_157 = _GEN_842 & _GEN_805 ? counter1[15:0] : counterRegs1_3_5; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_158 = _GEN_842 & _GEN_807 ? counter1[15:0] : counterRegs1_3_6; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_159 = _GEN_842 & _GEN_809 ? counter1[15:0] : counterRegs1_3_7; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_160 = _GEN_858 & _GEN_811 ? counter1[15:0] : counterRegs1_4_0; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_161 = _GEN_858 & _GEN_797 ? counter1[15:0] : counterRegs1_4_1; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_162 = _GEN_858 & _GEN_799 ? counter1[15:0] : counterRegs1_4_2; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_163 = _GEN_858 & _GEN_801 ? counter1[15:0] : counterRegs1_4_3; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_164 = _GEN_858 & _GEN_803 ? counter1[15:0] : counterRegs1_4_4; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_165 = _GEN_858 & _GEN_805 ? counter1[15:0] : counterRegs1_4_5; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_166 = _GEN_858 & _GEN_807 ? counter1[15:0] : counterRegs1_4_6; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_167 = _GEN_858 & _GEN_809 ? counter1[15:0] : counterRegs1_4_7; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_168 = _GEN_874 & _GEN_811 ? counter1[15:0] : counterRegs1_5_0; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_169 = _GEN_874 & _GEN_797 ? counter1[15:0] : counterRegs1_5_1; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_170 = _GEN_874 & _GEN_799 ? counter1[15:0] : counterRegs1_5_2; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_171 = _GEN_874 & _GEN_801 ? counter1[15:0] : counterRegs1_5_3; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_172 = _GEN_874 & _GEN_803 ? counter1[15:0] : counterRegs1_5_4; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_173 = _GEN_874 & _GEN_805 ? counter1[15:0] : counterRegs1_5_5; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_174 = _GEN_874 & _GEN_807 ? counter1[15:0] : counterRegs1_5_6; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_175 = _GEN_874 & _GEN_809 ? counter1[15:0] : counterRegs1_5_7; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_176 = _GEN_890 & _GEN_811 ? counter1[15:0] : counterRegs1_6_0; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_177 = _GEN_890 & _GEN_797 ? counter1[15:0] : counterRegs1_6_1; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_178 = _GEN_890 & _GEN_799 ? counter1[15:0] : counterRegs1_6_2; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_179 = _GEN_890 & _GEN_801 ? counter1[15:0] : counterRegs1_6_3; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_180 = _GEN_890 & _GEN_803 ? counter1[15:0] : counterRegs1_6_4; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_181 = _GEN_890 & _GEN_805 ? counter1[15:0] : counterRegs1_6_5; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_182 = _GEN_890 & _GEN_807 ? counter1[15:0] : counterRegs1_6_6; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_183 = _GEN_890 & _GEN_809 ? counter1[15:0] : counterRegs1_6_7; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_184 = _GEN_906 & _GEN_811 ? counter1[15:0] : counterRegs1_7_0; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_185 = _GEN_906 & _GEN_797 ? counter1[15:0] : counterRegs1_7_1; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_186 = _GEN_906 & _GEN_799 ? counter1[15:0] : counterRegs1_7_2; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_187 = _GEN_906 & _GEN_801 ? counter1[15:0] : counterRegs1_7_3; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_188 = _GEN_906 & _GEN_803 ? counter1[15:0] : counterRegs1_7_4; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_189 = _GEN_906 & _GEN_805 ? counter1[15:0] : counterRegs1_7_5; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_190 = _GEN_906 & _GEN_807 ? counter1[15:0] : counterRegs1_7_6; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_191 = _GEN_906 & _GEN_809 ? counter1[15:0] : counterRegs1_7_7; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [31:0] _counter1_T_1 = counter1 + 32'h1; // @[SourceDestination.scala 57:32]
  wire [31:0] _GEN_192 = ~_reg_i_T_2 ? _counter1_T_1 : counter1; // @[SourceDestination.scala 56:83 57:20 28:27]
  wire [15:0] _GEN_193 = _GEN_796 & _GEN_811 ? 16'h1 : counterRegs1_0_0; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_194 = _GEN_796 & _GEN_797 ? 16'h1 : counterRegs1_0_1; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_195 = _GEN_796 & _GEN_799 ? 16'h1 : counterRegs1_0_2; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_196 = _GEN_796 & _GEN_801 ? 16'h1 : counterRegs1_0_3; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_197 = _GEN_796 & _GEN_803 ? 16'h1 : counterRegs1_0_4; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_198 = _GEN_796 & _GEN_805 ? 16'h1 : counterRegs1_0_5; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_199 = _GEN_796 & _GEN_807 ? 16'h1 : counterRegs1_0_6; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_200 = _GEN_796 & _GEN_809 ? 16'h1 : counterRegs1_0_7; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_201 = _GEN_810 & _GEN_811 ? 16'h1 : counterRegs1_1_0; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_202 = _GEN_810 & _GEN_797 ? 16'h1 : counterRegs1_1_1; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_203 = _GEN_810 & _GEN_799 ? 16'h1 : counterRegs1_1_2; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_204 = _GEN_810 & _GEN_801 ? 16'h1 : counterRegs1_1_3; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_205 = _GEN_810 & _GEN_803 ? 16'h1 : counterRegs1_1_4; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_206 = _GEN_810 & _GEN_805 ? 16'h1 : counterRegs1_1_5; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_207 = _GEN_810 & _GEN_807 ? 16'h1 : counterRegs1_1_6; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_208 = _GEN_810 & _GEN_809 ? 16'h1 : counterRegs1_1_7; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_209 = _GEN_826 & _GEN_811 ? 16'h1 : counterRegs1_2_0; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_210 = _GEN_826 & _GEN_797 ? 16'h1 : counterRegs1_2_1; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_211 = _GEN_826 & _GEN_799 ? 16'h1 : counterRegs1_2_2; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_212 = _GEN_826 & _GEN_801 ? 16'h1 : counterRegs1_2_3; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_213 = _GEN_826 & _GEN_803 ? 16'h1 : counterRegs1_2_4; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_214 = _GEN_826 & _GEN_805 ? 16'h1 : counterRegs1_2_5; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_215 = _GEN_826 & _GEN_807 ? 16'h1 : counterRegs1_2_6; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_216 = _GEN_826 & _GEN_809 ? 16'h1 : counterRegs1_2_7; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_217 = _GEN_842 & _GEN_811 ? 16'h1 : counterRegs1_3_0; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_218 = _GEN_842 & _GEN_797 ? 16'h1 : counterRegs1_3_1; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_219 = _GEN_842 & _GEN_799 ? 16'h1 : counterRegs1_3_2; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_220 = _GEN_842 & _GEN_801 ? 16'h1 : counterRegs1_3_3; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_221 = _GEN_842 & _GEN_803 ? 16'h1 : counterRegs1_3_4; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_222 = _GEN_842 & _GEN_805 ? 16'h1 : counterRegs1_3_5; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_223 = _GEN_842 & _GEN_807 ? 16'h1 : counterRegs1_3_6; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_224 = _GEN_842 & _GEN_809 ? 16'h1 : counterRegs1_3_7; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_225 = _GEN_858 & _GEN_811 ? 16'h1 : counterRegs1_4_0; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_226 = _GEN_858 & _GEN_797 ? 16'h1 : counterRegs1_4_1; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_227 = _GEN_858 & _GEN_799 ? 16'h1 : counterRegs1_4_2; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_228 = _GEN_858 & _GEN_801 ? 16'h1 : counterRegs1_4_3; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_229 = _GEN_858 & _GEN_803 ? 16'h1 : counterRegs1_4_4; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_230 = _GEN_858 & _GEN_805 ? 16'h1 : counterRegs1_4_5; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_231 = _GEN_858 & _GEN_807 ? 16'h1 : counterRegs1_4_6; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_232 = _GEN_858 & _GEN_809 ? 16'h1 : counterRegs1_4_7; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_233 = _GEN_874 & _GEN_811 ? 16'h1 : counterRegs1_5_0; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_234 = _GEN_874 & _GEN_797 ? 16'h1 : counterRegs1_5_1; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_235 = _GEN_874 & _GEN_799 ? 16'h1 : counterRegs1_5_2; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_236 = _GEN_874 & _GEN_801 ? 16'h1 : counterRegs1_5_3; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_237 = _GEN_874 & _GEN_803 ? 16'h1 : counterRegs1_5_4; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_238 = _GEN_874 & _GEN_805 ? 16'h1 : counterRegs1_5_5; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_239 = _GEN_874 & _GEN_807 ? 16'h1 : counterRegs1_5_6; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_240 = _GEN_874 & _GEN_809 ? 16'h1 : counterRegs1_5_7; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_241 = _GEN_890 & _GEN_811 ? 16'h1 : counterRegs1_6_0; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_242 = _GEN_890 & _GEN_797 ? 16'h1 : counterRegs1_6_1; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_243 = _GEN_890 & _GEN_799 ? 16'h1 : counterRegs1_6_2; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_244 = _GEN_890 & _GEN_801 ? 16'h1 : counterRegs1_6_3; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_245 = _GEN_890 & _GEN_803 ? 16'h1 : counterRegs1_6_4; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_246 = _GEN_890 & _GEN_805 ? 16'h1 : counterRegs1_6_5; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_247 = _GEN_890 & _GEN_807 ? 16'h1 : counterRegs1_6_6; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_248 = _GEN_890 & _GEN_809 ? 16'h1 : counterRegs1_6_7; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_249 = _GEN_906 & _GEN_811 ? 16'h1 : counterRegs1_7_0; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_250 = _GEN_906 & _GEN_797 ? 16'h1 : counterRegs1_7_1; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_251 = _GEN_906 & _GEN_799 ? 16'h1 : counterRegs1_7_2; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_252 = _GEN_906 & _GEN_801 ? 16'h1 : counterRegs1_7_3; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_253 = _GEN_906 & _GEN_803 ? 16'h1 : counterRegs1_7_4; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_254 = _GEN_906 & _GEN_805 ? 16'h1 : counterRegs1_7_5; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_255 = _GEN_906 & _GEN_807 ? 16'h1 : counterRegs1_7_6; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_256 = _GEN_906 & _GEN_809 ? 16'h1 : counterRegs1_7_7; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_257 = counter1 < 32'h5 ? _GEN_128 : _GEN_193; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_258 = counter1 < 32'h5 ? _GEN_129 : _GEN_194; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_259 = counter1 < 32'h5 ? _GEN_130 : _GEN_195; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_260 = counter1 < 32'h5 ? _GEN_131 : _GEN_196; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_261 = counter1 < 32'h5 ? _GEN_132 : _GEN_197; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_262 = counter1 < 32'h5 ? _GEN_133 : _GEN_198; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_263 = counter1 < 32'h5 ? _GEN_134 : _GEN_199; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_264 = counter1 < 32'h5 ? _GEN_135 : _GEN_200; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_265 = counter1 < 32'h5 ? _GEN_136 : _GEN_201; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_266 = counter1 < 32'h5 ? _GEN_137 : _GEN_202; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_267 = counter1 < 32'h5 ? _GEN_138 : _GEN_203; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_268 = counter1 < 32'h5 ? _GEN_139 : _GEN_204; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_269 = counter1 < 32'h5 ? _GEN_140 : _GEN_205; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_270 = counter1 < 32'h5 ? _GEN_141 : _GEN_206; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_271 = counter1 < 32'h5 ? _GEN_142 : _GEN_207; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_272 = counter1 < 32'h5 ? _GEN_143 : _GEN_208; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_273 = counter1 < 32'h5 ? _GEN_144 : _GEN_209; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_274 = counter1 < 32'h5 ? _GEN_145 : _GEN_210; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_275 = counter1 < 32'h5 ? _GEN_146 : _GEN_211; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_276 = counter1 < 32'h5 ? _GEN_147 : _GEN_212; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_277 = counter1 < 32'h5 ? _GEN_148 : _GEN_213; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_278 = counter1 < 32'h5 ? _GEN_149 : _GEN_214; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_279 = counter1 < 32'h5 ? _GEN_150 : _GEN_215; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_280 = counter1 < 32'h5 ? _GEN_151 : _GEN_216; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_281 = counter1 < 32'h5 ? _GEN_152 : _GEN_217; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_282 = counter1 < 32'h5 ? _GEN_153 : _GEN_218; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_283 = counter1 < 32'h5 ? _GEN_154 : _GEN_219; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_284 = counter1 < 32'h5 ? _GEN_155 : _GEN_220; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_285 = counter1 < 32'h5 ? _GEN_156 : _GEN_221; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_286 = counter1 < 32'h5 ? _GEN_157 : _GEN_222; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_287 = counter1 < 32'h5 ? _GEN_158 : _GEN_223; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_288 = counter1 < 32'h5 ? _GEN_159 : _GEN_224; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_289 = counter1 < 32'h5 ? _GEN_160 : _GEN_225; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_290 = counter1 < 32'h5 ? _GEN_161 : _GEN_226; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_291 = counter1 < 32'h5 ? _GEN_162 : _GEN_227; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_292 = counter1 < 32'h5 ? _GEN_163 : _GEN_228; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_293 = counter1 < 32'h5 ? _GEN_164 : _GEN_229; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_294 = counter1 < 32'h5 ? _GEN_165 : _GEN_230; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_295 = counter1 < 32'h5 ? _GEN_166 : _GEN_231; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_296 = counter1 < 32'h5 ? _GEN_167 : _GEN_232; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_297 = counter1 < 32'h5 ? _GEN_168 : _GEN_233; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_298 = counter1 < 32'h5 ? _GEN_169 : _GEN_234; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_299 = counter1 < 32'h5 ? _GEN_170 : _GEN_235; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_300 = counter1 < 32'h5 ? _GEN_171 : _GEN_236; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_301 = counter1 < 32'h5 ? _GEN_172 : _GEN_237; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_302 = counter1 < 32'h5 ? _GEN_173 : _GEN_238; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_303 = counter1 < 32'h5 ? _GEN_174 : _GEN_239; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_304 = counter1 < 32'h5 ? _GEN_175 : _GEN_240; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_305 = counter1 < 32'h5 ? _GEN_176 : _GEN_241; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_306 = counter1 < 32'h5 ? _GEN_177 : _GEN_242; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_307 = counter1 < 32'h5 ? _GEN_178 : _GEN_243; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_308 = counter1 < 32'h5 ? _GEN_179 : _GEN_244; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_309 = counter1 < 32'h5 ? _GEN_180 : _GEN_245; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_310 = counter1 < 32'h5 ? _GEN_181 : _GEN_246; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_311 = counter1 < 32'h5 ? _GEN_182 : _GEN_247; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_312 = counter1 < 32'h5 ? _GEN_183 : _GEN_248; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_313 = counter1 < 32'h5 ? _GEN_184 : _GEN_249; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_314 = counter1 < 32'h5 ? _GEN_185 : _GEN_250; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_315 = counter1 < 32'h5 ? _GEN_186 : _GEN_251; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_316 = counter1 < 32'h5 ? _GEN_187 : _GEN_252; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_317 = counter1 < 32'h5 ? _GEN_188 : _GEN_253; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_318 = counter1 < 32'h5 ? _GEN_189 : _GEN_254; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_319 = counter1 < 32'h5 ? _GEN_190 : _GEN_255; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_320 = counter1 < 32'h5 ? _GEN_191 : _GEN_256; // @[SourceDestination.scala 54:48]
  wire [31:0] _GEN_321 = counter1 < 32'h5 ? _GEN_192 : 32'h2; // @[SourceDestination.scala 54:48 61:18]
  wire [15:0] _GEN_322 = _GEN_796 & _GEN_811 ? 16'h0 : counterRegs1_0_0; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_323 = _GEN_796 & _GEN_797 ? 16'h0 : counterRegs1_0_1; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_324 = _GEN_796 & _GEN_799 ? 16'h0 : counterRegs1_0_2; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_325 = _GEN_796 & _GEN_801 ? 16'h0 : counterRegs1_0_3; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_326 = _GEN_796 & _GEN_803 ? 16'h0 : counterRegs1_0_4; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_327 = _GEN_796 & _GEN_805 ? 16'h0 : counterRegs1_0_5; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_328 = _GEN_796 & _GEN_807 ? 16'h0 : counterRegs1_0_6; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_329 = _GEN_796 & _GEN_809 ? 16'h0 : counterRegs1_0_7; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_330 = _GEN_810 & _GEN_811 ? 16'h0 : counterRegs1_1_0; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_331 = _GEN_810 & _GEN_797 ? 16'h0 : counterRegs1_1_1; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_332 = _GEN_810 & _GEN_799 ? 16'h0 : counterRegs1_1_2; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_333 = _GEN_810 & _GEN_801 ? 16'h0 : counterRegs1_1_3; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_334 = _GEN_810 & _GEN_803 ? 16'h0 : counterRegs1_1_4; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_335 = _GEN_810 & _GEN_805 ? 16'h0 : counterRegs1_1_5; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_336 = _GEN_810 & _GEN_807 ? 16'h0 : counterRegs1_1_6; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_337 = _GEN_810 & _GEN_809 ? 16'h0 : counterRegs1_1_7; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_338 = _GEN_826 & _GEN_811 ? 16'h0 : counterRegs1_2_0; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_339 = _GEN_826 & _GEN_797 ? 16'h0 : counterRegs1_2_1; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_340 = _GEN_826 & _GEN_799 ? 16'h0 : counterRegs1_2_2; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_341 = _GEN_826 & _GEN_801 ? 16'h0 : counterRegs1_2_3; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_342 = _GEN_826 & _GEN_803 ? 16'h0 : counterRegs1_2_4; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_343 = _GEN_826 & _GEN_805 ? 16'h0 : counterRegs1_2_5; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_344 = _GEN_826 & _GEN_807 ? 16'h0 : counterRegs1_2_6; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_345 = _GEN_826 & _GEN_809 ? 16'h0 : counterRegs1_2_7; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_346 = _GEN_842 & _GEN_811 ? 16'h0 : counterRegs1_3_0; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_347 = _GEN_842 & _GEN_797 ? 16'h0 : counterRegs1_3_1; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_348 = _GEN_842 & _GEN_799 ? 16'h0 : counterRegs1_3_2; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_349 = _GEN_842 & _GEN_801 ? 16'h0 : counterRegs1_3_3; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_350 = _GEN_842 & _GEN_803 ? 16'h0 : counterRegs1_3_4; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_351 = _GEN_842 & _GEN_805 ? 16'h0 : counterRegs1_3_5; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_352 = _GEN_842 & _GEN_807 ? 16'h0 : counterRegs1_3_6; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_353 = _GEN_842 & _GEN_809 ? 16'h0 : counterRegs1_3_7; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_354 = _GEN_858 & _GEN_811 ? 16'h0 : counterRegs1_4_0; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_355 = _GEN_858 & _GEN_797 ? 16'h0 : counterRegs1_4_1; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_356 = _GEN_858 & _GEN_799 ? 16'h0 : counterRegs1_4_2; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_357 = _GEN_858 & _GEN_801 ? 16'h0 : counterRegs1_4_3; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_358 = _GEN_858 & _GEN_803 ? 16'h0 : counterRegs1_4_4; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_359 = _GEN_858 & _GEN_805 ? 16'h0 : counterRegs1_4_5; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_360 = _GEN_858 & _GEN_807 ? 16'h0 : counterRegs1_4_6; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_361 = _GEN_858 & _GEN_809 ? 16'h0 : counterRegs1_4_7; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_362 = _GEN_874 & _GEN_811 ? 16'h0 : counterRegs1_5_0; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_363 = _GEN_874 & _GEN_797 ? 16'h0 : counterRegs1_5_1; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_364 = _GEN_874 & _GEN_799 ? 16'h0 : counterRegs1_5_2; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_365 = _GEN_874 & _GEN_801 ? 16'h0 : counterRegs1_5_3; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_366 = _GEN_874 & _GEN_803 ? 16'h0 : counterRegs1_5_4; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_367 = _GEN_874 & _GEN_805 ? 16'h0 : counterRegs1_5_5; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_368 = _GEN_874 & _GEN_807 ? 16'h0 : counterRegs1_5_6; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_369 = _GEN_874 & _GEN_809 ? 16'h0 : counterRegs1_5_7; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_370 = _GEN_890 & _GEN_811 ? 16'h0 : counterRegs1_6_0; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_371 = _GEN_890 & _GEN_797 ? 16'h0 : counterRegs1_6_1; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_372 = _GEN_890 & _GEN_799 ? 16'h0 : counterRegs1_6_2; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_373 = _GEN_890 & _GEN_801 ? 16'h0 : counterRegs1_6_3; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_374 = _GEN_890 & _GEN_803 ? 16'h0 : counterRegs1_6_4; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_375 = _GEN_890 & _GEN_805 ? 16'h0 : counterRegs1_6_5; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_376 = _GEN_890 & _GEN_807 ? 16'h0 : counterRegs1_6_6; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_377 = _GEN_890 & _GEN_809 ? 16'h0 : counterRegs1_6_7; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_378 = _GEN_906 & _GEN_811 ? 16'h0 : counterRegs1_7_0; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_379 = _GEN_906 & _GEN_797 ? 16'h0 : counterRegs1_7_1; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_380 = _GEN_906 & _GEN_799 ? 16'h0 : counterRegs1_7_2; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_381 = _GEN_906 & _GEN_801 ? 16'h0 : counterRegs1_7_3; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_382 = _GEN_906 & _GEN_803 ? 16'h0 : counterRegs1_7_4; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_383 = _GEN_906 & _GEN_805 ? 16'h0 : counterRegs1_7_5; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_384 = _GEN_906 & _GEN_807 ? 16'h0 : counterRegs1_7_6; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_385 = _GEN_906 & _GEN_809 ? 16'h0 : counterRegs1_7_7; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_386 = _GEN_127 != 16'h0 ? _GEN_257 : _GEN_322; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_387 = _GEN_127 != 16'h0 ? _GEN_258 : _GEN_323; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_388 = _GEN_127 != 16'h0 ? _GEN_259 : _GEN_324; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_389 = _GEN_127 != 16'h0 ? _GEN_260 : _GEN_325; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_390 = _GEN_127 != 16'h0 ? _GEN_261 : _GEN_326; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_391 = _GEN_127 != 16'h0 ? _GEN_262 : _GEN_327; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_392 = _GEN_127 != 16'h0 ? _GEN_263 : _GEN_328; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_393 = _GEN_127 != 16'h0 ? _GEN_264 : _GEN_329; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_394 = _GEN_127 != 16'h0 ? _GEN_265 : _GEN_330; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_395 = _GEN_127 != 16'h0 ? _GEN_266 : _GEN_331; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_396 = _GEN_127 != 16'h0 ? _GEN_267 : _GEN_332; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_397 = _GEN_127 != 16'h0 ? _GEN_268 : _GEN_333; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_398 = _GEN_127 != 16'h0 ? _GEN_269 : _GEN_334; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_399 = _GEN_127 != 16'h0 ? _GEN_270 : _GEN_335; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_400 = _GEN_127 != 16'h0 ? _GEN_271 : _GEN_336; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_401 = _GEN_127 != 16'h0 ? _GEN_272 : _GEN_337; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_402 = _GEN_127 != 16'h0 ? _GEN_273 : _GEN_338; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_403 = _GEN_127 != 16'h0 ? _GEN_274 : _GEN_339; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_404 = _GEN_127 != 16'h0 ? _GEN_275 : _GEN_340; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_405 = _GEN_127 != 16'h0 ? _GEN_276 : _GEN_341; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_406 = _GEN_127 != 16'h0 ? _GEN_277 : _GEN_342; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_407 = _GEN_127 != 16'h0 ? _GEN_278 : _GEN_343; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_408 = _GEN_127 != 16'h0 ? _GEN_279 : _GEN_344; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_409 = _GEN_127 != 16'h0 ? _GEN_280 : _GEN_345; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_410 = _GEN_127 != 16'h0 ? _GEN_281 : _GEN_346; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_411 = _GEN_127 != 16'h0 ? _GEN_282 : _GEN_347; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_412 = _GEN_127 != 16'h0 ? _GEN_283 : _GEN_348; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_413 = _GEN_127 != 16'h0 ? _GEN_284 : _GEN_349; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_414 = _GEN_127 != 16'h0 ? _GEN_285 : _GEN_350; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_415 = _GEN_127 != 16'h0 ? _GEN_286 : _GEN_351; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_416 = _GEN_127 != 16'h0 ? _GEN_287 : _GEN_352; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_417 = _GEN_127 != 16'h0 ? _GEN_288 : _GEN_353; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_418 = _GEN_127 != 16'h0 ? _GEN_289 : _GEN_354; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_419 = _GEN_127 != 16'h0 ? _GEN_290 : _GEN_355; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_420 = _GEN_127 != 16'h0 ? _GEN_291 : _GEN_356; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_421 = _GEN_127 != 16'h0 ? _GEN_292 : _GEN_357; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_422 = _GEN_127 != 16'h0 ? _GEN_293 : _GEN_358; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_423 = _GEN_127 != 16'h0 ? _GEN_294 : _GEN_359; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_424 = _GEN_127 != 16'h0 ? _GEN_295 : _GEN_360; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_425 = _GEN_127 != 16'h0 ? _GEN_296 : _GEN_361; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_426 = _GEN_127 != 16'h0 ? _GEN_297 : _GEN_362; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_427 = _GEN_127 != 16'h0 ? _GEN_298 : _GEN_363; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_428 = _GEN_127 != 16'h0 ? _GEN_299 : _GEN_364; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_429 = _GEN_127 != 16'h0 ? _GEN_300 : _GEN_365; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_430 = _GEN_127 != 16'h0 ? _GEN_301 : _GEN_366; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_431 = _GEN_127 != 16'h0 ? _GEN_302 : _GEN_367; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_432 = _GEN_127 != 16'h0 ? _GEN_303 : _GEN_368; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_433 = _GEN_127 != 16'h0 ? _GEN_304 : _GEN_369; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_434 = _GEN_127 != 16'h0 ? _GEN_305 : _GEN_370; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_435 = _GEN_127 != 16'h0 ? _GEN_306 : _GEN_371; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_436 = _GEN_127 != 16'h0 ? _GEN_307 : _GEN_372; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_437 = _GEN_127 != 16'h0 ? _GEN_308 : _GEN_373; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_438 = _GEN_127 != 16'h0 ? _GEN_309 : _GEN_374; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_439 = _GEN_127 != 16'h0 ? _GEN_310 : _GEN_375; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_440 = _GEN_127 != 16'h0 ? _GEN_311 : _GEN_376; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_441 = _GEN_127 != 16'h0 ? _GEN_312 : _GEN_377; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_442 = _GEN_127 != 16'h0 ? _GEN_313 : _GEN_378; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_443 = _GEN_127 != 16'h0 ? _GEN_314 : _GEN_379; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_444 = _GEN_127 != 16'h0 ? _GEN_315 : _GEN_380; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_445 = _GEN_127 != 16'h0 ? _GEN_316 : _GEN_381; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_446 = _GEN_127 != 16'h0 ? _GEN_317 : _GEN_382; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_447 = _GEN_127 != 16'h0 ? _GEN_318 : _GEN_383; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_448 = _GEN_127 != 16'h0 ? _GEN_319 : _GEN_384; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_449 = _GEN_127 != 16'h0 ? _GEN_320 : _GEN_385; // @[SourceDestination.scala 53:47]
  wire [31:0] _GEN_450 = _GEN_127 != 16'h0 ? _GEN_321 : counter1; // @[SourceDestination.scala 28:27 53:47]
  wire [15:0] _GEN_452 = 3'h1 == k[2:0] ? io_Streaming_matrix_1 : io_Streaming_matrix_0; // @[SourceDestination.scala 67:{34,34}]
  wire [15:0] _GEN_453 = 3'h2 == k[2:0] ? io_Streaming_matrix_2 : _GEN_452; // @[SourceDestination.scala 67:{34,34}]
  wire [15:0] _GEN_454 = 3'h3 == k[2:0] ? io_Streaming_matrix_3 : _GEN_453; // @[SourceDestination.scala 67:{34,34}]
  wire [15:0] _GEN_455 = 3'h4 == k[2:0] ? io_Streaming_matrix_4 : _GEN_454; // @[SourceDestination.scala 67:{34,34}]
  wire [15:0] _GEN_456 = 3'h5 == k[2:0] ? io_Streaming_matrix_5 : _GEN_455; // @[SourceDestination.scala 67:{34,34}]
  wire [15:0] _GEN_457 = 3'h6 == k[2:0] ? io_Streaming_matrix_6 : _GEN_456; // @[SourceDestination.scala 67:{34,34}]
  wire [15:0] _GEN_458 = 3'h7 == k[2:0] ? io_Streaming_matrix_7 : _GEN_457; // @[SourceDestination.scala 67:{34,34}]
  wire [15:0] _GEN_459 = 3'h0 == k[2:0] ? counter2[15:0] : counterRegs2_0; // @[SourceDestination.scala 68:{23,23} 18:31]
  wire [15:0] _GEN_460 = 3'h1 == k[2:0] ? counter2[15:0] : counterRegs2_1; // @[SourceDestination.scala 68:{23,23} 18:31]
  wire [15:0] _GEN_461 = 3'h2 == k[2:0] ? counter2[15:0] : counterRegs2_2; // @[SourceDestination.scala 68:{23,23} 18:31]
  wire [15:0] _GEN_462 = 3'h3 == k[2:0] ? counter2[15:0] : counterRegs2_3; // @[SourceDestination.scala 68:{23,23} 18:31]
  wire [15:0] _GEN_463 = 3'h4 == k[2:0] ? counter2[15:0] : counterRegs2_4; // @[SourceDestination.scala 68:{23,23} 18:31]
  wire [15:0] _GEN_464 = 3'h5 == k[2:0] ? counter2[15:0] : counterRegs2_5; // @[SourceDestination.scala 68:{23,23} 18:31]
  wire [15:0] _GEN_465 = 3'h6 == k[2:0] ? counter2[15:0] : counterRegs2_6; // @[SourceDestination.scala 68:{23,23} 18:31]
  wire [15:0] _GEN_466 = 3'h7 == k[2:0] ? counter2[15:0] : counterRegs2_7; // @[SourceDestination.scala 68:{23,23} 18:31]
  wire [31:0] _counter2_T_1 = counter2 + 32'h1; // @[SourceDestination.scala 69:28]
  wire [15:0] _GEN_467 = _GEN_458 != 16'h0 ? _GEN_459 : counterRegs2_0; // @[SourceDestination.scala 18:31 67:43]
  wire [15:0] _GEN_468 = _GEN_458 != 16'h0 ? _GEN_460 : counterRegs2_1; // @[SourceDestination.scala 18:31 67:43]
  wire [15:0] _GEN_469 = _GEN_458 != 16'h0 ? _GEN_461 : counterRegs2_2; // @[SourceDestination.scala 18:31 67:43]
  wire [15:0] _GEN_470 = _GEN_458 != 16'h0 ? _GEN_462 : counterRegs2_3; // @[SourceDestination.scala 18:31 67:43]
  wire [15:0] _GEN_471 = _GEN_458 != 16'h0 ? _GEN_463 : counterRegs2_4; // @[SourceDestination.scala 18:31 67:43]
  wire [15:0] _GEN_472 = _GEN_458 != 16'h0 ? _GEN_464 : counterRegs2_5; // @[SourceDestination.scala 18:31 67:43]
  wire [15:0] _GEN_473 = _GEN_458 != 16'h0 ? _GEN_465 : counterRegs2_6; // @[SourceDestination.scala 18:31 67:43]
  wire [15:0] _GEN_474 = _GEN_458 != 16'h0 ? _GEN_466 : counterRegs2_7; // @[SourceDestination.scala 18:31 67:43]
  wire [31:0] _GEN_475 = _GEN_458 != 16'h0 ? _counter2_T_1 : counter2; // @[SourceDestination.scala 67:43 69:16 29:27]
  wire [31:0] _k_T_1 = k + 32'h1; // @[SourceDestination.scala 77:16]
  wire [31:0] _GEN_477 = k == 32'h7 ? k : _k_T_1; // @[SourceDestination.scala 73:37 74:9]
  wire [31:0] _GEN_478 = k == 32'h7 ? counter2 : _GEN_475; // @[SourceDestination.scala 73:37 75:16]
  wire [31:0] _j_T_1 = j + 32'h1; // @[SourceDestination.scala 81:16]
  wire [31:0] _i_T_1 = i + 32'h1; // @[SourceDestination.scala 87:18]
  wire [31:0] _GEN_479 = i < 32'h7 ? _i_T_1 : i; // @[SourceDestination.scala 86:42 87:13 20:20]
  wire [31:0] _GEN_481 = _reg_i_T_2 ? j : 32'h0; // @[SourceDestination.scala 21:20 82:83 85:11]
  wire [31:0] _GEN_482 = _reg_i_T_2 ? i : _GEN_479; // @[SourceDestination.scala 20:20 82:83]
  wire  _GEN_484 = j < 32'h7 ? 1'h0 : _reg_i_T_2; // @[SourceDestination.scala 49:12 80:40]
  wire  _GEN_564 = ~jValid & _GEN_484; // @[SourceDestination.scala 49:12 79:26]
  wire [31:0] _GEN_724 = io_start ? {{16'd0}, counterRegs1_0_0} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_725 = io_start ? {{16'd0}, counterRegs1_0_1} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_726 = io_start ? {{16'd0}, counterRegs1_0_2} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_727 = io_start ? {{16'd0}, counterRegs1_0_3} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_728 = io_start ? {{16'd0}, counterRegs1_0_4} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_729 = io_start ? {{16'd0}, counterRegs1_0_5} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_730 = io_start ? {{16'd0}, counterRegs1_0_6} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_731 = io_start ? {{16'd0}, counterRegs1_0_7} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_732 = io_start ? {{16'd0}, counterRegs1_1_0} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_733 = io_start ? {{16'd0}, counterRegs1_1_1} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_734 = io_start ? {{16'd0}, counterRegs1_1_2} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_735 = io_start ? {{16'd0}, counterRegs1_1_3} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_736 = io_start ? {{16'd0}, counterRegs1_1_4} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_737 = io_start ? {{16'd0}, counterRegs1_1_5} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_738 = io_start ? {{16'd0}, counterRegs1_1_6} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_739 = io_start ? {{16'd0}, counterRegs1_1_7} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_740 = io_start ? {{16'd0}, counterRegs1_2_0} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_741 = io_start ? {{16'd0}, counterRegs1_2_1} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_742 = io_start ? {{16'd0}, counterRegs1_2_2} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_743 = io_start ? {{16'd0}, counterRegs1_2_3} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_744 = io_start ? {{16'd0}, counterRegs1_2_4} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_745 = io_start ? {{16'd0}, counterRegs1_2_5} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_746 = io_start ? {{16'd0}, counterRegs1_2_6} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_747 = io_start ? {{16'd0}, counterRegs1_2_7} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_748 = io_start ? {{16'd0}, counterRegs1_3_0} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_749 = io_start ? {{16'd0}, counterRegs1_3_1} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_750 = io_start ? {{16'd0}, counterRegs1_3_2} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_751 = io_start ? {{16'd0}, counterRegs1_3_3} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_752 = io_start ? {{16'd0}, counterRegs1_3_4} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_753 = io_start ? {{16'd0}, counterRegs1_3_5} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_754 = io_start ? {{16'd0}, counterRegs1_3_6} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_755 = io_start ? {{16'd0}, counterRegs1_3_7} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_756 = io_start ? {{16'd0}, counterRegs1_4_0} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_757 = io_start ? {{16'd0}, counterRegs1_4_1} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_758 = io_start ? {{16'd0}, counterRegs1_4_2} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_759 = io_start ? {{16'd0}, counterRegs1_4_3} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_760 = io_start ? {{16'd0}, counterRegs1_4_4} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_761 = io_start ? {{16'd0}, counterRegs1_4_5} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_762 = io_start ? {{16'd0}, counterRegs1_4_6} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_763 = io_start ? {{16'd0}, counterRegs1_4_7} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_764 = io_start ? {{16'd0}, counterRegs1_5_0} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_765 = io_start ? {{16'd0}, counterRegs1_5_1} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_766 = io_start ? {{16'd0}, counterRegs1_5_2} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_767 = io_start ? {{16'd0}, counterRegs1_5_3} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_768 = io_start ? {{16'd0}, counterRegs1_5_4} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_769 = io_start ? {{16'd0}, counterRegs1_5_5} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_770 = io_start ? {{16'd0}, counterRegs1_5_6} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_771 = io_start ? {{16'd0}, counterRegs1_5_7} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_772 = io_start ? {{16'd0}, counterRegs1_6_0} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_773 = io_start ? {{16'd0}, counterRegs1_6_1} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_774 = io_start ? {{16'd0}, counterRegs1_6_2} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_775 = io_start ? {{16'd0}, counterRegs1_6_3} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_776 = io_start ? {{16'd0}, counterRegs1_6_4} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_777 = io_start ? {{16'd0}, counterRegs1_6_5} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_778 = io_start ? {{16'd0}, counterRegs1_6_6} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_779 = io_start ? {{16'd0}, counterRegs1_6_7} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_780 = io_start ? {{16'd0}, counterRegs1_7_0} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_781 = io_start ? {{16'd0}, counterRegs1_7_1} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_782 = io_start ? {{16'd0}, counterRegs1_7_2} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_783 = io_start ? {{16'd0}, counterRegs1_7_3} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_784 = io_start ? {{16'd0}, counterRegs1_7_4} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_785 = io_start ? {{16'd0}, counterRegs1_7_5} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_786 = io_start ? {{16'd0}, counterRegs1_7_6} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_787 = io_start ? {{16'd0}, counterRegs1_7_7} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_788 = io_start ? {{16'd0}, counterRegs2_0} : 32'h0; // @[SourceDestination.scala 34:17 115:28 119:26]
  wire [31:0] _GEN_789 = io_start ? {{16'd0}, counterRegs2_1} : 32'h0; // @[SourceDestination.scala 34:17 115:28 119:26]
  wire [31:0] _GEN_790 = io_start ? {{16'd0}, counterRegs2_2} : 32'h0; // @[SourceDestination.scala 34:17 115:28 119:26]
  wire [31:0] _GEN_791 = io_start ? {{16'd0}, counterRegs2_3} : 32'h0; // @[SourceDestination.scala 34:17 115:28 119:26]
  wire [31:0] _GEN_792 = io_start ? {{16'd0}, counterRegs2_4} : 32'h0; // @[SourceDestination.scala 34:17 115:28 119:26]
  wire [31:0] _GEN_793 = io_start ? {{16'd0}, counterRegs2_5} : 32'h0; // @[SourceDestination.scala 34:17 115:28 119:26]
  wire [31:0] _GEN_794 = io_start ? {{16'd0}, counterRegs2_6} : 32'h0; // @[SourceDestination.scala 34:17 115:28 119:26]
  wire [31:0] _GEN_795 = io_start ? {{16'd0}, counterRegs2_7} : 32'h0; // @[SourceDestination.scala 34:17 115:28 119:26]
  assign io_counterMatrix1_bits_0_0 = _GEN_724[15:0];
  assign io_counterMatrix1_bits_0_1 = _GEN_725[15:0];
  assign io_counterMatrix1_bits_0_2 = _GEN_726[15:0];
  assign io_counterMatrix1_bits_0_3 = _GEN_727[15:0];
  assign io_counterMatrix1_bits_0_4 = _GEN_728[15:0];
  assign io_counterMatrix1_bits_0_5 = _GEN_729[15:0];
  assign io_counterMatrix1_bits_0_6 = _GEN_730[15:0];
  assign io_counterMatrix1_bits_0_7 = _GEN_731[15:0];
  assign io_counterMatrix1_bits_1_0 = _GEN_732[15:0];
  assign io_counterMatrix1_bits_1_1 = _GEN_733[15:0];
  assign io_counterMatrix1_bits_1_2 = _GEN_734[15:0];
  assign io_counterMatrix1_bits_1_3 = _GEN_735[15:0];
  assign io_counterMatrix1_bits_1_4 = _GEN_736[15:0];
  assign io_counterMatrix1_bits_1_5 = _GEN_737[15:0];
  assign io_counterMatrix1_bits_1_6 = _GEN_738[15:0];
  assign io_counterMatrix1_bits_1_7 = _GEN_739[15:0];
  assign io_counterMatrix1_bits_2_0 = _GEN_740[15:0];
  assign io_counterMatrix1_bits_2_1 = _GEN_741[15:0];
  assign io_counterMatrix1_bits_2_2 = _GEN_742[15:0];
  assign io_counterMatrix1_bits_2_3 = _GEN_743[15:0];
  assign io_counterMatrix1_bits_2_4 = _GEN_744[15:0];
  assign io_counterMatrix1_bits_2_5 = _GEN_745[15:0];
  assign io_counterMatrix1_bits_2_6 = _GEN_746[15:0];
  assign io_counterMatrix1_bits_2_7 = _GEN_747[15:0];
  assign io_counterMatrix1_bits_3_0 = _GEN_748[15:0];
  assign io_counterMatrix1_bits_3_1 = _GEN_749[15:0];
  assign io_counterMatrix1_bits_3_2 = _GEN_750[15:0];
  assign io_counterMatrix1_bits_3_3 = _GEN_751[15:0];
  assign io_counterMatrix1_bits_3_4 = _GEN_752[15:0];
  assign io_counterMatrix1_bits_3_5 = _GEN_753[15:0];
  assign io_counterMatrix1_bits_3_6 = _GEN_754[15:0];
  assign io_counterMatrix1_bits_3_7 = _GEN_755[15:0];
  assign io_counterMatrix1_bits_4_0 = _GEN_756[15:0];
  assign io_counterMatrix1_bits_4_1 = _GEN_757[15:0];
  assign io_counterMatrix1_bits_4_2 = _GEN_758[15:0];
  assign io_counterMatrix1_bits_4_3 = _GEN_759[15:0];
  assign io_counterMatrix1_bits_4_4 = _GEN_760[15:0];
  assign io_counterMatrix1_bits_4_5 = _GEN_761[15:0];
  assign io_counterMatrix1_bits_4_6 = _GEN_762[15:0];
  assign io_counterMatrix1_bits_4_7 = _GEN_763[15:0];
  assign io_counterMatrix1_bits_5_0 = _GEN_764[15:0];
  assign io_counterMatrix1_bits_5_1 = _GEN_765[15:0];
  assign io_counterMatrix1_bits_5_2 = _GEN_766[15:0];
  assign io_counterMatrix1_bits_5_3 = _GEN_767[15:0];
  assign io_counterMatrix1_bits_5_4 = _GEN_768[15:0];
  assign io_counterMatrix1_bits_5_5 = _GEN_769[15:0];
  assign io_counterMatrix1_bits_5_6 = _GEN_770[15:0];
  assign io_counterMatrix1_bits_5_7 = _GEN_771[15:0];
  assign io_counterMatrix1_bits_6_0 = _GEN_772[15:0];
  assign io_counterMatrix1_bits_6_1 = _GEN_773[15:0];
  assign io_counterMatrix1_bits_6_2 = _GEN_774[15:0];
  assign io_counterMatrix1_bits_6_3 = _GEN_775[15:0];
  assign io_counterMatrix1_bits_6_4 = _GEN_776[15:0];
  assign io_counterMatrix1_bits_6_5 = _GEN_777[15:0];
  assign io_counterMatrix1_bits_6_6 = _GEN_778[15:0];
  assign io_counterMatrix1_bits_6_7 = _GEN_779[15:0];
  assign io_counterMatrix1_bits_7_0 = _GEN_780[15:0];
  assign io_counterMatrix1_bits_7_1 = _GEN_781[15:0];
  assign io_counterMatrix1_bits_7_2 = _GEN_782[15:0];
  assign io_counterMatrix1_bits_7_3 = _GEN_783[15:0];
  assign io_counterMatrix1_bits_7_4 = _GEN_784[15:0];
  assign io_counterMatrix1_bits_7_5 = _GEN_785[15:0];
  assign io_counterMatrix1_bits_7_6 = _GEN_786[15:0];
  assign io_counterMatrix1_bits_7_7 = _GEN_787[15:0];
  assign io_counterMatrix2_bits_0 = _GEN_788[15:0];
  assign io_counterMatrix2_bits_1 = _GEN_789[15:0];
  assign io_counterMatrix2_bits_2 = _GEN_790[15:0];
  assign io_counterMatrix2_bits_3 = _GEN_791[15:0];
  assign io_counterMatrix2_bits_4 = _GEN_792[15:0];
  assign io_counterMatrix2_bits_5 = _GEN_793[15:0];
  assign io_counterMatrix2_bits_6 = _GEN_794[15:0];
  assign io_counterMatrix2_bits_7 = _GEN_795[15:0];
  assign io_valid = io_start & (i == 32'h3 & j == 32'h3); // @[SourceDestination.scala 104:14 122:12 34:17]
  always @(posedge clock) begin
    prevStationary_matrix_0_0 <= io_Stationary_matrix_0_0; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_0_1 <= io_Stationary_matrix_0_1; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_0_2 <= io_Stationary_matrix_0_2; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_0_3 <= io_Stationary_matrix_0_3; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_0_4 <= io_Stationary_matrix_0_4; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_0_5 <= io_Stationary_matrix_0_5; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_0_6 <= io_Stationary_matrix_0_6; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_0_7 <= io_Stationary_matrix_0_7; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_1_0 <= io_Stationary_matrix_1_0; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_1_1 <= io_Stationary_matrix_1_1; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_1_2 <= io_Stationary_matrix_1_2; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_1_3 <= io_Stationary_matrix_1_3; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_1_4 <= io_Stationary_matrix_1_4; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_1_5 <= io_Stationary_matrix_1_5; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_1_6 <= io_Stationary_matrix_1_6; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_1_7 <= io_Stationary_matrix_1_7; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_2_0 <= io_Stationary_matrix_2_0; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_2_1 <= io_Stationary_matrix_2_1; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_2_2 <= io_Stationary_matrix_2_2; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_2_3 <= io_Stationary_matrix_2_3; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_2_4 <= io_Stationary_matrix_2_4; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_2_5 <= io_Stationary_matrix_2_5; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_2_6 <= io_Stationary_matrix_2_6; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_2_7 <= io_Stationary_matrix_2_7; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_3_0 <= io_Stationary_matrix_3_0; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_3_1 <= io_Stationary_matrix_3_1; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_3_2 <= io_Stationary_matrix_3_2; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_3_3 <= io_Stationary_matrix_3_3; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_3_4 <= io_Stationary_matrix_3_4; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_3_5 <= io_Stationary_matrix_3_5; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_3_6 <= io_Stationary_matrix_3_6; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_3_7 <= io_Stationary_matrix_3_7; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_4_0 <= io_Stationary_matrix_4_0; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_4_1 <= io_Stationary_matrix_4_1; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_4_2 <= io_Stationary_matrix_4_2; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_4_3 <= io_Stationary_matrix_4_3; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_4_4 <= io_Stationary_matrix_4_4; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_4_5 <= io_Stationary_matrix_4_5; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_4_6 <= io_Stationary_matrix_4_6; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_4_7 <= io_Stationary_matrix_4_7; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_5_0 <= io_Stationary_matrix_5_0; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_5_1 <= io_Stationary_matrix_5_1; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_5_2 <= io_Stationary_matrix_5_2; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_5_3 <= io_Stationary_matrix_5_3; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_5_4 <= io_Stationary_matrix_5_4; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_5_5 <= io_Stationary_matrix_5_5; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_5_6 <= io_Stationary_matrix_5_6; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_5_7 <= io_Stationary_matrix_5_7; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_6_0 <= io_Stationary_matrix_6_0; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_6_1 <= io_Stationary_matrix_6_1; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_6_2 <= io_Stationary_matrix_6_2; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_6_3 <= io_Stationary_matrix_6_3; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_6_4 <= io_Stationary_matrix_6_4; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_6_5 <= io_Stationary_matrix_6_5; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_6_6 <= io_Stationary_matrix_6_6; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_6_7 <= io_Stationary_matrix_6_7; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_7_0 <= io_Stationary_matrix_7_0; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_7_1 <= io_Stationary_matrix_7_1; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_7_2 <= io_Stationary_matrix_7_2; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_7_3 <= io_Stationary_matrix_7_3; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_7_4 <= io_Stationary_matrix_7_4; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_7_5 <= io_Stationary_matrix_7_5; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_7_6 <= io_Stationary_matrix_7_6; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_7_7 <= io_Stationary_matrix_7_7; // @[SourceDestination.scala 15:40]
    if (io_start) begin // @[SourceDestination.scala 34:17]
      if (io_Stationary_matrix_7_7 != prevStationary_matrix_7_7) begin // @[SourceDestination.scala 40:74]
        matricesAreEqual <= 1'h0; // @[SourceDestination.scala 41:28]
      end else if (io_Stationary_matrix_7_6 != prevStationary_matrix_7_6) begin // @[SourceDestination.scala 40:74]
        matricesAreEqual <= 1'h0; // @[SourceDestination.scala 41:28]
      end else if (io_Stationary_matrix_7_5 != prevStationary_matrix_7_5) begin // @[SourceDestination.scala 40:74]
        matricesAreEqual <= 1'h0; // @[SourceDestination.scala 41:28]
      end else begin
        matricesAreEqual <= _GEN_60;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_0_0 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_0_0 <= _GEN_386;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_0_0 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_0_0 <= _GEN_386;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_0_1 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_0_1 <= _GEN_387;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_0_1 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_0_1 <= _GEN_387;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_0_2 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_0_2 <= _GEN_388;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_0_2 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_0_2 <= _GEN_388;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_0_3 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_0_3 <= _GEN_389;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_0_3 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_0_3 <= _GEN_389;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_0_4 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_0_4 <= _GEN_390;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_0_4 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_0_4 <= _GEN_390;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_0_5 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_0_5 <= _GEN_391;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_0_5 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_0_5 <= _GEN_391;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_0_6 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_0_6 <= _GEN_392;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_0_6 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_0_6 <= _GEN_392;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_0_7 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_0_7 <= _GEN_393;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_0_7 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_0_7 <= _GEN_393;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_1_0 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_1_0 <= _GEN_394;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_1_0 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_1_0 <= _GEN_394;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_1_1 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_1_1 <= _GEN_395;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_1_1 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_1_1 <= _GEN_395;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_1_2 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_1_2 <= _GEN_396;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_1_2 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_1_2 <= _GEN_396;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_1_3 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_1_3 <= _GEN_397;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_1_3 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_1_3 <= _GEN_397;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_1_4 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_1_4 <= _GEN_398;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_1_4 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_1_4 <= _GEN_398;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_1_5 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_1_5 <= _GEN_399;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_1_5 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_1_5 <= _GEN_399;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_1_6 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_1_6 <= _GEN_400;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_1_6 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_1_6 <= _GEN_400;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_1_7 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_1_7 <= _GEN_401;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_1_7 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_1_7 <= _GEN_401;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_2_0 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_2_0 <= _GEN_402;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_2_0 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_2_0 <= _GEN_402;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_2_1 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_2_1 <= _GEN_403;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_2_1 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_2_1 <= _GEN_403;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_2_2 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_2_2 <= _GEN_404;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_2_2 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_2_2 <= _GEN_404;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_2_3 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_2_3 <= _GEN_405;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_2_3 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_2_3 <= _GEN_405;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_2_4 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_2_4 <= _GEN_406;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_2_4 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_2_4 <= _GEN_406;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_2_5 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_2_5 <= _GEN_407;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_2_5 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_2_5 <= _GEN_407;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_2_6 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_2_6 <= _GEN_408;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_2_6 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_2_6 <= _GEN_408;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_2_7 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_2_7 <= _GEN_409;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_2_7 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_2_7 <= _GEN_409;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_3_0 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_3_0 <= _GEN_410;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_3_0 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_3_0 <= _GEN_410;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_3_1 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_3_1 <= _GEN_411;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_3_1 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_3_1 <= _GEN_411;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_3_2 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_3_2 <= _GEN_412;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_3_2 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_3_2 <= _GEN_412;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_3_3 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_3_3 <= _GEN_413;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_3_3 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_3_3 <= _GEN_413;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_3_4 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_3_4 <= _GEN_414;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_3_4 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_3_4 <= _GEN_414;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_3_5 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_3_5 <= _GEN_415;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_3_5 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_3_5 <= _GEN_415;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_3_6 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_3_6 <= _GEN_416;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_3_6 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_3_6 <= _GEN_416;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_3_7 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_3_7 <= _GEN_417;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_3_7 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_3_7 <= _GEN_417;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_4_0 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_4_0 <= _GEN_418;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_4_0 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_4_0 <= _GEN_418;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_4_1 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_4_1 <= _GEN_419;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_4_1 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_4_1 <= _GEN_419;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_4_2 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_4_2 <= _GEN_420;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_4_2 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_4_2 <= _GEN_420;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_4_3 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_4_3 <= _GEN_421;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_4_3 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_4_3 <= _GEN_421;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_4_4 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_4_4 <= _GEN_422;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_4_4 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_4_4 <= _GEN_422;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_4_5 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_4_5 <= _GEN_423;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_4_5 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_4_5 <= _GEN_423;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_4_6 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_4_6 <= _GEN_424;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_4_6 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_4_6 <= _GEN_424;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_4_7 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_4_7 <= _GEN_425;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_4_7 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_4_7 <= _GEN_425;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_5_0 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_5_0 <= _GEN_426;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_5_0 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_5_0 <= _GEN_426;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_5_1 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_5_1 <= _GEN_427;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_5_1 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_5_1 <= _GEN_427;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_5_2 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_5_2 <= _GEN_428;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_5_2 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_5_2 <= _GEN_428;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_5_3 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_5_3 <= _GEN_429;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_5_3 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_5_3 <= _GEN_429;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_5_4 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_5_4 <= _GEN_430;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_5_4 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_5_4 <= _GEN_430;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_5_5 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_5_5 <= _GEN_431;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_5_5 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_5_5 <= _GEN_431;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_5_6 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_5_6 <= _GEN_432;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_5_6 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_5_6 <= _GEN_432;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_5_7 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_5_7 <= _GEN_433;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_5_7 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_5_7 <= _GEN_433;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_6_0 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_6_0 <= _GEN_434;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_6_0 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_6_0 <= _GEN_434;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_6_1 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_6_1 <= _GEN_435;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_6_1 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_6_1 <= _GEN_435;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_6_2 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_6_2 <= _GEN_436;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_6_2 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_6_2 <= _GEN_436;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_6_3 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_6_3 <= _GEN_437;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_6_3 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_6_3 <= _GEN_437;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_6_4 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_6_4 <= _GEN_438;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_6_4 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_6_4 <= _GEN_438;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_6_5 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_6_5 <= _GEN_439;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_6_5 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_6_5 <= _GEN_439;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_6_6 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_6_6 <= _GEN_440;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_6_6 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_6_6 <= _GEN_440;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_6_7 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_6_7 <= _GEN_441;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_6_7 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_6_7 <= _GEN_441;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_7_0 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_7_0 <= _GEN_442;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_7_0 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_7_0 <= _GEN_442;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_7_1 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_7_1 <= _GEN_443;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_7_1 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_7_1 <= _GEN_443;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_7_2 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_7_2 <= _GEN_444;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_7_2 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_7_2 <= _GEN_444;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_7_3 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_7_3 <= _GEN_445;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_7_3 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_7_3 <= _GEN_445;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_7_4 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_7_4 <= _GEN_446;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_7_4 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_7_4 <= _GEN_446;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_7_5 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_7_5 <= _GEN_447;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_7_5 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_7_5 <= _GEN_447;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_7_6 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_7_6 <= _GEN_448;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_7_6 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_7_6 <= _GEN_448;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_7_7 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_7_7 <= _GEN_449;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_7_7 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_7_7 <= _GEN_449;
      end
    end
    if (reset) begin // @[SourceDestination.scala 18:31]
      counterRegs2_0 <= 16'h0; // @[SourceDestination.scala 18:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs2_0 <= _GEN_467;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs2_0 <= 16'h0; // @[SourceDestination.scala 100:25]
      end else begin
        counterRegs2_0 <= _GEN_467;
      end
    end
    if (reset) begin // @[SourceDestination.scala 18:31]
      counterRegs2_1 <= 16'h0; // @[SourceDestination.scala 18:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs2_1 <= _GEN_468;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs2_1 <= 16'h0; // @[SourceDestination.scala 100:25]
      end else begin
        counterRegs2_1 <= _GEN_468;
      end
    end
    if (reset) begin // @[SourceDestination.scala 18:31]
      counterRegs2_2 <= 16'h0; // @[SourceDestination.scala 18:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs2_2 <= _GEN_469;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs2_2 <= 16'h0; // @[SourceDestination.scala 100:25]
      end else begin
        counterRegs2_2 <= _GEN_469;
      end
    end
    if (reset) begin // @[SourceDestination.scala 18:31]
      counterRegs2_3 <= 16'h0; // @[SourceDestination.scala 18:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs2_3 <= _GEN_470;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs2_3 <= 16'h0; // @[SourceDestination.scala 100:25]
      end else begin
        counterRegs2_3 <= _GEN_470;
      end
    end
    if (reset) begin // @[SourceDestination.scala 18:31]
      counterRegs2_4 <= 16'h0; // @[SourceDestination.scala 18:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs2_4 <= _GEN_471;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs2_4 <= 16'h0; // @[SourceDestination.scala 100:25]
      end else begin
        counterRegs2_4 <= _GEN_471;
      end
    end
    if (reset) begin // @[SourceDestination.scala 18:31]
      counterRegs2_5 <= 16'h0; // @[SourceDestination.scala 18:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs2_5 <= _GEN_472;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs2_5 <= 16'h0; // @[SourceDestination.scala 100:25]
      end else begin
        counterRegs2_5 <= _GEN_472;
      end
    end
    if (reset) begin // @[SourceDestination.scala 18:31]
      counterRegs2_6 <= 16'h0; // @[SourceDestination.scala 18:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs2_6 <= _GEN_473;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs2_6 <= 16'h0; // @[SourceDestination.scala 100:25]
      end else begin
        counterRegs2_6 <= _GEN_473;
      end
    end
    if (reset) begin // @[SourceDestination.scala 18:31]
      counterRegs2_7 <= 16'h0; // @[SourceDestination.scala 18:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs2_7 <= _GEN_474;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs2_7 <= 16'h0; // @[SourceDestination.scala 100:25]
      end else begin
        counterRegs2_7 <= _GEN_474;
      end
    end
    if (reset) begin // @[SourceDestination.scala 20:20]
      i <= 32'h0; // @[SourceDestination.scala 20:20]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        if (!(j < 32'h7)) begin // @[SourceDestination.scala 80:40]
          i <= _GEN_482;
        end
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        i <= 32'h0; // @[SourceDestination.scala 91:9]
      end
    end
    if (reset) begin // @[SourceDestination.scala 21:20]
      j <= 32'h0; // @[SourceDestination.scala 21:20]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        if (j < 32'h7) begin // @[SourceDestination.scala 80:40]
          j <= _j_T_1; // @[SourceDestination.scala 81:11]
        end else begin
          j <= _GEN_481;
        end
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        j <= 32'h0; // @[SourceDestination.scala 92:9]
      end
    end
    if (io_start) begin // @[SourceDestination.scala 34:17]
      jValid <= _GEN_564;
    end
    if (reset) begin // @[SourceDestination.scala 26:20]
      k <= 32'h0; // @[SourceDestination.scala 26:20]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        k <= _GEN_477;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        k <= 32'h0; // @[SourceDestination.scala 93:9]
      end else begin
        k <= _GEN_477;
      end
    end
    if (reset) begin // @[SourceDestination.scala 28:27]
      counter1 <= 32'h1; // @[SourceDestination.scala 28:27]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counter1 <= _GEN_450;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counter1 <= 32'h1; // @[SourceDestination.scala 94:16]
      end else begin
        counter1 <= _GEN_450;
      end
    end
    if (reset) begin // @[SourceDestination.scala 29:27]
      counter2 <= 32'h1; // @[SourceDestination.scala 29:27]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counter2 <= _GEN_478;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counter2 <= 32'h1; // @[SourceDestination.scala 95:16]
      end else begin
        counter2 <= _GEN_478;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  prevStationary_matrix_0_0 = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  prevStationary_matrix_0_1 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  prevStationary_matrix_0_2 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  prevStationary_matrix_0_3 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  prevStationary_matrix_0_4 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  prevStationary_matrix_0_5 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  prevStationary_matrix_0_6 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  prevStationary_matrix_0_7 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  prevStationary_matrix_1_0 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  prevStationary_matrix_1_1 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  prevStationary_matrix_1_2 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  prevStationary_matrix_1_3 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  prevStationary_matrix_1_4 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  prevStationary_matrix_1_5 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  prevStationary_matrix_1_6 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  prevStationary_matrix_1_7 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  prevStationary_matrix_2_0 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  prevStationary_matrix_2_1 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  prevStationary_matrix_2_2 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  prevStationary_matrix_2_3 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  prevStationary_matrix_2_4 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  prevStationary_matrix_2_5 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  prevStationary_matrix_2_6 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  prevStationary_matrix_2_7 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  prevStationary_matrix_3_0 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  prevStationary_matrix_3_1 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  prevStationary_matrix_3_2 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  prevStationary_matrix_3_3 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  prevStationary_matrix_3_4 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  prevStationary_matrix_3_5 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  prevStationary_matrix_3_6 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  prevStationary_matrix_3_7 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  prevStationary_matrix_4_0 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  prevStationary_matrix_4_1 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  prevStationary_matrix_4_2 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  prevStationary_matrix_4_3 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  prevStationary_matrix_4_4 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  prevStationary_matrix_4_5 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  prevStationary_matrix_4_6 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  prevStationary_matrix_4_7 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  prevStationary_matrix_5_0 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  prevStationary_matrix_5_1 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  prevStationary_matrix_5_2 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  prevStationary_matrix_5_3 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  prevStationary_matrix_5_4 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  prevStationary_matrix_5_5 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  prevStationary_matrix_5_6 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  prevStationary_matrix_5_7 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  prevStationary_matrix_6_0 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  prevStationary_matrix_6_1 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  prevStationary_matrix_6_2 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  prevStationary_matrix_6_3 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  prevStationary_matrix_6_4 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  prevStationary_matrix_6_5 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  prevStationary_matrix_6_6 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  prevStationary_matrix_6_7 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  prevStationary_matrix_7_0 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  prevStationary_matrix_7_1 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  prevStationary_matrix_7_2 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  prevStationary_matrix_7_3 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  prevStationary_matrix_7_4 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  prevStationary_matrix_7_5 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  prevStationary_matrix_7_6 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  prevStationary_matrix_7_7 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  matricesAreEqual = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  counterRegs1_0_0 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  counterRegs1_0_1 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  counterRegs1_0_2 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  counterRegs1_0_3 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  counterRegs1_0_4 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  counterRegs1_0_5 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  counterRegs1_0_6 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  counterRegs1_0_7 = _RAND_72[15:0];
  _RAND_73 = {1{`RANDOM}};
  counterRegs1_1_0 = _RAND_73[15:0];
  _RAND_74 = {1{`RANDOM}};
  counterRegs1_1_1 = _RAND_74[15:0];
  _RAND_75 = {1{`RANDOM}};
  counterRegs1_1_2 = _RAND_75[15:0];
  _RAND_76 = {1{`RANDOM}};
  counterRegs1_1_3 = _RAND_76[15:0];
  _RAND_77 = {1{`RANDOM}};
  counterRegs1_1_4 = _RAND_77[15:0];
  _RAND_78 = {1{`RANDOM}};
  counterRegs1_1_5 = _RAND_78[15:0];
  _RAND_79 = {1{`RANDOM}};
  counterRegs1_1_6 = _RAND_79[15:0];
  _RAND_80 = {1{`RANDOM}};
  counterRegs1_1_7 = _RAND_80[15:0];
  _RAND_81 = {1{`RANDOM}};
  counterRegs1_2_0 = _RAND_81[15:0];
  _RAND_82 = {1{`RANDOM}};
  counterRegs1_2_1 = _RAND_82[15:0];
  _RAND_83 = {1{`RANDOM}};
  counterRegs1_2_2 = _RAND_83[15:0];
  _RAND_84 = {1{`RANDOM}};
  counterRegs1_2_3 = _RAND_84[15:0];
  _RAND_85 = {1{`RANDOM}};
  counterRegs1_2_4 = _RAND_85[15:0];
  _RAND_86 = {1{`RANDOM}};
  counterRegs1_2_5 = _RAND_86[15:0];
  _RAND_87 = {1{`RANDOM}};
  counterRegs1_2_6 = _RAND_87[15:0];
  _RAND_88 = {1{`RANDOM}};
  counterRegs1_2_7 = _RAND_88[15:0];
  _RAND_89 = {1{`RANDOM}};
  counterRegs1_3_0 = _RAND_89[15:0];
  _RAND_90 = {1{`RANDOM}};
  counterRegs1_3_1 = _RAND_90[15:0];
  _RAND_91 = {1{`RANDOM}};
  counterRegs1_3_2 = _RAND_91[15:0];
  _RAND_92 = {1{`RANDOM}};
  counterRegs1_3_3 = _RAND_92[15:0];
  _RAND_93 = {1{`RANDOM}};
  counterRegs1_3_4 = _RAND_93[15:0];
  _RAND_94 = {1{`RANDOM}};
  counterRegs1_3_5 = _RAND_94[15:0];
  _RAND_95 = {1{`RANDOM}};
  counterRegs1_3_6 = _RAND_95[15:0];
  _RAND_96 = {1{`RANDOM}};
  counterRegs1_3_7 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  counterRegs1_4_0 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  counterRegs1_4_1 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  counterRegs1_4_2 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  counterRegs1_4_3 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  counterRegs1_4_4 = _RAND_101[15:0];
  _RAND_102 = {1{`RANDOM}};
  counterRegs1_4_5 = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  counterRegs1_4_6 = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  counterRegs1_4_7 = _RAND_104[15:0];
  _RAND_105 = {1{`RANDOM}};
  counterRegs1_5_0 = _RAND_105[15:0];
  _RAND_106 = {1{`RANDOM}};
  counterRegs1_5_1 = _RAND_106[15:0];
  _RAND_107 = {1{`RANDOM}};
  counterRegs1_5_2 = _RAND_107[15:0];
  _RAND_108 = {1{`RANDOM}};
  counterRegs1_5_3 = _RAND_108[15:0];
  _RAND_109 = {1{`RANDOM}};
  counterRegs1_5_4 = _RAND_109[15:0];
  _RAND_110 = {1{`RANDOM}};
  counterRegs1_5_5 = _RAND_110[15:0];
  _RAND_111 = {1{`RANDOM}};
  counterRegs1_5_6 = _RAND_111[15:0];
  _RAND_112 = {1{`RANDOM}};
  counterRegs1_5_7 = _RAND_112[15:0];
  _RAND_113 = {1{`RANDOM}};
  counterRegs1_6_0 = _RAND_113[15:0];
  _RAND_114 = {1{`RANDOM}};
  counterRegs1_6_1 = _RAND_114[15:0];
  _RAND_115 = {1{`RANDOM}};
  counterRegs1_6_2 = _RAND_115[15:0];
  _RAND_116 = {1{`RANDOM}};
  counterRegs1_6_3 = _RAND_116[15:0];
  _RAND_117 = {1{`RANDOM}};
  counterRegs1_6_4 = _RAND_117[15:0];
  _RAND_118 = {1{`RANDOM}};
  counterRegs1_6_5 = _RAND_118[15:0];
  _RAND_119 = {1{`RANDOM}};
  counterRegs1_6_6 = _RAND_119[15:0];
  _RAND_120 = {1{`RANDOM}};
  counterRegs1_6_7 = _RAND_120[15:0];
  _RAND_121 = {1{`RANDOM}};
  counterRegs1_7_0 = _RAND_121[15:0];
  _RAND_122 = {1{`RANDOM}};
  counterRegs1_7_1 = _RAND_122[15:0];
  _RAND_123 = {1{`RANDOM}};
  counterRegs1_7_2 = _RAND_123[15:0];
  _RAND_124 = {1{`RANDOM}};
  counterRegs1_7_3 = _RAND_124[15:0];
  _RAND_125 = {1{`RANDOM}};
  counterRegs1_7_4 = _RAND_125[15:0];
  _RAND_126 = {1{`RANDOM}};
  counterRegs1_7_5 = _RAND_126[15:0];
  _RAND_127 = {1{`RANDOM}};
  counterRegs1_7_6 = _RAND_127[15:0];
  _RAND_128 = {1{`RANDOM}};
  counterRegs1_7_7 = _RAND_128[15:0];
  _RAND_129 = {1{`RANDOM}};
  counterRegs2_0 = _RAND_129[15:0];
  _RAND_130 = {1{`RANDOM}};
  counterRegs2_1 = _RAND_130[15:0];
  _RAND_131 = {1{`RANDOM}};
  counterRegs2_2 = _RAND_131[15:0];
  _RAND_132 = {1{`RANDOM}};
  counterRegs2_3 = _RAND_132[15:0];
  _RAND_133 = {1{`RANDOM}};
  counterRegs2_4 = _RAND_133[15:0];
  _RAND_134 = {1{`RANDOM}};
  counterRegs2_5 = _RAND_134[15:0];
  _RAND_135 = {1{`RANDOM}};
  counterRegs2_6 = _RAND_135[15:0];
  _RAND_136 = {1{`RANDOM}};
  counterRegs2_7 = _RAND_136[15:0];
  _RAND_137 = {1{`RANDOM}};
  i = _RAND_137[31:0];
  _RAND_138 = {1{`RANDOM}};
  j = _RAND_138[31:0];
  _RAND_139 = {1{`RANDOM}};
  jValid = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  k = _RAND_140[31:0];
  _RAND_141 = {1{`RANDOM}};
  counter1 = _RAND_141[31:0];
  _RAND_142 = {1{`RANDOM}};
  counter2 = _RAND_142[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module abc2(
  input         clock,
  input         reset,
  input  [31:0] io_IDex,
  input  [31:0] io_JDex,
  input         io_valid,
  input  [31:0] io_mat_0_0,
  input  [31:0] io_mat_0_1,
  input  [31:0] io_mat_0_2,
  input  [31:0] io_mat_0_3,
  input  [31:0] io_mat_0_4,
  input  [31:0] io_mat_0_5,
  input  [31:0] io_mat_0_6,
  input  [31:0] io_mat_0_7,
  input  [31:0] io_mat_1_0,
  input  [31:0] io_mat_1_1,
  input  [31:0] io_mat_1_2,
  input  [31:0] io_mat_1_3,
  input  [31:0] io_mat_1_4,
  input  [31:0] io_mat_1_5,
  input  [31:0] io_mat_1_6,
  input  [31:0] io_mat_1_7,
  input  [31:0] io_mat_2_0,
  input  [31:0] io_mat_2_1,
  input  [31:0] io_mat_2_2,
  input  [31:0] io_mat_2_3,
  input  [31:0] io_mat_2_4,
  input  [31:0] io_mat_2_5,
  input  [31:0] io_mat_2_6,
  input  [31:0] io_mat_2_7,
  input  [31:0] io_mat_3_0,
  input  [31:0] io_mat_3_1,
  input  [31:0] io_mat_3_2,
  input  [31:0] io_mat_3_3,
  input  [31:0] io_mat_3_4,
  input  [31:0] io_mat_3_5,
  input  [31:0] io_mat_3_6,
  input  [31:0] io_mat_3_7,
  input  [31:0] io_mat_4_0,
  input  [31:0] io_mat_4_1,
  input  [31:0] io_mat_4_2,
  input  [31:0] io_mat_4_3,
  input  [31:0] io_mat_4_4,
  input  [31:0] io_mat_4_5,
  input  [31:0] io_mat_4_6,
  input  [31:0] io_mat_4_7,
  input  [31:0] io_mat_5_0,
  input  [31:0] io_mat_5_1,
  input  [31:0] io_mat_5_2,
  input  [31:0] io_mat_5_3,
  input  [31:0] io_mat_5_4,
  input  [31:0] io_mat_5_5,
  input  [31:0] io_mat_5_6,
  input  [31:0] io_mat_5_7,
  input  [31:0] io_mat_6_0,
  input  [31:0] io_mat_6_1,
  input  [31:0] io_mat_6_2,
  input  [31:0] io_mat_6_3,
  input  [31:0] io_mat_6_4,
  input  [31:0] io_mat_6_5,
  input  [31:0] io_mat_6_6,
  input  [31:0] io_mat_6_7,
  input  [31:0] io_mat_7_0,
  input  [31:0] io_mat_7_1,
  input  [31:0] io_mat_7_2,
  input  [31:0] io_mat_7_3,
  input  [31:0] io_mat_7_4,
  input  [31:0] io_mat_7_5,
  input  [31:0] io_mat_7_6,
  input  [31:0] io_mat_7_7,
  output [31:0] io_OutMat_0_0,
  output [31:0] io_OutMat_0_1,
  output [31:0] io_OutMat_0_2,
  output [31:0] io_OutMat_0_3,
  output [31:0] io_OutMat_0_4,
  output [31:0] io_OutMat_0_5,
  output [31:0] io_OutMat_0_6,
  output [31:0] io_OutMat_0_7,
  output [31:0] io_OutMat_1_0,
  output [31:0] io_OutMat_1_1,
  output [31:0] io_OutMat_1_2,
  output [31:0] io_OutMat_1_3,
  output [31:0] io_OutMat_1_4,
  output [31:0] io_OutMat_1_5,
  output [31:0] io_OutMat_1_6,
  output [31:0] io_OutMat_1_7,
  output [31:0] io_OutMat_2_0,
  output [31:0] io_OutMat_2_1,
  output [31:0] io_OutMat_2_2,
  output [31:0] io_OutMat_2_3,
  output [31:0] io_OutMat_2_4,
  output [31:0] io_OutMat_2_5,
  output [31:0] io_OutMat_2_6,
  output [31:0] io_OutMat_2_7,
  output [31:0] io_OutMat_3_0,
  output [31:0] io_OutMat_3_1,
  output [31:0] io_OutMat_3_2,
  output [31:0] io_OutMat_3_3,
  output [31:0] io_OutMat_3_4,
  output [31:0] io_OutMat_3_5,
  output [31:0] io_OutMat_3_6,
  output [31:0] io_OutMat_3_7,
  output [31:0] io_OutMat_4_0,
  output [31:0] io_OutMat_4_1,
  output [31:0] io_OutMat_4_2,
  output [31:0] io_OutMat_4_3,
  output [31:0] io_OutMat_4_4,
  output [31:0] io_OutMat_4_5,
  output [31:0] io_OutMat_4_6,
  output [31:0] io_OutMat_4_7,
  output [31:0] io_OutMat_5_0,
  output [31:0] io_OutMat_5_1,
  output [31:0] io_OutMat_5_2,
  output [31:0] io_OutMat_5_3,
  output [31:0] io_OutMat_5_4,
  output [31:0] io_OutMat_5_5,
  output [31:0] io_OutMat_5_6,
  output [31:0] io_OutMat_5_7,
  output [31:0] io_OutMat_6_0,
  output [31:0] io_OutMat_6_1,
  output [31:0] io_OutMat_6_2,
  output [31:0] io_OutMat_6_3,
  output [31:0] io_OutMat_6_4,
  output [31:0] io_OutMat_6_5,
  output [31:0] io_OutMat_6_6,
  output [31:0] io_OutMat_6_7,
  output [31:0] io_OutMat_7_0,
  output [31:0] io_OutMat_7_1,
  output [31:0] io_OutMat_7_2,
  output [31:0] io_OutMat_7_3,
  output [31:0] io_OutMat_7_4,
  output [31:0] io_OutMat_7_5,
  output [31:0] io_OutMat_7_6,
  output [31:0] io_OutMat_7_7,
  output        io_Ovalid,
  output        io_ProcessValid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] b_0_0; // @[singleLoop.scala 19:20]
  reg [31:0] b_0_1; // @[singleLoop.scala 19:20]
  reg [31:0] b_0_2; // @[singleLoop.scala 19:20]
  reg [31:0] b_0_3; // @[singleLoop.scala 19:20]
  reg [31:0] b_0_4; // @[singleLoop.scala 19:20]
  reg [31:0] b_0_5; // @[singleLoop.scala 19:20]
  reg [31:0] b_0_6; // @[singleLoop.scala 19:20]
  reg [31:0] b_0_7; // @[singleLoop.scala 19:20]
  reg [31:0] b_1_0; // @[singleLoop.scala 19:20]
  reg [31:0] b_1_1; // @[singleLoop.scala 19:20]
  reg [31:0] b_1_2; // @[singleLoop.scala 19:20]
  reg [31:0] b_1_3; // @[singleLoop.scala 19:20]
  reg [31:0] b_1_4; // @[singleLoop.scala 19:20]
  reg [31:0] b_1_5; // @[singleLoop.scala 19:20]
  reg [31:0] b_1_6; // @[singleLoop.scala 19:20]
  reg [31:0] b_1_7; // @[singleLoop.scala 19:20]
  reg [31:0] b_2_0; // @[singleLoop.scala 19:20]
  reg [31:0] b_2_1; // @[singleLoop.scala 19:20]
  reg [31:0] b_2_2; // @[singleLoop.scala 19:20]
  reg [31:0] b_2_3; // @[singleLoop.scala 19:20]
  reg [31:0] b_2_4; // @[singleLoop.scala 19:20]
  reg [31:0] b_2_5; // @[singleLoop.scala 19:20]
  reg [31:0] b_2_6; // @[singleLoop.scala 19:20]
  reg [31:0] b_2_7; // @[singleLoop.scala 19:20]
  reg [31:0] b_3_0; // @[singleLoop.scala 19:20]
  reg [31:0] b_3_1; // @[singleLoop.scala 19:20]
  reg [31:0] b_3_2; // @[singleLoop.scala 19:20]
  reg [31:0] b_3_3; // @[singleLoop.scala 19:20]
  reg [31:0] b_3_4; // @[singleLoop.scala 19:20]
  reg [31:0] b_3_5; // @[singleLoop.scala 19:20]
  reg [31:0] b_3_6; // @[singleLoop.scala 19:20]
  reg [31:0] b_3_7; // @[singleLoop.scala 19:20]
  reg [31:0] b_4_0; // @[singleLoop.scala 19:20]
  reg [31:0] b_4_1; // @[singleLoop.scala 19:20]
  reg [31:0] b_4_2; // @[singleLoop.scala 19:20]
  reg [31:0] b_4_3; // @[singleLoop.scala 19:20]
  reg [31:0] b_4_4; // @[singleLoop.scala 19:20]
  reg [31:0] b_4_5; // @[singleLoop.scala 19:20]
  reg [31:0] b_4_6; // @[singleLoop.scala 19:20]
  reg [31:0] b_4_7; // @[singleLoop.scala 19:20]
  reg [31:0] b_5_0; // @[singleLoop.scala 19:20]
  reg [31:0] b_5_1; // @[singleLoop.scala 19:20]
  reg [31:0] b_5_2; // @[singleLoop.scala 19:20]
  reg [31:0] b_5_3; // @[singleLoop.scala 19:20]
  reg [31:0] b_5_4; // @[singleLoop.scala 19:20]
  reg [31:0] b_5_5; // @[singleLoop.scala 19:20]
  reg [31:0] b_5_6; // @[singleLoop.scala 19:20]
  reg [31:0] b_5_7; // @[singleLoop.scala 19:20]
  reg [31:0] b_6_0; // @[singleLoop.scala 19:20]
  reg [31:0] b_6_1; // @[singleLoop.scala 19:20]
  reg [31:0] b_6_2; // @[singleLoop.scala 19:20]
  reg [31:0] b_6_3; // @[singleLoop.scala 19:20]
  reg [31:0] b_6_4; // @[singleLoop.scala 19:20]
  reg [31:0] b_6_5; // @[singleLoop.scala 19:20]
  reg [31:0] b_6_6; // @[singleLoop.scala 19:20]
  reg [31:0] b_6_7; // @[singleLoop.scala 19:20]
  reg [31:0] b_7_0; // @[singleLoop.scala 19:20]
  reg [31:0] b_7_1; // @[singleLoop.scala 19:20]
  reg [31:0] b_7_2; // @[singleLoop.scala 19:20]
  reg [31:0] b_7_3; // @[singleLoop.scala 19:20]
  reg [31:0] b_7_4; // @[singleLoop.scala 19:20]
  reg [31:0] b_7_5; // @[singleLoop.scala 19:20]
  reg [31:0] b_7_6; // @[singleLoop.scala 19:20]
  reg [31:0] b_7_7; // @[singleLoop.scala 19:20]
  reg [31:0] j; // @[singleLoop.scala 21:16]
  reg [31:0] a; // @[singleLoop.scala 23:20]
  wire  _T_1 = io_valid & a != 32'h0; // @[singleLoop.scala 24:19]
  wire [31:0] _GEN_65 = 3'h0 == io_IDex[2:0] & 3'h1 == j[2:0] ? io_mat_0_1 : io_mat_0_0; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_66 = 3'h0 == io_IDex[2:0] & 3'h2 == j[2:0] ? io_mat_0_2 : _GEN_65; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_67 = 3'h0 == io_IDex[2:0] & 3'h3 == j[2:0] ? io_mat_0_3 : _GEN_66; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_68 = 3'h0 == io_IDex[2:0] & 3'h4 == j[2:0] ? io_mat_0_4 : _GEN_67; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_69 = 3'h0 == io_IDex[2:0] & 3'h5 == j[2:0] ? io_mat_0_5 : _GEN_68; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_70 = 3'h0 == io_IDex[2:0] & 3'h6 == j[2:0] ? io_mat_0_6 : _GEN_69; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_71 = 3'h0 == io_IDex[2:0] & 3'h7 == j[2:0] ? io_mat_0_7 : _GEN_70; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_72 = 3'h1 == io_IDex[2:0] & 3'h0 == j[2:0] ? io_mat_1_0 : _GEN_71; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_73 = 3'h1 == io_IDex[2:0] & 3'h1 == j[2:0] ? io_mat_1_1 : _GEN_72; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_74 = 3'h1 == io_IDex[2:0] & 3'h2 == j[2:0] ? io_mat_1_2 : _GEN_73; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_75 = 3'h1 == io_IDex[2:0] & 3'h3 == j[2:0] ? io_mat_1_3 : _GEN_74; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_76 = 3'h1 == io_IDex[2:0] & 3'h4 == j[2:0] ? io_mat_1_4 : _GEN_75; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_77 = 3'h1 == io_IDex[2:0] & 3'h5 == j[2:0] ? io_mat_1_5 : _GEN_76; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_78 = 3'h1 == io_IDex[2:0] & 3'h6 == j[2:0] ? io_mat_1_6 : _GEN_77; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_79 = 3'h1 == io_IDex[2:0] & 3'h7 == j[2:0] ? io_mat_1_7 : _GEN_78; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_80 = 3'h2 == io_IDex[2:0] & 3'h0 == j[2:0] ? io_mat_2_0 : _GEN_79; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_81 = 3'h2 == io_IDex[2:0] & 3'h1 == j[2:0] ? io_mat_2_1 : _GEN_80; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_82 = 3'h2 == io_IDex[2:0] & 3'h2 == j[2:0] ? io_mat_2_2 : _GEN_81; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_83 = 3'h2 == io_IDex[2:0] & 3'h3 == j[2:0] ? io_mat_2_3 : _GEN_82; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_84 = 3'h2 == io_IDex[2:0] & 3'h4 == j[2:0] ? io_mat_2_4 : _GEN_83; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_85 = 3'h2 == io_IDex[2:0] & 3'h5 == j[2:0] ? io_mat_2_5 : _GEN_84; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_86 = 3'h2 == io_IDex[2:0] & 3'h6 == j[2:0] ? io_mat_2_6 : _GEN_85; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_87 = 3'h2 == io_IDex[2:0] & 3'h7 == j[2:0] ? io_mat_2_7 : _GEN_86; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_88 = 3'h3 == io_IDex[2:0] & 3'h0 == j[2:0] ? io_mat_3_0 : _GEN_87; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_89 = 3'h3 == io_IDex[2:0] & 3'h1 == j[2:0] ? io_mat_3_1 : _GEN_88; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_90 = 3'h3 == io_IDex[2:0] & 3'h2 == j[2:0] ? io_mat_3_2 : _GEN_89; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_91 = 3'h3 == io_IDex[2:0] & 3'h3 == j[2:0] ? io_mat_3_3 : _GEN_90; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_92 = 3'h3 == io_IDex[2:0] & 3'h4 == j[2:0] ? io_mat_3_4 : _GEN_91; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_93 = 3'h3 == io_IDex[2:0] & 3'h5 == j[2:0] ? io_mat_3_5 : _GEN_92; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_94 = 3'h3 == io_IDex[2:0] & 3'h6 == j[2:0] ? io_mat_3_6 : _GEN_93; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_95 = 3'h3 == io_IDex[2:0] & 3'h7 == j[2:0] ? io_mat_3_7 : _GEN_94; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_96 = 3'h4 == io_IDex[2:0] & 3'h0 == j[2:0] ? io_mat_4_0 : _GEN_95; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_97 = 3'h4 == io_IDex[2:0] & 3'h1 == j[2:0] ? io_mat_4_1 : _GEN_96; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_98 = 3'h4 == io_IDex[2:0] & 3'h2 == j[2:0] ? io_mat_4_2 : _GEN_97; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_99 = 3'h4 == io_IDex[2:0] & 3'h3 == j[2:0] ? io_mat_4_3 : _GEN_98; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_100 = 3'h4 == io_IDex[2:0] & 3'h4 == j[2:0] ? io_mat_4_4 : _GEN_99; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_101 = 3'h4 == io_IDex[2:0] & 3'h5 == j[2:0] ? io_mat_4_5 : _GEN_100; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_102 = 3'h4 == io_IDex[2:0] & 3'h6 == j[2:0] ? io_mat_4_6 : _GEN_101; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_103 = 3'h4 == io_IDex[2:0] & 3'h7 == j[2:0] ? io_mat_4_7 : _GEN_102; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_104 = 3'h5 == io_IDex[2:0] & 3'h0 == j[2:0] ? io_mat_5_0 : _GEN_103; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_105 = 3'h5 == io_IDex[2:0] & 3'h1 == j[2:0] ? io_mat_5_1 : _GEN_104; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_106 = 3'h5 == io_IDex[2:0] & 3'h2 == j[2:0] ? io_mat_5_2 : _GEN_105; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_107 = 3'h5 == io_IDex[2:0] & 3'h3 == j[2:0] ? io_mat_5_3 : _GEN_106; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_108 = 3'h5 == io_IDex[2:0] & 3'h4 == j[2:0] ? io_mat_5_4 : _GEN_107; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_109 = 3'h5 == io_IDex[2:0] & 3'h5 == j[2:0] ? io_mat_5_5 : _GEN_108; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_110 = 3'h5 == io_IDex[2:0] & 3'h6 == j[2:0] ? io_mat_5_6 : _GEN_109; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_111 = 3'h5 == io_IDex[2:0] & 3'h7 == j[2:0] ? io_mat_5_7 : _GEN_110; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_112 = 3'h6 == io_IDex[2:0] & 3'h0 == j[2:0] ? io_mat_6_0 : _GEN_111; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_113 = 3'h6 == io_IDex[2:0] & 3'h1 == j[2:0] ? io_mat_6_1 : _GEN_112; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_114 = 3'h6 == io_IDex[2:0] & 3'h2 == j[2:0] ? io_mat_6_2 : _GEN_113; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_115 = 3'h6 == io_IDex[2:0] & 3'h3 == j[2:0] ? io_mat_6_3 : _GEN_114; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_116 = 3'h6 == io_IDex[2:0] & 3'h4 == j[2:0] ? io_mat_6_4 : _GEN_115; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_117 = 3'h6 == io_IDex[2:0] & 3'h5 == j[2:0] ? io_mat_6_5 : _GEN_116; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_118 = 3'h6 == io_IDex[2:0] & 3'h6 == j[2:0] ? io_mat_6_6 : _GEN_117; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_119 = 3'h6 == io_IDex[2:0] & 3'h7 == j[2:0] ? io_mat_6_7 : _GEN_118; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_120 = 3'h7 == io_IDex[2:0] & 3'h0 == j[2:0] ? io_mat_7_0 : _GEN_119; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_121 = 3'h7 == io_IDex[2:0] & 3'h1 == j[2:0] ? io_mat_7_1 : _GEN_120; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_122 = 3'h7 == io_IDex[2:0] & 3'h2 == j[2:0] ? io_mat_7_2 : _GEN_121; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_123 = 3'h7 == io_IDex[2:0] & 3'h3 == j[2:0] ? io_mat_7_3 : _GEN_122; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_124 = 3'h7 == io_IDex[2:0] & 3'h4 == j[2:0] ? io_mat_7_4 : _GEN_123; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_125 = 3'h7 == io_IDex[2:0] & 3'h5 == j[2:0] ? io_mat_7_5 : _GEN_124; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_126 = 3'h7 == io_IDex[2:0] & 3'h6 == j[2:0] ? io_mat_7_6 : _GEN_125; // @[singleLoop.scala 25:{19,19}]
  wire [31:0] _GEN_193 = 3'h1 == io_IDex[2:0] ? io_mat_1_3 : io_mat_0_3; // @[singleLoop.scala 27:{45,45}]
  wire [31:0] _GEN_194 = 3'h2 == io_IDex[2:0] ? io_mat_2_3 : _GEN_193; // @[singleLoop.scala 27:{45,45}]
  wire [31:0] _GEN_195 = 3'h3 == io_IDex[2:0] ? io_mat_3_3 : _GEN_194; // @[singleLoop.scala 27:{45,45}]
  wire [31:0] _GEN_196 = 3'h4 == io_IDex[2:0] ? io_mat_4_3 : _GEN_195; // @[singleLoop.scala 27:{45,45}]
  wire [31:0] _GEN_197 = 3'h5 == io_IDex[2:0] ? io_mat_5_3 : _GEN_196; // @[singleLoop.scala 27:{45,45}]
  wire [31:0] _GEN_198 = 3'h6 == io_IDex[2:0] ? io_mat_6_3 : _GEN_197; // @[singleLoop.scala 27:{45,45}]
  wire [31:0] _GEN_199 = 3'h7 == io_IDex[2:0] ? io_mat_7_3 : _GEN_198; // @[singleLoop.scala 27:{45,45}]
  reg  io_Ovalid_REG; // @[singleLoop.scala 27:25]
  wire  _io_ProcessValid_T = j == 32'h7; // @[singleLoop.scala 31:35]
  wire [31:0] _a_T_1 = a + 32'h1; // @[singleLoop.scala 46:12]
  wire [31:0] _j_T_1 = j + 32'h1; // @[singleLoop.scala 49:16]
  assign io_OutMat_0_0 = b_0_0; // @[singleLoop.scala 20:15]
  assign io_OutMat_0_1 = b_0_1; // @[singleLoop.scala 20:15]
  assign io_OutMat_0_2 = b_0_2; // @[singleLoop.scala 20:15]
  assign io_OutMat_0_3 = b_0_3; // @[singleLoop.scala 20:15]
  assign io_OutMat_0_4 = b_0_4; // @[singleLoop.scala 20:15]
  assign io_OutMat_0_5 = b_0_5; // @[singleLoop.scala 20:15]
  assign io_OutMat_0_6 = b_0_6; // @[singleLoop.scala 20:15]
  assign io_OutMat_0_7 = b_0_7; // @[singleLoop.scala 20:15]
  assign io_OutMat_1_0 = b_1_0; // @[singleLoop.scala 20:15]
  assign io_OutMat_1_1 = b_1_1; // @[singleLoop.scala 20:15]
  assign io_OutMat_1_2 = b_1_2; // @[singleLoop.scala 20:15]
  assign io_OutMat_1_3 = b_1_3; // @[singleLoop.scala 20:15]
  assign io_OutMat_1_4 = b_1_4; // @[singleLoop.scala 20:15]
  assign io_OutMat_1_5 = b_1_5; // @[singleLoop.scala 20:15]
  assign io_OutMat_1_6 = b_1_6; // @[singleLoop.scala 20:15]
  assign io_OutMat_1_7 = b_1_7; // @[singleLoop.scala 20:15]
  assign io_OutMat_2_0 = b_2_0; // @[singleLoop.scala 20:15]
  assign io_OutMat_2_1 = b_2_1; // @[singleLoop.scala 20:15]
  assign io_OutMat_2_2 = b_2_2; // @[singleLoop.scala 20:15]
  assign io_OutMat_2_3 = b_2_3; // @[singleLoop.scala 20:15]
  assign io_OutMat_2_4 = b_2_4; // @[singleLoop.scala 20:15]
  assign io_OutMat_2_5 = b_2_5; // @[singleLoop.scala 20:15]
  assign io_OutMat_2_6 = b_2_6; // @[singleLoop.scala 20:15]
  assign io_OutMat_2_7 = b_2_7; // @[singleLoop.scala 20:15]
  assign io_OutMat_3_0 = b_3_0; // @[singleLoop.scala 20:15]
  assign io_OutMat_3_1 = b_3_1; // @[singleLoop.scala 20:15]
  assign io_OutMat_3_2 = b_3_2; // @[singleLoop.scala 20:15]
  assign io_OutMat_3_3 = b_3_3; // @[singleLoop.scala 20:15]
  assign io_OutMat_3_4 = b_3_4; // @[singleLoop.scala 20:15]
  assign io_OutMat_3_5 = b_3_5; // @[singleLoop.scala 20:15]
  assign io_OutMat_3_6 = b_3_6; // @[singleLoop.scala 20:15]
  assign io_OutMat_3_7 = b_3_7; // @[singleLoop.scala 20:15]
  assign io_OutMat_4_0 = b_4_0; // @[singleLoop.scala 20:15]
  assign io_OutMat_4_1 = b_4_1; // @[singleLoop.scala 20:15]
  assign io_OutMat_4_2 = b_4_2; // @[singleLoop.scala 20:15]
  assign io_OutMat_4_3 = b_4_3; // @[singleLoop.scala 20:15]
  assign io_OutMat_4_4 = b_4_4; // @[singleLoop.scala 20:15]
  assign io_OutMat_4_5 = b_4_5; // @[singleLoop.scala 20:15]
  assign io_OutMat_4_6 = b_4_6; // @[singleLoop.scala 20:15]
  assign io_OutMat_4_7 = b_4_7; // @[singleLoop.scala 20:15]
  assign io_OutMat_5_0 = b_5_0; // @[singleLoop.scala 20:15]
  assign io_OutMat_5_1 = b_5_1; // @[singleLoop.scala 20:15]
  assign io_OutMat_5_2 = b_5_2; // @[singleLoop.scala 20:15]
  assign io_OutMat_5_3 = b_5_3; // @[singleLoop.scala 20:15]
  assign io_OutMat_5_4 = b_5_4; // @[singleLoop.scala 20:15]
  assign io_OutMat_5_5 = b_5_5; // @[singleLoop.scala 20:15]
  assign io_OutMat_5_6 = b_5_6; // @[singleLoop.scala 20:15]
  assign io_OutMat_5_7 = b_5_7; // @[singleLoop.scala 20:15]
  assign io_OutMat_6_0 = b_6_0; // @[singleLoop.scala 20:15]
  assign io_OutMat_6_1 = b_6_1; // @[singleLoop.scala 20:15]
  assign io_OutMat_6_2 = b_6_2; // @[singleLoop.scala 20:15]
  assign io_OutMat_6_3 = b_6_3; // @[singleLoop.scala 20:15]
  assign io_OutMat_6_4 = b_6_4; // @[singleLoop.scala 20:15]
  assign io_OutMat_6_5 = b_6_5; // @[singleLoop.scala 20:15]
  assign io_OutMat_6_6 = b_6_6; // @[singleLoop.scala 20:15]
  assign io_OutMat_6_7 = b_6_7; // @[singleLoop.scala 20:15]
  assign io_OutMat_7_0 = b_7_0; // @[singleLoop.scala 20:15]
  assign io_OutMat_7_1 = b_7_1; // @[singleLoop.scala 20:15]
  assign io_OutMat_7_2 = b_7_2; // @[singleLoop.scala 20:15]
  assign io_OutMat_7_3 = b_7_3; // @[singleLoop.scala 20:15]
  assign io_OutMat_7_4 = b_7_4; // @[singleLoop.scala 20:15]
  assign io_OutMat_7_5 = b_7_5; // @[singleLoop.scala 20:15]
  assign io_OutMat_7_6 = b_7_6; // @[singleLoop.scala 20:15]
  assign io_OutMat_7_7 = b_7_7; // @[singleLoop.scala 20:15]
  assign io_Ovalid = j == 32'h3 & io_Ovalid_REG; // @[singleLoop.scala 26:21 27:15 29:19]
  assign io_ProcessValid = j == 32'h7; // @[singleLoop.scala 31:35]
  always @(posedge clock) begin
    if (reset) begin // @[singleLoop.scala 19:20]
      b_0_0 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h0 == io_IDex[2:0] & 3'h0 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_0_0 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_0_0 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_0_1 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h0 == io_IDex[2:0] & 3'h1 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_0_1 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_0_1 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_0_2 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h0 == io_IDex[2:0] & 3'h2 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_0_2 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_0_2 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_0_3 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h0 == io_IDex[2:0] & 3'h3 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_0_3 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_0_3 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_0_4 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h0 == io_IDex[2:0] & 3'h4 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_0_4 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_0_4 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_0_5 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h0 == io_IDex[2:0] & 3'h5 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_0_5 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_0_5 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_0_6 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h0 == io_IDex[2:0] & 3'h6 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_0_6 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_0_6 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_0_7 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h0 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_0_7 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_0_7 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_1_0 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h1 == io_IDex[2:0] & 3'h0 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_1_0 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_1_0 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_1_1 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h1 == io_IDex[2:0] & 3'h1 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_1_1 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_1_1 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_1_2 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h1 == io_IDex[2:0] & 3'h2 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_1_2 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_1_2 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_1_3 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h1 == io_IDex[2:0] & 3'h3 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_1_3 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_1_3 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_1_4 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h1 == io_IDex[2:0] & 3'h4 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_1_4 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_1_4 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_1_5 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h1 == io_IDex[2:0] & 3'h5 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_1_5 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_1_5 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_1_6 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h1 == io_IDex[2:0] & 3'h6 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_1_6 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_1_6 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_1_7 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h1 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_1_7 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_1_7 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_2_0 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h2 == io_IDex[2:0] & 3'h0 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_2_0 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_2_0 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_2_1 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h2 == io_IDex[2:0] & 3'h1 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_2_1 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_2_1 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_2_2 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h2 == io_IDex[2:0] & 3'h2 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_2_2 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_2_2 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_2_3 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h2 == io_IDex[2:0] & 3'h3 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_2_3 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_2_3 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_2_4 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h2 == io_IDex[2:0] & 3'h4 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_2_4 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_2_4 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_2_5 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h2 == io_IDex[2:0] & 3'h5 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_2_5 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_2_5 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_2_6 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h2 == io_IDex[2:0] & 3'h6 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_2_6 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_2_6 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_2_7 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h2 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_2_7 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_2_7 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_3_0 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h3 == io_IDex[2:0] & 3'h0 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_3_0 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_3_0 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_3_1 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h3 == io_IDex[2:0] & 3'h1 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_3_1 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_3_1 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_3_2 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h3 == io_IDex[2:0] & 3'h2 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_3_2 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_3_2 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_3_3 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h3 == io_IDex[2:0] & 3'h3 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_3_3 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_3_3 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_3_4 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h3 == io_IDex[2:0] & 3'h4 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_3_4 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_3_4 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_3_5 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h3 == io_IDex[2:0] & 3'h5 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_3_5 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_3_5 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_3_6 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h3 == io_IDex[2:0] & 3'h6 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_3_6 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_3_6 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_3_7 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h3 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_3_7 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_3_7 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_4_0 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h4 == io_IDex[2:0] & 3'h0 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_4_0 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_4_0 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_4_1 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h4 == io_IDex[2:0] & 3'h1 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_4_1 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_4_1 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_4_2 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h4 == io_IDex[2:0] & 3'h2 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_4_2 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_4_2 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_4_3 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h4 == io_IDex[2:0] & 3'h3 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_4_3 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_4_3 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_4_4 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h4 == io_IDex[2:0] & 3'h4 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_4_4 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_4_4 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_4_5 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h4 == io_IDex[2:0] & 3'h5 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_4_5 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_4_5 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_4_6 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h4 == io_IDex[2:0] & 3'h6 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_4_6 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_4_6 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_4_7 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h4 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_4_7 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_4_7 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_5_0 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h5 == io_IDex[2:0] & 3'h0 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_5_0 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_5_0 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_5_1 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h5 == io_IDex[2:0] & 3'h1 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_5_1 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_5_1 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_5_2 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h5 == io_IDex[2:0] & 3'h2 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_5_2 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_5_2 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_5_3 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h5 == io_IDex[2:0] & 3'h3 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_5_3 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_5_3 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_5_4 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h5 == io_IDex[2:0] & 3'h4 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_5_4 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_5_4 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_5_5 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h5 == io_IDex[2:0] & 3'h5 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_5_5 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_5_5 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_5_6 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h5 == io_IDex[2:0] & 3'h6 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_5_6 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_5_6 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_5_7 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h5 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_5_7 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_5_7 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_6_0 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h6 == io_IDex[2:0] & 3'h0 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_6_0 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_6_0 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_6_1 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h6 == io_IDex[2:0] & 3'h1 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_6_1 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_6_1 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_6_2 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h6 == io_IDex[2:0] & 3'h2 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_6_2 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_6_2 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_6_3 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h6 == io_IDex[2:0] & 3'h3 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_6_3 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_6_3 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_6_4 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h6 == io_IDex[2:0] & 3'h4 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_6_4 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_6_4 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_6_5 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h6 == io_IDex[2:0] & 3'h5 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_6_5 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_6_5 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_6_6 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h6 == io_IDex[2:0] & 3'h6 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_6_6 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_6_6 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_6_7 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h6 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_6_7 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_6_7 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_7_0 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h7 == io_IDex[2:0] & 3'h0 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_7_0 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_7_0 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_7_1 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h7 == io_IDex[2:0] & 3'h1 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_7_1 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_7_1 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_7_2 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h7 == io_IDex[2:0] & 3'h2 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_7_2 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_7_2 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_7_3 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h7 == io_IDex[2:0] & 3'h3 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_7_3 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_7_3 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_7_4 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h7 == io_IDex[2:0] & 3'h4 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_7_4 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_7_4 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_7_5 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h7 == io_IDex[2:0] & 3'h5 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_7_5 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_7_5 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_7_6 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h7 == io_IDex[2:0] & 3'h6 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_7_6 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_7_6 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[singleLoop.scala 19:20]
      b_7_7 <= 32'h0; // @[singleLoop.scala 19:20]
    end else if (io_valid & a != 32'h0) begin // @[singleLoop.scala 24:34]
      if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[singleLoop.scala 25:19]
          b_7_7 <= io_mat_7_7; // @[singleLoop.scala 25:19]
        end else begin
          b_7_7 <= _GEN_126;
        end
      end
    end
    if (_T_1 & j < 32'h7) begin // @[singleLoop.scala 48:65]
      j <= _j_T_1; // @[singleLoop.scala 49:11]
    end else if (!(_io_ProcessValid_T)) begin // @[singleLoop.scala 50:43]
      j <= io_JDex; // @[singleLoop.scala 22:7]
    end
    if (reset) begin // @[singleLoop.scala 23:20]
      a <= 32'h0; // @[singleLoop.scala 23:20]
    end else if (io_valid) begin // @[singleLoop.scala 45:20]
      a <= _a_T_1; // @[singleLoop.scala 46:7]
    end
    io_Ovalid_REG <= _GEN_199 == 32'h4; // @[singleLoop.scala 27:45]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  b_0_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  b_0_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  b_0_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  b_0_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  b_0_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  b_0_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  b_0_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  b_0_7 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  b_1_0 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  b_1_1 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  b_1_2 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  b_1_3 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  b_1_4 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  b_1_5 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  b_1_6 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  b_1_7 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  b_2_0 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  b_2_1 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  b_2_2 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  b_2_3 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  b_2_4 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  b_2_5 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  b_2_6 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  b_2_7 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  b_3_0 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  b_3_1 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  b_3_2 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  b_3_3 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  b_3_4 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  b_3_5 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  b_3_6 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  b_3_7 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  b_4_0 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  b_4_1 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  b_4_2 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  b_4_3 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  b_4_4 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  b_4_5 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  b_4_6 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  b_4_7 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  b_5_0 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  b_5_1 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  b_5_2 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  b_5_3 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  b_5_4 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  b_5_5 = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  b_5_6 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  b_5_7 = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  b_6_0 = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  b_6_1 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  b_6_2 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  b_6_3 = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  b_6_4 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  b_6_5 = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  b_6_6 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  b_6_7 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  b_7_0 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  b_7_1 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  b_7_2 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  b_7_3 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  b_7_4 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  b_7_5 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  b_7_6 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  b_7_7 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  j = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  a = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  io_Ovalid_REG = _RAND_66[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module abc3(
  input         clock,
  input         reset,
  input  [31:0] io_PreMat_0_0,
  input  [31:0] io_PreMat_0_1,
  input  [31:0] io_PreMat_0_2,
  input  [31:0] io_PreMat_0_3,
  input  [31:0] io_PreMat_0_4,
  input  [31:0] io_PreMat_0_5,
  input  [31:0] io_PreMat_0_6,
  input  [31:0] io_PreMat_0_7,
  input  [31:0] io_PreMat_1_0,
  input  [31:0] io_PreMat_1_1,
  input  [31:0] io_PreMat_1_2,
  input  [31:0] io_PreMat_1_3,
  input  [31:0] io_PreMat_1_4,
  input  [31:0] io_PreMat_1_5,
  input  [31:0] io_PreMat_1_6,
  input  [31:0] io_PreMat_1_7,
  input  [31:0] io_PreMat_2_0,
  input  [31:0] io_PreMat_2_1,
  input  [31:0] io_PreMat_2_2,
  input  [31:0] io_PreMat_2_3,
  input  [31:0] io_PreMat_2_4,
  input  [31:0] io_PreMat_2_5,
  input  [31:0] io_PreMat_2_6,
  input  [31:0] io_PreMat_2_7,
  input  [31:0] io_PreMat_3_0,
  input  [31:0] io_PreMat_3_1,
  input  [31:0] io_PreMat_3_2,
  input  [31:0] io_PreMat_3_3,
  input  [31:0] io_PreMat_3_4,
  input  [31:0] io_PreMat_3_5,
  input  [31:0] io_PreMat_3_6,
  input  [31:0] io_PreMat_3_7,
  input  [31:0] io_PreMat_4_0,
  input  [31:0] io_PreMat_4_1,
  input  [31:0] io_PreMat_4_2,
  input  [31:0] io_PreMat_4_3,
  input  [31:0] io_PreMat_4_4,
  input  [31:0] io_PreMat_4_5,
  input  [31:0] io_PreMat_4_6,
  input  [31:0] io_PreMat_4_7,
  input  [31:0] io_PreMat_5_0,
  input  [31:0] io_PreMat_5_1,
  input  [31:0] io_PreMat_5_2,
  input  [31:0] io_PreMat_5_3,
  input  [31:0] io_PreMat_5_4,
  input  [31:0] io_PreMat_5_5,
  input  [31:0] io_PreMat_5_6,
  input  [31:0] io_PreMat_5_7,
  input  [31:0] io_PreMat_6_0,
  input  [31:0] io_PreMat_6_1,
  input  [31:0] io_PreMat_6_2,
  input  [31:0] io_PreMat_6_3,
  input  [31:0] io_PreMat_6_4,
  input  [31:0] io_PreMat_6_5,
  input  [31:0] io_PreMat_6_6,
  input  [31:0] io_PreMat_6_7,
  input  [31:0] io_PreMat_7_0,
  input  [31:0] io_PreMat_7_1,
  input  [31:0] io_PreMat_7_2,
  input  [31:0] io_PreMat_7_3,
  input  [31:0] io_PreMat_7_4,
  input  [31:0] io_PreMat_7_5,
  input  [31:0] io_PreMat_7_6,
  input  [31:0] io_PreMat_7_7,
  input  [31:0] io_IDex,
  input  [31:0] io_mat_0_0,
  input  [31:0] io_mat_0_1,
  input  [31:0] io_mat_0_2,
  input  [31:0] io_mat_0_3,
  input  [31:0] io_mat_0_4,
  input  [31:0] io_mat_0_5,
  input  [31:0] io_mat_0_6,
  input  [31:0] io_mat_0_7,
  input  [31:0] io_mat_1_0,
  input  [31:0] io_mat_1_1,
  input  [31:0] io_mat_1_2,
  input  [31:0] io_mat_1_3,
  input  [31:0] io_mat_1_4,
  input  [31:0] io_mat_1_5,
  input  [31:0] io_mat_1_6,
  input  [31:0] io_mat_1_7,
  input  [31:0] io_mat_2_0,
  input  [31:0] io_mat_2_1,
  input  [31:0] io_mat_2_2,
  input  [31:0] io_mat_2_3,
  input  [31:0] io_mat_2_4,
  input  [31:0] io_mat_2_5,
  input  [31:0] io_mat_2_6,
  input  [31:0] io_mat_2_7,
  input  [31:0] io_mat_3_0,
  input  [31:0] io_mat_3_1,
  input  [31:0] io_mat_3_2,
  input  [31:0] io_mat_3_3,
  input  [31:0] io_mat_3_4,
  input  [31:0] io_mat_3_5,
  input  [31:0] io_mat_3_6,
  input  [31:0] io_mat_3_7,
  input  [31:0] io_mat_4_0,
  input  [31:0] io_mat_4_1,
  input  [31:0] io_mat_4_2,
  input  [31:0] io_mat_4_3,
  input  [31:0] io_mat_4_4,
  input  [31:0] io_mat_4_5,
  input  [31:0] io_mat_4_6,
  input  [31:0] io_mat_4_7,
  input  [31:0] io_mat_5_0,
  input  [31:0] io_mat_5_1,
  input  [31:0] io_mat_5_2,
  input  [31:0] io_mat_5_3,
  input  [31:0] io_mat_5_4,
  input  [31:0] io_mat_5_5,
  input  [31:0] io_mat_5_6,
  input  [31:0] io_mat_5_7,
  input  [31:0] io_mat_6_0,
  input  [31:0] io_mat_6_1,
  input  [31:0] io_mat_6_2,
  input  [31:0] io_mat_6_3,
  input  [31:0] io_mat_6_4,
  input  [31:0] io_mat_6_5,
  input  [31:0] io_mat_6_6,
  input  [31:0] io_mat_6_7,
  input  [31:0] io_mat_7_0,
  input  [31:0] io_mat_7_1,
  input  [31:0] io_mat_7_2,
  input  [31:0] io_mat_7_3,
  input  [31:0] io_mat_7_4,
  input  [31:0] io_mat_7_5,
  input  [31:0] io_mat_7_6,
  input  [31:0] io_mat_7_7,
  input         io_i_valid,
  output        io_valid,
  output [31:0] io_Omat_0_0,
  output [31:0] io_Omat_0_1,
  output [31:0] io_Omat_0_2,
  output [31:0] io_Omat_0_3,
  output [31:0] io_Omat_0_4,
  output [31:0] io_Omat_0_5,
  output [31:0] io_Omat_0_6,
  output [31:0] io_Omat_0_7,
  output [31:0] io_Omat_1_0,
  output [31:0] io_Omat_1_1,
  output [31:0] io_Omat_1_2,
  output [31:0] io_Omat_1_3,
  output [31:0] io_Omat_1_4,
  output [31:0] io_Omat_1_5,
  output [31:0] io_Omat_1_6,
  output [31:0] io_Omat_1_7,
  output [31:0] io_Omat_2_0,
  output [31:0] io_Omat_2_1,
  output [31:0] io_Omat_2_2,
  output [31:0] io_Omat_2_3,
  output [31:0] io_Omat_2_4,
  output [31:0] io_Omat_2_5,
  output [31:0] io_Omat_2_6,
  output [31:0] io_Omat_2_7,
  output [31:0] io_Omat_3_0,
  output [31:0] io_Omat_3_1,
  output [31:0] io_Omat_3_2,
  output [31:0] io_Omat_3_3,
  output [31:0] io_Omat_3_4,
  output [31:0] io_Omat_3_5,
  output [31:0] io_Omat_3_6,
  output [31:0] io_Omat_3_7,
  output [31:0] io_Omat_4_0,
  output [31:0] io_Omat_4_1,
  output [31:0] io_Omat_4_2,
  output [31:0] io_Omat_4_3,
  output [31:0] io_Omat_4_4,
  output [31:0] io_Omat_4_5,
  output [31:0] io_Omat_4_6,
  output [31:0] io_Omat_4_7,
  output [31:0] io_Omat_5_0,
  output [31:0] io_Omat_5_1,
  output [31:0] io_Omat_5_2,
  output [31:0] io_Omat_5_3,
  output [31:0] io_Omat_5_4,
  output [31:0] io_Omat_5_5,
  output [31:0] io_Omat_5_6,
  output [31:0] io_Omat_5_7,
  output [31:0] io_Omat_6_0,
  output [31:0] io_Omat_6_1,
  output [31:0] io_Omat_6_2,
  output [31:0] io_Omat_6_3,
  output [31:0] io_Omat_6_4,
  output [31:0] io_Omat_6_5,
  output [31:0] io_Omat_6_6,
  output [31:0] io_Omat_6_7,
  output [31:0] io_Omat_7_0,
  output [31:0] io_Omat_7_1,
  output [31:0] io_Omat_7_2,
  output [31:0] io_Omat_7_3,
  output [31:0] io_Omat_7_4,
  output [31:0] io_Omat_7_5,
  output [31:0] io_Omat_7_6,
  output [31:0] io_Omat_7_7,
  input         io_merge
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] b_0_0; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_0_1; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_0_2; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_0_3; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_0_4; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_0_5; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_0_6; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_0_7; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_1_0; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_1_1; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_1_2; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_1_3; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_1_4; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_1_5; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_1_6; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_1_7; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_2_0; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_2_1; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_2_2; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_2_3; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_2_4; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_2_5; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_2_6; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_2_7; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_3_0; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_3_1; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_3_2; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_3_3; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_3_4; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_3_5; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_3_6; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_3_7; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_4_0; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_4_1; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_4_2; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_4_3; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_4_4; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_4_5; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_4_6; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_4_7; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_5_0; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_5_1; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_5_2; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_5_3; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_5_4; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_5_5; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_5_6; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_5_7; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_6_0; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_6_1; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_6_2; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_6_3; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_6_4; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_6_5; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_6_6; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_6_7; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_7_0; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_7_1; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_7_2; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_7_3; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_7_4; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_7_5; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_7_6; // @[MergeDIstribution.scala 18:20]
  reg [31:0] b_7_7; // @[MergeDIstribution.scala 18:20]
  reg [31:0] check; // @[MergeDIstribution.scala 20:24]
  reg [31:0] i; // @[MergeDIstribution.scala 22:20]
  reg [31:0] j; // @[MergeDIstribution.scala 23:20]
  reg [31:0] k; // @[MergeDIstribution.scala 26:20]
  reg [31:0] l; // @[MergeDIstribution.scala 27:20]
  reg [31:0] delay; // @[MergeDIstribution.scala 29:24]
  wire [31:0] _delay_T_1 = delay + 32'h1; // @[MergeDIstribution.scala 32:24]
  wire [31:0] _k_T_1 = k + 32'h1; // @[MergeDIstribution.scala 44:16]
  wire [31:0] _l_T_1 = l + 32'h1; // @[MergeDIstribution.scala 47:16]
  wire [31:0] _GEN_70 = 3'h0 == k[2:0] & 3'h1 == l[2:0] ? io_PreMat_0_1 : io_PreMat_0_0; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_71 = 3'h0 == k[2:0] & 3'h2 == l[2:0] ? io_PreMat_0_2 : _GEN_70; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_72 = 3'h0 == k[2:0] & 3'h3 == l[2:0] ? io_PreMat_0_3 : _GEN_71; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_73 = 3'h0 == k[2:0] & 3'h4 == l[2:0] ? io_PreMat_0_4 : _GEN_72; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_74 = 3'h0 == k[2:0] & 3'h5 == l[2:0] ? io_PreMat_0_5 : _GEN_73; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_75 = 3'h0 == k[2:0] & 3'h6 == l[2:0] ? io_PreMat_0_6 : _GEN_74; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_76 = 3'h0 == k[2:0] & 3'h7 == l[2:0] ? io_PreMat_0_7 : _GEN_75; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_77 = 3'h1 == k[2:0] & 3'h0 == l[2:0] ? io_PreMat_1_0 : _GEN_76; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_78 = 3'h1 == k[2:0] & 3'h1 == l[2:0] ? io_PreMat_1_1 : _GEN_77; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_79 = 3'h1 == k[2:0] & 3'h2 == l[2:0] ? io_PreMat_1_2 : _GEN_78; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_80 = 3'h1 == k[2:0] & 3'h3 == l[2:0] ? io_PreMat_1_3 : _GEN_79; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_81 = 3'h1 == k[2:0] & 3'h4 == l[2:0] ? io_PreMat_1_4 : _GEN_80; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_82 = 3'h1 == k[2:0] & 3'h5 == l[2:0] ? io_PreMat_1_5 : _GEN_81; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_83 = 3'h1 == k[2:0] & 3'h6 == l[2:0] ? io_PreMat_1_6 : _GEN_82; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_84 = 3'h1 == k[2:0] & 3'h7 == l[2:0] ? io_PreMat_1_7 : _GEN_83; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_85 = 3'h2 == k[2:0] & 3'h0 == l[2:0] ? io_PreMat_2_0 : _GEN_84; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_86 = 3'h2 == k[2:0] & 3'h1 == l[2:0] ? io_PreMat_2_1 : _GEN_85; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_87 = 3'h2 == k[2:0] & 3'h2 == l[2:0] ? io_PreMat_2_2 : _GEN_86; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_88 = 3'h2 == k[2:0] & 3'h3 == l[2:0] ? io_PreMat_2_3 : _GEN_87; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_89 = 3'h2 == k[2:0] & 3'h4 == l[2:0] ? io_PreMat_2_4 : _GEN_88; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_90 = 3'h2 == k[2:0] & 3'h5 == l[2:0] ? io_PreMat_2_5 : _GEN_89; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_91 = 3'h2 == k[2:0] & 3'h6 == l[2:0] ? io_PreMat_2_6 : _GEN_90; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_92 = 3'h2 == k[2:0] & 3'h7 == l[2:0] ? io_PreMat_2_7 : _GEN_91; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_93 = 3'h3 == k[2:0] & 3'h0 == l[2:0] ? io_PreMat_3_0 : _GEN_92; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_94 = 3'h3 == k[2:0] & 3'h1 == l[2:0] ? io_PreMat_3_1 : _GEN_93; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_95 = 3'h3 == k[2:0] & 3'h2 == l[2:0] ? io_PreMat_3_2 : _GEN_94; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_96 = 3'h3 == k[2:0] & 3'h3 == l[2:0] ? io_PreMat_3_3 : _GEN_95; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_97 = 3'h3 == k[2:0] & 3'h4 == l[2:0] ? io_PreMat_3_4 : _GEN_96; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_98 = 3'h3 == k[2:0] & 3'h5 == l[2:0] ? io_PreMat_3_5 : _GEN_97; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_99 = 3'h3 == k[2:0] & 3'h6 == l[2:0] ? io_PreMat_3_6 : _GEN_98; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_100 = 3'h3 == k[2:0] & 3'h7 == l[2:0] ? io_PreMat_3_7 : _GEN_99; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_101 = 3'h4 == k[2:0] & 3'h0 == l[2:0] ? io_PreMat_4_0 : _GEN_100; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_102 = 3'h4 == k[2:0] & 3'h1 == l[2:0] ? io_PreMat_4_1 : _GEN_101; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_103 = 3'h4 == k[2:0] & 3'h2 == l[2:0] ? io_PreMat_4_2 : _GEN_102; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_104 = 3'h4 == k[2:0] & 3'h3 == l[2:0] ? io_PreMat_4_3 : _GEN_103; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_105 = 3'h4 == k[2:0] & 3'h4 == l[2:0] ? io_PreMat_4_4 : _GEN_104; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_106 = 3'h4 == k[2:0] & 3'h5 == l[2:0] ? io_PreMat_4_5 : _GEN_105; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_107 = 3'h4 == k[2:0] & 3'h6 == l[2:0] ? io_PreMat_4_6 : _GEN_106; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_108 = 3'h4 == k[2:0] & 3'h7 == l[2:0] ? io_PreMat_4_7 : _GEN_107; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_109 = 3'h5 == k[2:0] & 3'h0 == l[2:0] ? io_PreMat_5_0 : _GEN_108; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_110 = 3'h5 == k[2:0] & 3'h1 == l[2:0] ? io_PreMat_5_1 : _GEN_109; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_111 = 3'h5 == k[2:0] & 3'h2 == l[2:0] ? io_PreMat_5_2 : _GEN_110; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_112 = 3'h5 == k[2:0] & 3'h3 == l[2:0] ? io_PreMat_5_3 : _GEN_111; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_113 = 3'h5 == k[2:0] & 3'h4 == l[2:0] ? io_PreMat_5_4 : _GEN_112; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_114 = 3'h5 == k[2:0] & 3'h5 == l[2:0] ? io_PreMat_5_5 : _GEN_113; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_115 = 3'h5 == k[2:0] & 3'h6 == l[2:0] ? io_PreMat_5_6 : _GEN_114; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_116 = 3'h5 == k[2:0] & 3'h7 == l[2:0] ? io_PreMat_5_7 : _GEN_115; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_117 = 3'h6 == k[2:0] & 3'h0 == l[2:0] ? io_PreMat_6_0 : _GEN_116; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_118 = 3'h6 == k[2:0] & 3'h1 == l[2:0] ? io_PreMat_6_1 : _GEN_117; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_119 = 3'h6 == k[2:0] & 3'h2 == l[2:0] ? io_PreMat_6_2 : _GEN_118; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_120 = 3'h6 == k[2:0] & 3'h3 == l[2:0] ? io_PreMat_6_3 : _GEN_119; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_121 = 3'h6 == k[2:0] & 3'h4 == l[2:0] ? io_PreMat_6_4 : _GEN_120; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_122 = 3'h6 == k[2:0] & 3'h5 == l[2:0] ? io_PreMat_6_5 : _GEN_121; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_123 = 3'h6 == k[2:0] & 3'h6 == l[2:0] ? io_PreMat_6_6 : _GEN_122; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_124 = 3'h6 == k[2:0] & 3'h7 == l[2:0] ? io_PreMat_6_7 : _GEN_123; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_125 = 3'h7 == k[2:0] & 3'h0 == l[2:0] ? io_PreMat_7_0 : _GEN_124; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_126 = 3'h7 == k[2:0] & 3'h1 == l[2:0] ? io_PreMat_7_1 : _GEN_125; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_127 = 3'h7 == k[2:0] & 3'h2 == l[2:0] ? io_PreMat_7_2 : _GEN_126; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_128 = 3'h7 == k[2:0] & 3'h3 == l[2:0] ? io_PreMat_7_3 : _GEN_127; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_129 = 3'h7 == k[2:0] & 3'h4 == l[2:0] ? io_PreMat_7_4 : _GEN_128; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_130 = 3'h7 == k[2:0] & 3'h5 == l[2:0] ? io_PreMat_7_5 : _GEN_129; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_131 = 3'h7 == k[2:0] & 3'h6 == l[2:0] ? io_PreMat_7_6 : _GEN_130; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_132 = 3'h7 == k[2:0] & 3'h7 == l[2:0] ? io_PreMat_7_7 : _GEN_131; // @[MergeDIstribution.scala 52:{13,13}]
  wire [31:0] _GEN_5 = 3'h0 == k[2:0] & 3'h0 == l[2:0] ? _GEN_132 : b_0_0; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_6 = 3'h0 == k[2:0] & 3'h1 == l[2:0] ? _GEN_132 : b_0_1; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_7 = 3'h0 == k[2:0] & 3'h2 == l[2:0] ? _GEN_132 : b_0_2; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_8 = 3'h0 == k[2:0] & 3'h3 == l[2:0] ? _GEN_132 : b_0_3; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_9 = 3'h0 == k[2:0] & 3'h4 == l[2:0] ? _GEN_132 : b_0_4; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_10 = 3'h0 == k[2:0] & 3'h5 == l[2:0] ? _GEN_132 : b_0_5; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_11 = 3'h0 == k[2:0] & 3'h6 == l[2:0] ? _GEN_132 : b_0_6; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_12 = 3'h0 == k[2:0] & 3'h7 == l[2:0] ? _GEN_132 : b_0_7; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_13 = 3'h1 == k[2:0] & 3'h0 == l[2:0] ? _GEN_132 : b_1_0; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_14 = 3'h1 == k[2:0] & 3'h1 == l[2:0] ? _GEN_132 : b_1_1; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_15 = 3'h1 == k[2:0] & 3'h2 == l[2:0] ? _GEN_132 : b_1_2; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_16 = 3'h1 == k[2:0] & 3'h3 == l[2:0] ? _GEN_132 : b_1_3; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_17 = 3'h1 == k[2:0] & 3'h4 == l[2:0] ? _GEN_132 : b_1_4; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_18 = 3'h1 == k[2:0] & 3'h5 == l[2:0] ? _GEN_132 : b_1_5; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_19 = 3'h1 == k[2:0] & 3'h6 == l[2:0] ? _GEN_132 : b_1_6; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_20 = 3'h1 == k[2:0] & 3'h7 == l[2:0] ? _GEN_132 : b_1_7; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_21 = 3'h2 == k[2:0] & 3'h0 == l[2:0] ? _GEN_132 : b_2_0; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_22 = 3'h2 == k[2:0] & 3'h1 == l[2:0] ? _GEN_132 : b_2_1; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_23 = 3'h2 == k[2:0] & 3'h2 == l[2:0] ? _GEN_132 : b_2_2; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_24 = 3'h2 == k[2:0] & 3'h3 == l[2:0] ? _GEN_132 : b_2_3; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_25 = 3'h2 == k[2:0] & 3'h4 == l[2:0] ? _GEN_132 : b_2_4; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_26 = 3'h2 == k[2:0] & 3'h5 == l[2:0] ? _GEN_132 : b_2_5; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_27 = 3'h2 == k[2:0] & 3'h6 == l[2:0] ? _GEN_132 : b_2_6; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_28 = 3'h2 == k[2:0] & 3'h7 == l[2:0] ? _GEN_132 : b_2_7; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_29 = 3'h3 == k[2:0] & 3'h0 == l[2:0] ? _GEN_132 : b_3_0; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_30 = 3'h3 == k[2:0] & 3'h1 == l[2:0] ? _GEN_132 : b_3_1; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_31 = 3'h3 == k[2:0] & 3'h2 == l[2:0] ? _GEN_132 : b_3_2; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_32 = 3'h3 == k[2:0] & 3'h3 == l[2:0] ? _GEN_132 : b_3_3; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_33 = 3'h3 == k[2:0] & 3'h4 == l[2:0] ? _GEN_132 : b_3_4; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_34 = 3'h3 == k[2:0] & 3'h5 == l[2:0] ? _GEN_132 : b_3_5; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_35 = 3'h3 == k[2:0] & 3'h6 == l[2:0] ? _GEN_132 : b_3_6; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_36 = 3'h3 == k[2:0] & 3'h7 == l[2:0] ? _GEN_132 : b_3_7; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_37 = 3'h4 == k[2:0] & 3'h0 == l[2:0] ? _GEN_132 : b_4_0; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_38 = 3'h4 == k[2:0] & 3'h1 == l[2:0] ? _GEN_132 : b_4_1; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_39 = 3'h4 == k[2:0] & 3'h2 == l[2:0] ? _GEN_132 : b_4_2; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_40 = 3'h4 == k[2:0] & 3'h3 == l[2:0] ? _GEN_132 : b_4_3; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_41 = 3'h4 == k[2:0] & 3'h4 == l[2:0] ? _GEN_132 : b_4_4; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_42 = 3'h4 == k[2:0] & 3'h5 == l[2:0] ? _GEN_132 : b_4_5; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_43 = 3'h4 == k[2:0] & 3'h6 == l[2:0] ? _GEN_132 : b_4_6; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_44 = 3'h4 == k[2:0] & 3'h7 == l[2:0] ? _GEN_132 : b_4_7; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_45 = 3'h5 == k[2:0] & 3'h0 == l[2:0] ? _GEN_132 : b_5_0; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_46 = 3'h5 == k[2:0] & 3'h1 == l[2:0] ? _GEN_132 : b_5_1; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_47 = 3'h5 == k[2:0] & 3'h2 == l[2:0] ? _GEN_132 : b_5_2; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_48 = 3'h5 == k[2:0] & 3'h3 == l[2:0] ? _GEN_132 : b_5_3; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_49 = 3'h5 == k[2:0] & 3'h4 == l[2:0] ? _GEN_132 : b_5_4; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_50 = 3'h5 == k[2:0] & 3'h5 == l[2:0] ? _GEN_132 : b_5_5; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_51 = 3'h5 == k[2:0] & 3'h6 == l[2:0] ? _GEN_132 : b_5_6; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_52 = 3'h5 == k[2:0] & 3'h7 == l[2:0] ? _GEN_132 : b_5_7; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_53 = 3'h6 == k[2:0] & 3'h0 == l[2:0] ? _GEN_132 : b_6_0; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_54 = 3'h6 == k[2:0] & 3'h1 == l[2:0] ? _GEN_132 : b_6_1; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_55 = 3'h6 == k[2:0] & 3'h2 == l[2:0] ? _GEN_132 : b_6_2; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_56 = 3'h6 == k[2:0] & 3'h3 == l[2:0] ? _GEN_132 : b_6_3; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_57 = 3'h6 == k[2:0] & 3'h4 == l[2:0] ? _GEN_132 : b_6_4; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_58 = 3'h6 == k[2:0] & 3'h5 == l[2:0] ? _GEN_132 : b_6_5; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_59 = 3'h6 == k[2:0] & 3'h6 == l[2:0] ? _GEN_132 : b_6_6; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_60 = 3'h6 == k[2:0] & 3'h7 == l[2:0] ? _GEN_132 : b_6_7; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_61 = 3'h7 == k[2:0] & 3'h0 == l[2:0] ? _GEN_132 : b_7_0; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_62 = 3'h7 == k[2:0] & 3'h1 == l[2:0] ? _GEN_132 : b_7_1; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_63 = 3'h7 == k[2:0] & 3'h2 == l[2:0] ? _GEN_132 : b_7_2; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_64 = 3'h7 == k[2:0] & 3'h3 == l[2:0] ? _GEN_132 : b_7_3; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_65 = 3'h7 == k[2:0] & 3'h4 == l[2:0] ? _GEN_132 : b_7_4; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_66 = 3'h7 == k[2:0] & 3'h5 == l[2:0] ? _GEN_132 : b_7_5; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_67 = 3'h7 == k[2:0] & 3'h6 == l[2:0] ? _GEN_132 : b_7_6; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_68 = 3'h7 == k[2:0] & 3'h7 == l[2:0] ? _GEN_132 : b_7_7; // @[MergeDIstribution.scala 52:{13,13} 18:20]
  wire [31:0] _GEN_135 = io_merge & delay == 32'h8 ? _GEN_5 : b_0_0; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_136 = io_merge & delay == 32'h8 ? _GEN_6 : b_0_1; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_137 = io_merge & delay == 32'h8 ? _GEN_7 : b_0_2; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_138 = io_merge & delay == 32'h8 ? _GEN_8 : b_0_3; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_139 = io_merge & delay == 32'h8 ? _GEN_9 : b_0_4; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_140 = io_merge & delay == 32'h8 ? _GEN_10 : b_0_5; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_141 = io_merge & delay == 32'h8 ? _GEN_11 : b_0_6; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_142 = io_merge & delay == 32'h8 ? _GEN_12 : b_0_7; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_143 = io_merge & delay == 32'h8 ? _GEN_13 : b_1_0; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_144 = io_merge & delay == 32'h8 ? _GEN_14 : b_1_1; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_145 = io_merge & delay == 32'h8 ? _GEN_15 : b_1_2; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_146 = io_merge & delay == 32'h8 ? _GEN_16 : b_1_3; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_147 = io_merge & delay == 32'h8 ? _GEN_17 : b_1_4; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_148 = io_merge & delay == 32'h8 ? _GEN_18 : b_1_5; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_149 = io_merge & delay == 32'h8 ? _GEN_19 : b_1_6; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_150 = io_merge & delay == 32'h8 ? _GEN_20 : b_1_7; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_151 = io_merge & delay == 32'h8 ? _GEN_21 : b_2_0; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_152 = io_merge & delay == 32'h8 ? _GEN_22 : b_2_1; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_153 = io_merge & delay == 32'h8 ? _GEN_23 : b_2_2; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_154 = io_merge & delay == 32'h8 ? _GEN_24 : b_2_3; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_155 = io_merge & delay == 32'h8 ? _GEN_25 : b_2_4; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_156 = io_merge & delay == 32'h8 ? _GEN_26 : b_2_5; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_157 = io_merge & delay == 32'h8 ? _GEN_27 : b_2_6; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_158 = io_merge & delay == 32'h8 ? _GEN_28 : b_2_7; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_159 = io_merge & delay == 32'h8 ? _GEN_29 : b_3_0; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_160 = io_merge & delay == 32'h8 ? _GEN_30 : b_3_1; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_161 = io_merge & delay == 32'h8 ? _GEN_31 : b_3_2; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_162 = io_merge & delay == 32'h8 ? _GEN_32 : b_3_3; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_163 = io_merge & delay == 32'h8 ? _GEN_33 : b_3_4; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_164 = io_merge & delay == 32'h8 ? _GEN_34 : b_3_5; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_165 = io_merge & delay == 32'h8 ? _GEN_35 : b_3_6; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_166 = io_merge & delay == 32'h8 ? _GEN_36 : b_3_7; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_167 = io_merge & delay == 32'h8 ? _GEN_37 : b_4_0; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_168 = io_merge & delay == 32'h8 ? _GEN_38 : b_4_1; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_169 = io_merge & delay == 32'h8 ? _GEN_39 : b_4_2; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_170 = io_merge & delay == 32'h8 ? _GEN_40 : b_4_3; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_171 = io_merge & delay == 32'h8 ? _GEN_41 : b_4_4; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_172 = io_merge & delay == 32'h8 ? _GEN_42 : b_4_5; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_173 = io_merge & delay == 32'h8 ? _GEN_43 : b_4_6; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_174 = io_merge & delay == 32'h8 ? _GEN_44 : b_4_7; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_175 = io_merge & delay == 32'h8 ? _GEN_45 : b_5_0; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_176 = io_merge & delay == 32'h8 ? _GEN_46 : b_5_1; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_177 = io_merge & delay == 32'h8 ? _GEN_47 : b_5_2; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_178 = io_merge & delay == 32'h8 ? _GEN_48 : b_5_3; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_179 = io_merge & delay == 32'h8 ? _GEN_49 : b_5_4; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_180 = io_merge & delay == 32'h8 ? _GEN_50 : b_5_5; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_181 = io_merge & delay == 32'h8 ? _GEN_51 : b_5_6; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_182 = io_merge & delay == 32'h8 ? _GEN_52 : b_5_7; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_183 = io_merge & delay == 32'h8 ? _GEN_53 : b_6_0; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_184 = io_merge & delay == 32'h8 ? _GEN_54 : b_6_1; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_185 = io_merge & delay == 32'h8 ? _GEN_55 : b_6_2; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_186 = io_merge & delay == 32'h8 ? _GEN_56 : b_6_3; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_187 = io_merge & delay == 32'h8 ? _GEN_57 : b_6_4; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_188 = io_merge & delay == 32'h8 ? _GEN_58 : b_6_5; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_189 = io_merge & delay == 32'h8 ? _GEN_59 : b_6_6; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_190 = io_merge & delay == 32'h8 ? _GEN_60 : b_6_7; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_191 = io_merge & delay == 32'h8 ? _GEN_61 : b_7_0; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_192 = io_merge & delay == 32'h8 ? _GEN_62 : b_7_1; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_193 = io_merge & delay == 32'h8 ? _GEN_63 : b_7_2; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_194 = io_merge & delay == 32'h8 ? _GEN_64 : b_7_3; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_195 = io_merge & delay == 32'h8 ? _GEN_65 : b_7_4; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_196 = io_merge & delay == 32'h8 ? _GEN_66 : b_7_5; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_197 = io_merge & delay == 32'h8 ? _GEN_67 : b_7_6; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _GEN_198 = io_merge & delay == 32'h8 ? _GEN_68 : b_7_7; // @[MergeDIstribution.scala 18:20 41:53]
  wire [31:0] _i_T_1 = io_IDex + 32'h1; // @[MergeDIstribution.scala 55:22]
  wire [31:0] _check_T_1 = check + 32'h1; // @[MergeDIstribution.scala 57:24]
  wire [31:0] _GEN_199 = io_i_valid & i == 32'h0 & j == 32'h0 ? _i_T_1 : i; // @[MergeDIstribution.scala 54:53 55:11 22:20]
  wire [31:0] _GEN_200 = io_i_valid & i == 32'h0 & j == 32'h0 ? 32'h0 : j; // @[MergeDIstribution.scala 54:53 56:11 23:20]
  wire  _GEN_202 = check >= 32'h1; // @[MergeDIstribution.scala 60:17]
  wire [31:0] _GEN_269 = 3'h0 == i[2:0] & 3'h1 == j[2:0] ? io_mat_0_1 : io_mat_0_0; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_270 = 3'h0 == i[2:0] & 3'h2 == j[2:0] ? io_mat_0_2 : _GEN_269; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_271 = 3'h0 == i[2:0] & 3'h3 == j[2:0] ? io_mat_0_3 : _GEN_270; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_272 = 3'h0 == i[2:0] & 3'h4 == j[2:0] ? io_mat_0_4 : _GEN_271; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_273 = 3'h0 == i[2:0] & 3'h5 == j[2:0] ? io_mat_0_5 : _GEN_272; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_274 = 3'h0 == i[2:0] & 3'h6 == j[2:0] ? io_mat_0_6 : _GEN_273; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_275 = 3'h0 == i[2:0] & 3'h7 == j[2:0] ? io_mat_0_7 : _GEN_274; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_276 = 3'h1 == i[2:0] & 3'h0 == j[2:0] ? io_mat_1_0 : _GEN_275; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_277 = 3'h1 == i[2:0] & 3'h1 == j[2:0] ? io_mat_1_1 : _GEN_276; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_278 = 3'h1 == i[2:0] & 3'h2 == j[2:0] ? io_mat_1_2 : _GEN_277; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_279 = 3'h1 == i[2:0] & 3'h3 == j[2:0] ? io_mat_1_3 : _GEN_278; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_280 = 3'h1 == i[2:0] & 3'h4 == j[2:0] ? io_mat_1_4 : _GEN_279; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_281 = 3'h1 == i[2:0] & 3'h5 == j[2:0] ? io_mat_1_5 : _GEN_280; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_282 = 3'h1 == i[2:0] & 3'h6 == j[2:0] ? io_mat_1_6 : _GEN_281; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_283 = 3'h1 == i[2:0] & 3'h7 == j[2:0] ? io_mat_1_7 : _GEN_282; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_284 = 3'h2 == i[2:0] & 3'h0 == j[2:0] ? io_mat_2_0 : _GEN_283; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_285 = 3'h2 == i[2:0] & 3'h1 == j[2:0] ? io_mat_2_1 : _GEN_284; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_286 = 3'h2 == i[2:0] & 3'h2 == j[2:0] ? io_mat_2_2 : _GEN_285; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_287 = 3'h2 == i[2:0] & 3'h3 == j[2:0] ? io_mat_2_3 : _GEN_286; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_288 = 3'h2 == i[2:0] & 3'h4 == j[2:0] ? io_mat_2_4 : _GEN_287; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_289 = 3'h2 == i[2:0] & 3'h5 == j[2:0] ? io_mat_2_5 : _GEN_288; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_290 = 3'h2 == i[2:0] & 3'h6 == j[2:0] ? io_mat_2_6 : _GEN_289; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_291 = 3'h2 == i[2:0] & 3'h7 == j[2:0] ? io_mat_2_7 : _GEN_290; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_292 = 3'h3 == i[2:0] & 3'h0 == j[2:0] ? io_mat_3_0 : _GEN_291; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_293 = 3'h3 == i[2:0] & 3'h1 == j[2:0] ? io_mat_3_1 : _GEN_292; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_294 = 3'h3 == i[2:0] & 3'h2 == j[2:0] ? io_mat_3_2 : _GEN_293; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_295 = 3'h3 == i[2:0] & 3'h3 == j[2:0] ? io_mat_3_3 : _GEN_294; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_296 = 3'h3 == i[2:0] & 3'h4 == j[2:0] ? io_mat_3_4 : _GEN_295; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_297 = 3'h3 == i[2:0] & 3'h5 == j[2:0] ? io_mat_3_5 : _GEN_296; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_298 = 3'h3 == i[2:0] & 3'h6 == j[2:0] ? io_mat_3_6 : _GEN_297; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_299 = 3'h3 == i[2:0] & 3'h7 == j[2:0] ? io_mat_3_7 : _GEN_298; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_300 = 3'h4 == i[2:0] & 3'h0 == j[2:0] ? io_mat_4_0 : _GEN_299; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_301 = 3'h4 == i[2:0] & 3'h1 == j[2:0] ? io_mat_4_1 : _GEN_300; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_302 = 3'h4 == i[2:0] & 3'h2 == j[2:0] ? io_mat_4_2 : _GEN_301; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_303 = 3'h4 == i[2:0] & 3'h3 == j[2:0] ? io_mat_4_3 : _GEN_302; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_304 = 3'h4 == i[2:0] & 3'h4 == j[2:0] ? io_mat_4_4 : _GEN_303; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_305 = 3'h4 == i[2:0] & 3'h5 == j[2:0] ? io_mat_4_5 : _GEN_304; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_306 = 3'h4 == i[2:0] & 3'h6 == j[2:0] ? io_mat_4_6 : _GEN_305; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_307 = 3'h4 == i[2:0] & 3'h7 == j[2:0] ? io_mat_4_7 : _GEN_306; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_308 = 3'h5 == i[2:0] & 3'h0 == j[2:0] ? io_mat_5_0 : _GEN_307; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_309 = 3'h5 == i[2:0] & 3'h1 == j[2:0] ? io_mat_5_1 : _GEN_308; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_310 = 3'h5 == i[2:0] & 3'h2 == j[2:0] ? io_mat_5_2 : _GEN_309; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_311 = 3'h5 == i[2:0] & 3'h3 == j[2:0] ? io_mat_5_3 : _GEN_310; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_312 = 3'h5 == i[2:0] & 3'h4 == j[2:0] ? io_mat_5_4 : _GEN_311; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_313 = 3'h5 == i[2:0] & 3'h5 == j[2:0] ? io_mat_5_5 : _GEN_312; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_314 = 3'h5 == i[2:0] & 3'h6 == j[2:0] ? io_mat_5_6 : _GEN_313; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_315 = 3'h5 == i[2:0] & 3'h7 == j[2:0] ? io_mat_5_7 : _GEN_314; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_316 = 3'h6 == i[2:0] & 3'h0 == j[2:0] ? io_mat_6_0 : _GEN_315; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_317 = 3'h6 == i[2:0] & 3'h1 == j[2:0] ? io_mat_6_1 : _GEN_316; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_318 = 3'h6 == i[2:0] & 3'h2 == j[2:0] ? io_mat_6_2 : _GEN_317; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_319 = 3'h6 == i[2:0] & 3'h3 == j[2:0] ? io_mat_6_3 : _GEN_318; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_320 = 3'h6 == i[2:0] & 3'h4 == j[2:0] ? io_mat_6_4 : _GEN_319; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_321 = 3'h6 == i[2:0] & 3'h5 == j[2:0] ? io_mat_6_5 : _GEN_320; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_322 = 3'h6 == i[2:0] & 3'h6 == j[2:0] ? io_mat_6_6 : _GEN_321; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_323 = 3'h6 == i[2:0] & 3'h7 == j[2:0] ? io_mat_6_7 : _GEN_322; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_324 = 3'h7 == i[2:0] & 3'h0 == j[2:0] ? io_mat_7_0 : _GEN_323; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_325 = 3'h7 == i[2:0] & 3'h1 == j[2:0] ? io_mat_7_1 : _GEN_324; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_326 = 3'h7 == i[2:0] & 3'h2 == j[2:0] ? io_mat_7_2 : _GEN_325; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_327 = 3'h7 == i[2:0] & 3'h3 == j[2:0] ? io_mat_7_3 : _GEN_326; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_328 = 3'h7 == i[2:0] & 3'h4 == j[2:0] ? io_mat_7_4 : _GEN_327; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_329 = 3'h7 == i[2:0] & 3'h5 == j[2:0] ? io_mat_7_5 : _GEN_328; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_330 = 3'h7 == i[2:0] & 3'h6 == j[2:0] ? io_mat_7_6 : _GEN_329; // @[MergeDIstribution.scala 68:{13,13}]
  wire [31:0] _GEN_331 = 3'h7 == i[2:0] & 3'h7 == j[2:0] ? io_mat_7_7 : _GEN_330; // @[MergeDIstribution.scala 68:{13,13}]
  wire  _T_26 = j == 32'h7; // @[MergeDIstribution.scala 104:49]
  wire [31:0] _i_T_3 = i + 32'h1; // @[MergeDIstribution.scala 105:16]
  wire [31:0] _j_T_1 = j + 32'h1; // @[MergeDIstribution.scala 108:16]
  wire [31:0] _GEN_460 = i == 32'h7 & _T_26 ? j : _GEN_200; // @[MergeDIstribution.scala 109:75 110:11]
  wire [31:0] _GEN_461 = i <= 32'h7 & j < 32'h7 ? _j_T_1 : _GEN_460; // @[MergeDIstribution.scala 107:74 108:11]
  wire  _GEN_466 = _GEN_331 == 32'h4 | i == 32'h3 & j == 32'h3; // @[MergeDIstribution.scala 100:44 103:18 24:14]
  wire  counter = check >= 32'h1; // @[MergeDIstribution.scala 60:17]
  assign io_valid = _GEN_202 ? _GEN_466 : i == 32'h3 & j == 32'h3; // @[MergeDIstribution.scala 24:14 97:14]
  assign io_Omat_0_0 = b_0_0; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_0_1 = b_0_1; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_0_2 = b_0_2; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_0_3 = b_0_3; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_0_4 = b_0_4; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_0_5 = b_0_5; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_0_6 = b_0_6; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_0_7 = b_0_7; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_1_0 = b_1_0; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_1_1 = b_1_1; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_1_2 = b_1_2; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_1_3 = b_1_3; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_1_4 = b_1_4; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_1_5 = b_1_5; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_1_6 = b_1_6; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_1_7 = b_1_7; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_2_0 = b_2_0; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_2_1 = b_2_1; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_2_2 = b_2_2; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_2_3 = b_2_3; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_2_4 = b_2_4; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_2_5 = b_2_5; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_2_6 = b_2_6; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_2_7 = b_2_7; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_3_0 = b_3_0; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_3_1 = b_3_1; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_3_2 = b_3_2; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_3_3 = b_3_3; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_3_4 = b_3_4; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_3_5 = b_3_5; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_3_6 = b_3_6; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_3_7 = b_3_7; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_4_0 = b_4_0; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_4_1 = b_4_1; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_4_2 = b_4_2; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_4_3 = b_4_3; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_4_4 = b_4_4; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_4_5 = b_4_5; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_4_6 = b_4_6; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_4_7 = b_4_7; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_5_0 = b_5_0; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_5_1 = b_5_1; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_5_2 = b_5_2; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_5_3 = b_5_3; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_5_4 = b_5_4; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_5_5 = b_5_5; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_5_6 = b_5_6; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_5_7 = b_5_7; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_6_0 = b_6_0; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_6_1 = b_6_1; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_6_2 = b_6_2; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_6_3 = b_6_3; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_6_4 = b_6_4; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_6_5 = b_6_5; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_6_6 = b_6_6; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_6_7 = b_6_7; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_7_0 = b_7_0; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_7_1 = b_7_1; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_7_2 = b_7_2; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_7_3 = b_7_3; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_7_4 = b_7_4; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_7_5 = b_7_5; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_7_6 = b_7_6; // @[MergeDIstribution.scala 19:13]
  assign io_Omat_7_7 = b_7_7; // @[MergeDIstribution.scala 19:13]
  always @(posedge clock) begin
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_0_0 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h0 == i[2:0] & 3'h0 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_0_0 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_0_0 <= _GEN_330;
        end
      end else begin
        b_0_0 <= _GEN_135;
      end
    end else begin
      b_0_0 <= _GEN_135;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_0_1 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h0 == i[2:0] & 3'h1 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_0_1 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_0_1 <= _GEN_330;
        end
      end else begin
        b_0_1 <= _GEN_136;
      end
    end else begin
      b_0_1 <= _GEN_136;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_0_2 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h0 == i[2:0] & 3'h2 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_0_2 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_0_2 <= _GEN_330;
        end
      end else begin
        b_0_2 <= _GEN_137;
      end
    end else begin
      b_0_2 <= _GEN_137;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_0_3 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h0 == i[2:0] & 3'h3 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_0_3 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_0_3 <= _GEN_330;
        end
      end else begin
        b_0_3 <= _GEN_138;
      end
    end else begin
      b_0_3 <= _GEN_138;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_0_4 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h0 == i[2:0] & 3'h4 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_0_4 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_0_4 <= _GEN_330;
        end
      end else begin
        b_0_4 <= _GEN_139;
      end
    end else begin
      b_0_4 <= _GEN_139;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_0_5 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h0 == i[2:0] & 3'h5 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_0_5 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_0_5 <= _GEN_330;
        end
      end else begin
        b_0_5 <= _GEN_140;
      end
    end else begin
      b_0_5 <= _GEN_140;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_0_6 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h0 == i[2:0] & 3'h6 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_0_6 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_0_6 <= _GEN_330;
        end
      end else begin
        b_0_6 <= _GEN_141;
      end
    end else begin
      b_0_6 <= _GEN_141;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_0_7 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h0 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_0_7 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_0_7 <= _GEN_330;
        end
      end else begin
        b_0_7 <= _GEN_142;
      end
    end else begin
      b_0_7 <= _GEN_142;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_1_0 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h1 == i[2:0] & 3'h0 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_1_0 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_1_0 <= _GEN_330;
        end
      end else begin
        b_1_0 <= _GEN_143;
      end
    end else begin
      b_1_0 <= _GEN_143;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_1_1 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h1 == i[2:0] & 3'h1 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_1_1 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_1_1 <= _GEN_330;
        end
      end else begin
        b_1_1 <= _GEN_144;
      end
    end else begin
      b_1_1 <= _GEN_144;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_1_2 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h1 == i[2:0] & 3'h2 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_1_2 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_1_2 <= _GEN_330;
        end
      end else begin
        b_1_2 <= _GEN_145;
      end
    end else begin
      b_1_2 <= _GEN_145;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_1_3 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h1 == i[2:0] & 3'h3 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_1_3 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_1_3 <= _GEN_330;
        end
      end else begin
        b_1_3 <= _GEN_146;
      end
    end else begin
      b_1_3 <= _GEN_146;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_1_4 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h1 == i[2:0] & 3'h4 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_1_4 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_1_4 <= _GEN_330;
        end
      end else begin
        b_1_4 <= _GEN_147;
      end
    end else begin
      b_1_4 <= _GEN_147;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_1_5 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h1 == i[2:0] & 3'h5 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_1_5 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_1_5 <= _GEN_330;
        end
      end else begin
        b_1_5 <= _GEN_148;
      end
    end else begin
      b_1_5 <= _GEN_148;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_1_6 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h1 == i[2:0] & 3'h6 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_1_6 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_1_6 <= _GEN_330;
        end
      end else begin
        b_1_6 <= _GEN_149;
      end
    end else begin
      b_1_6 <= _GEN_149;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_1_7 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h1 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_1_7 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_1_7 <= _GEN_330;
        end
      end else begin
        b_1_7 <= _GEN_150;
      end
    end else begin
      b_1_7 <= _GEN_150;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_2_0 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h2 == i[2:0] & 3'h0 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_2_0 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_2_0 <= _GEN_330;
        end
      end else begin
        b_2_0 <= _GEN_151;
      end
    end else begin
      b_2_0 <= _GEN_151;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_2_1 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h2 == i[2:0] & 3'h1 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_2_1 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_2_1 <= _GEN_330;
        end
      end else begin
        b_2_1 <= _GEN_152;
      end
    end else begin
      b_2_1 <= _GEN_152;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_2_2 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h2 == i[2:0] & 3'h2 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_2_2 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_2_2 <= _GEN_330;
        end
      end else begin
        b_2_2 <= _GEN_153;
      end
    end else begin
      b_2_2 <= _GEN_153;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_2_3 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h2 == i[2:0] & 3'h3 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_2_3 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_2_3 <= _GEN_330;
        end
      end else begin
        b_2_3 <= _GEN_154;
      end
    end else begin
      b_2_3 <= _GEN_154;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_2_4 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h2 == i[2:0] & 3'h4 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_2_4 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_2_4 <= _GEN_330;
        end
      end else begin
        b_2_4 <= _GEN_155;
      end
    end else begin
      b_2_4 <= _GEN_155;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_2_5 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h2 == i[2:0] & 3'h5 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_2_5 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_2_5 <= _GEN_330;
        end
      end else begin
        b_2_5 <= _GEN_156;
      end
    end else begin
      b_2_5 <= _GEN_156;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_2_6 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h2 == i[2:0] & 3'h6 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_2_6 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_2_6 <= _GEN_330;
        end
      end else begin
        b_2_6 <= _GEN_157;
      end
    end else begin
      b_2_6 <= _GEN_157;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_2_7 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h2 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_2_7 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_2_7 <= _GEN_330;
        end
      end else begin
        b_2_7 <= _GEN_158;
      end
    end else begin
      b_2_7 <= _GEN_158;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_3_0 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h3 == i[2:0] & 3'h0 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_3_0 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_3_0 <= _GEN_330;
        end
      end else begin
        b_3_0 <= _GEN_159;
      end
    end else begin
      b_3_0 <= _GEN_159;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_3_1 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h3 == i[2:0] & 3'h1 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_3_1 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_3_1 <= _GEN_330;
        end
      end else begin
        b_3_1 <= _GEN_160;
      end
    end else begin
      b_3_1 <= _GEN_160;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_3_2 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h3 == i[2:0] & 3'h2 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_3_2 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_3_2 <= _GEN_330;
        end
      end else begin
        b_3_2 <= _GEN_161;
      end
    end else begin
      b_3_2 <= _GEN_161;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_3_3 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h3 == i[2:0] & 3'h3 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_3_3 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_3_3 <= _GEN_330;
        end
      end else begin
        b_3_3 <= _GEN_162;
      end
    end else begin
      b_3_3 <= _GEN_162;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_3_4 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h3 == i[2:0] & 3'h4 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_3_4 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_3_4 <= _GEN_330;
        end
      end else begin
        b_3_4 <= _GEN_163;
      end
    end else begin
      b_3_4 <= _GEN_163;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_3_5 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h3 == i[2:0] & 3'h5 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_3_5 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_3_5 <= _GEN_330;
        end
      end else begin
        b_3_5 <= _GEN_164;
      end
    end else begin
      b_3_5 <= _GEN_164;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_3_6 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h3 == i[2:0] & 3'h6 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_3_6 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_3_6 <= _GEN_330;
        end
      end else begin
        b_3_6 <= _GEN_165;
      end
    end else begin
      b_3_6 <= _GEN_165;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_3_7 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h3 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_3_7 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_3_7 <= _GEN_330;
        end
      end else begin
        b_3_7 <= _GEN_166;
      end
    end else begin
      b_3_7 <= _GEN_166;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_4_0 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h4 == i[2:0] & 3'h0 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_4_0 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_4_0 <= _GEN_330;
        end
      end else begin
        b_4_0 <= _GEN_167;
      end
    end else begin
      b_4_0 <= _GEN_167;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_4_1 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h4 == i[2:0] & 3'h1 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_4_1 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_4_1 <= _GEN_330;
        end
      end else begin
        b_4_1 <= _GEN_168;
      end
    end else begin
      b_4_1 <= _GEN_168;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_4_2 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h4 == i[2:0] & 3'h2 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_4_2 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_4_2 <= _GEN_330;
        end
      end else begin
        b_4_2 <= _GEN_169;
      end
    end else begin
      b_4_2 <= _GEN_169;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_4_3 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h4 == i[2:0] & 3'h3 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_4_3 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_4_3 <= _GEN_330;
        end
      end else begin
        b_4_3 <= _GEN_170;
      end
    end else begin
      b_4_3 <= _GEN_170;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_4_4 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h4 == i[2:0] & 3'h4 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_4_4 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_4_4 <= _GEN_330;
        end
      end else begin
        b_4_4 <= _GEN_171;
      end
    end else begin
      b_4_4 <= _GEN_171;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_4_5 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h4 == i[2:0] & 3'h5 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_4_5 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_4_5 <= _GEN_330;
        end
      end else begin
        b_4_5 <= _GEN_172;
      end
    end else begin
      b_4_5 <= _GEN_172;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_4_6 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h4 == i[2:0] & 3'h6 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_4_6 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_4_6 <= _GEN_330;
        end
      end else begin
        b_4_6 <= _GEN_173;
      end
    end else begin
      b_4_6 <= _GEN_173;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_4_7 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h4 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_4_7 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_4_7 <= _GEN_330;
        end
      end else begin
        b_4_7 <= _GEN_174;
      end
    end else begin
      b_4_7 <= _GEN_174;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_5_0 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h5 == i[2:0] & 3'h0 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_5_0 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_5_0 <= _GEN_330;
        end
      end else begin
        b_5_0 <= _GEN_175;
      end
    end else begin
      b_5_0 <= _GEN_175;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_5_1 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h5 == i[2:0] & 3'h1 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_5_1 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_5_1 <= _GEN_330;
        end
      end else begin
        b_5_1 <= _GEN_176;
      end
    end else begin
      b_5_1 <= _GEN_176;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_5_2 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h5 == i[2:0] & 3'h2 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_5_2 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_5_2 <= _GEN_330;
        end
      end else begin
        b_5_2 <= _GEN_177;
      end
    end else begin
      b_5_2 <= _GEN_177;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_5_3 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h5 == i[2:0] & 3'h3 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_5_3 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_5_3 <= _GEN_330;
        end
      end else begin
        b_5_3 <= _GEN_178;
      end
    end else begin
      b_5_3 <= _GEN_178;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_5_4 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h5 == i[2:0] & 3'h4 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_5_4 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_5_4 <= _GEN_330;
        end
      end else begin
        b_5_4 <= _GEN_179;
      end
    end else begin
      b_5_4 <= _GEN_179;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_5_5 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h5 == i[2:0] & 3'h5 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_5_5 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_5_5 <= _GEN_330;
        end
      end else begin
        b_5_5 <= _GEN_180;
      end
    end else begin
      b_5_5 <= _GEN_180;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_5_6 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h5 == i[2:0] & 3'h6 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_5_6 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_5_6 <= _GEN_330;
        end
      end else begin
        b_5_6 <= _GEN_181;
      end
    end else begin
      b_5_6 <= _GEN_181;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_5_7 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h5 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_5_7 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_5_7 <= _GEN_330;
        end
      end else begin
        b_5_7 <= _GEN_182;
      end
    end else begin
      b_5_7 <= _GEN_182;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_6_0 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h6 == i[2:0] & 3'h0 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_6_0 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_6_0 <= _GEN_330;
        end
      end else begin
        b_6_0 <= _GEN_183;
      end
    end else begin
      b_6_0 <= _GEN_183;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_6_1 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h6 == i[2:0] & 3'h1 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_6_1 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_6_1 <= _GEN_330;
        end
      end else begin
        b_6_1 <= _GEN_184;
      end
    end else begin
      b_6_1 <= _GEN_184;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_6_2 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h6 == i[2:0] & 3'h2 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_6_2 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_6_2 <= _GEN_330;
        end
      end else begin
        b_6_2 <= _GEN_185;
      end
    end else begin
      b_6_2 <= _GEN_185;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_6_3 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h6 == i[2:0] & 3'h3 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_6_3 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_6_3 <= _GEN_330;
        end
      end else begin
        b_6_3 <= _GEN_186;
      end
    end else begin
      b_6_3 <= _GEN_186;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_6_4 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h6 == i[2:0] & 3'h4 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_6_4 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_6_4 <= _GEN_330;
        end
      end else begin
        b_6_4 <= _GEN_187;
      end
    end else begin
      b_6_4 <= _GEN_187;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_6_5 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h6 == i[2:0] & 3'h5 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_6_5 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_6_5 <= _GEN_330;
        end
      end else begin
        b_6_5 <= _GEN_188;
      end
    end else begin
      b_6_5 <= _GEN_188;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_6_6 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h6 == i[2:0] & 3'h6 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_6_6 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_6_6 <= _GEN_330;
        end
      end else begin
        b_6_6 <= _GEN_189;
      end
    end else begin
      b_6_6 <= _GEN_189;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_6_7 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h6 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_6_7 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_6_7 <= _GEN_330;
        end
      end else begin
        b_6_7 <= _GEN_190;
      end
    end else begin
      b_6_7 <= _GEN_190;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_7_0 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h7 == i[2:0] & 3'h0 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_7_0 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_7_0 <= _GEN_330;
        end
      end else begin
        b_7_0 <= _GEN_191;
      end
    end else begin
      b_7_0 <= _GEN_191;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_7_1 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h7 == i[2:0] & 3'h1 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_7_1 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_7_1 <= _GEN_330;
        end
      end else begin
        b_7_1 <= _GEN_192;
      end
    end else begin
      b_7_1 <= _GEN_192;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_7_2 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h7 == i[2:0] & 3'h2 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_7_2 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_7_2 <= _GEN_330;
        end
      end else begin
        b_7_2 <= _GEN_193;
      end
    end else begin
      b_7_2 <= _GEN_193;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_7_3 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h7 == i[2:0] & 3'h3 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_7_3 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_7_3 <= _GEN_330;
        end
      end else begin
        b_7_3 <= _GEN_194;
      end
    end else begin
      b_7_3 <= _GEN_194;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_7_4 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h7 == i[2:0] & 3'h4 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_7_4 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_7_4 <= _GEN_330;
        end
      end else begin
        b_7_4 <= _GEN_195;
      end
    end else begin
      b_7_4 <= _GEN_195;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_7_5 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h7 == i[2:0] & 3'h5 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_7_5 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_7_5 <= _GEN_330;
        end
      end else begin
        b_7_5 <= _GEN_196;
      end
    end else begin
      b_7_5 <= _GEN_196;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_7_6 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h7 == i[2:0] & 3'h6 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_7_6 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_7_6 <= _GEN_330;
        end
      end else begin
        b_7_6 <= _GEN_197;
      end
    end else begin
      b_7_6 <= _GEN_197;
    end
    if (reset) begin // @[MergeDIstribution.scala 18:20]
      b_7_7 <= 32'h0; // @[MergeDIstribution.scala 18:20]
    end else if (io_merge) begin // @[MergeDIstribution.scala 67:19]
      if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDIstribution.scala 68:13]
          b_7_7 <= io_mat_7_7; // @[MergeDIstribution.scala 68:13]
        end else begin
          b_7_7 <= _GEN_330;
        end
      end else begin
        b_7_7 <= _GEN_198;
      end
    end else begin
      b_7_7 <= _GEN_198;
    end
    if (reset) begin // @[MergeDIstribution.scala 20:24]
      check <= 32'h0; // @[MergeDIstribution.scala 20:24]
    end else if (check >= 32'h1) begin // @[MergeDIstribution.scala 60:24]
      check <= _check_T_1; // @[MergeDIstribution.scala 62:15]
    end else if (io_i_valid & i == 32'h0 & j == 32'h0) begin // @[MergeDIstribution.scala 54:53]
      check <= _check_T_1; // @[MergeDIstribution.scala 57:15]
    end
    if (reset) begin // @[MergeDIstribution.scala 22:20]
      i <= 32'h0; // @[MergeDIstribution.scala 22:20]
    end else if (_GEN_202) begin // @[MergeDIstribution.scala 97:14]
      if (!(_GEN_331 == 32'h4)) begin // @[MergeDIstribution.scala 100:44]
        if (i < 32'h7 & j == 32'h7) begin // @[MergeDIstribution.scala 104:75]
          i <= _i_T_3; // @[MergeDIstribution.scala 105:11]
        end else begin
          i <= _GEN_199;
        end
      end
    end else begin
      i <= _GEN_199;
    end
    if (reset) begin // @[MergeDIstribution.scala 23:20]
      j <= 32'h0; // @[MergeDIstribution.scala 23:20]
    end else if (_GEN_202) begin // @[MergeDIstribution.scala 97:14]
      if (!(_GEN_331 == 32'h4)) begin // @[MergeDIstribution.scala 100:44]
        if (i < 32'h7 & j == 32'h7) begin // @[MergeDIstribution.scala 104:75]
          j <= 32'h0; // @[MergeDIstribution.scala 106:11]
        end else begin
          j <= _GEN_461;
        end
      end
    end else if (io_i_valid & i == 32'h0 & j == 32'h0) begin // @[MergeDIstribution.scala 54:53]
      j <= 32'h0; // @[MergeDIstribution.scala 56:11]
    end
    if (reset) begin // @[MergeDIstribution.scala 26:20]
      k <= 32'h0; // @[MergeDIstribution.scala 26:20]
    end else if (io_merge & delay == 32'h8) begin // @[MergeDIstribution.scala 41:53]
      if (k < io_IDex & l == 32'h7) begin // @[MergeDIstribution.scala 43:56]
        k <= _k_T_1; // @[MergeDIstribution.scala 44:11]
      end
    end
    if (reset) begin // @[MergeDIstribution.scala 27:20]
      l <= 32'h0; // @[MergeDIstribution.scala 27:20]
    end else if (io_merge & delay == 32'h8) begin // @[MergeDIstribution.scala 41:53]
      if (k < io_IDex & l == 32'h7) begin // @[MergeDIstribution.scala 43:56]
        l <= 32'h0; // @[MergeDIstribution.scala 45:11]
      end else if (k <= io_IDex & l < 32'h7) begin // @[MergeDIstribution.scala 46:61]
        l <= _l_T_1; // @[MergeDIstribution.scala 47:11]
      end
    end
    if (reset) begin // @[MergeDIstribution.scala 29:24]
      delay <= 32'h0; // @[MergeDIstribution.scala 29:24]
    end else if (delay <= 32'h7 & io_merge) begin // @[MergeDIstribution.scala 31:53]
      delay <= _delay_T_1; // @[MergeDIstribution.scala 32:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  b_0_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  b_0_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  b_0_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  b_0_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  b_0_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  b_0_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  b_0_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  b_0_7 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  b_1_0 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  b_1_1 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  b_1_2 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  b_1_3 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  b_1_4 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  b_1_5 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  b_1_6 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  b_1_7 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  b_2_0 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  b_2_1 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  b_2_2 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  b_2_3 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  b_2_4 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  b_2_5 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  b_2_6 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  b_2_7 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  b_3_0 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  b_3_1 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  b_3_2 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  b_3_3 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  b_3_4 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  b_3_5 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  b_3_6 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  b_3_7 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  b_4_0 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  b_4_1 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  b_4_2 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  b_4_3 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  b_4_4 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  b_4_5 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  b_4_6 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  b_4_7 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  b_5_0 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  b_5_1 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  b_5_2 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  b_5_3 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  b_5_4 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  b_5_5 = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  b_5_6 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  b_5_7 = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  b_6_0 = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  b_6_1 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  b_6_2 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  b_6_3 = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  b_6_4 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  b_6_5 = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  b_6_6 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  b_6_7 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  b_7_0 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  b_7_1 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  b_7_2 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  b_7_3 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  b_7_4 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  b_7_5 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  b_7_6 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  b_7_7 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  check = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  i = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  j = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  k = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  l = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  delay = _RAND_69[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Distribution(
  input         clock,
  input         reset,
  input  [31:0] io_matrix_0_0,
  input  [31:0] io_matrix_0_1,
  input  [31:0] io_matrix_0_2,
  input  [31:0] io_matrix_0_3,
  input  [31:0] io_matrix_0_4,
  input  [31:0] io_matrix_0_5,
  input  [31:0] io_matrix_0_6,
  input  [31:0] io_matrix_0_7,
  input  [31:0] io_matrix_1_0,
  input  [31:0] io_matrix_1_1,
  input  [31:0] io_matrix_1_2,
  input  [31:0] io_matrix_1_3,
  input  [31:0] io_matrix_1_4,
  input  [31:0] io_matrix_1_5,
  input  [31:0] io_matrix_1_6,
  input  [31:0] io_matrix_1_7,
  input  [31:0] io_matrix_2_0,
  input  [31:0] io_matrix_2_1,
  input  [31:0] io_matrix_2_2,
  input  [31:0] io_matrix_2_3,
  input  [31:0] io_matrix_2_4,
  input  [31:0] io_matrix_2_5,
  input  [31:0] io_matrix_2_6,
  input  [31:0] io_matrix_2_7,
  input  [31:0] io_matrix_3_0,
  input  [31:0] io_matrix_3_1,
  input  [31:0] io_matrix_3_2,
  input  [31:0] io_matrix_3_3,
  input  [31:0] io_matrix_3_4,
  input  [31:0] io_matrix_3_5,
  input  [31:0] io_matrix_3_6,
  input  [31:0] io_matrix_3_7,
  input  [31:0] io_matrix_4_0,
  input  [31:0] io_matrix_4_1,
  input  [31:0] io_matrix_4_2,
  input  [31:0] io_matrix_4_3,
  input  [31:0] io_matrix_4_4,
  input  [31:0] io_matrix_4_5,
  input  [31:0] io_matrix_4_6,
  input  [31:0] io_matrix_4_7,
  input  [31:0] io_matrix_5_0,
  input  [31:0] io_matrix_5_1,
  input  [31:0] io_matrix_5_2,
  input  [31:0] io_matrix_5_3,
  input  [31:0] io_matrix_5_4,
  input  [31:0] io_matrix_5_5,
  input  [31:0] io_matrix_5_6,
  input  [31:0] io_matrix_5_7,
  input  [31:0] io_matrix_6_0,
  input  [31:0] io_matrix_6_1,
  input  [31:0] io_matrix_6_2,
  input  [31:0] io_matrix_6_3,
  input  [31:0] io_matrix_6_4,
  input  [31:0] io_matrix_6_5,
  input  [31:0] io_matrix_6_6,
  input  [31:0] io_matrix_6_7,
  input  [31:0] io_matrix_7_0,
  input  [31:0] io_matrix_7_1,
  input  [31:0] io_matrix_7_2,
  input  [31:0] io_matrix_7_3,
  input  [31:0] io_matrix_7_4,
  input  [31:0] io_matrix_7_5,
  input  [31:0] io_matrix_7_6,
  input  [31:0] io_matrix_7_7,
  input  [31:0] io_s,
  output [31:0] io_out_0_0,
  output [31:0] io_out_0_1,
  output [31:0] io_out_0_2,
  output [31:0] io_out_0_3,
  output [31:0] io_out_0_4,
  output [31:0] io_out_0_5,
  output [31:0] io_out_0_6,
  output [31:0] io_out_0_7,
  output [31:0] io_out_1_0,
  output [31:0] io_out_1_1,
  output [31:0] io_out_1_2,
  output [31:0] io_out_1_3,
  output [31:0] io_out_1_4,
  output [31:0] io_out_1_5,
  output [31:0] io_out_1_6,
  output [31:0] io_out_1_7,
  output [31:0] io_out_2_0,
  output [31:0] io_out_2_1,
  output [31:0] io_out_2_2,
  output [31:0] io_out_2_3,
  output [31:0] io_out_2_4,
  output [31:0] io_out_2_5,
  output [31:0] io_out_2_6,
  output [31:0] io_out_2_7,
  output [31:0] io_out_3_0,
  output [31:0] io_out_3_1,
  output [31:0] io_out_3_2,
  output [31:0] io_out_3_3,
  output [31:0] io_out_3_4,
  output [31:0] io_out_3_5,
  output [31:0] io_out_3_6,
  output [31:0] io_out_3_7,
  output [31:0] io_out_4_0,
  output [31:0] io_out_4_1,
  output [31:0] io_out_4_2,
  output [31:0] io_out_4_3,
  output [31:0] io_out_4_4,
  output [31:0] io_out_4_5,
  output [31:0] io_out_4_6,
  output [31:0] io_out_4_7,
  output [31:0] io_out_5_0,
  output [31:0] io_out_5_1,
  output [31:0] io_out_5_2,
  output [31:0] io_out_5_3,
  output [31:0] io_out_5_4,
  output [31:0] io_out_5_5,
  output [31:0] io_out_5_6,
  output [31:0] io_out_5_7,
  output [31:0] io_out_6_0,
  output [31:0] io_out_6_1,
  output [31:0] io_out_6_2,
  output [31:0] io_out_6_3,
  output [31:0] io_out_6_4,
  output [31:0] io_out_6_5,
  output [31:0] io_out_6_6,
  output [31:0] io_out_6_7,
  output [31:0] io_out_7_0,
  output [31:0] io_out_7_1,
  output [31:0] io_out_7_2,
  output [31:0] io_out_7_3,
  output [31:0] io_out_7_4,
  output [31:0] io_out_7_5,
  output [31:0] io_out_7_6,
  output [31:0] io_out_7_7,
  output        io_ProcessValid,
  input         io_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
`endif // RANDOMIZE_REG_INIT
  wire  part2_clock; // @[DIstribution.scala 55:19]
  wire  part2_reset; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_IDex; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_JDex; // @[DIstribution.scala 55:19]
  wire  part2_io_valid; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_0_0; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_0_1; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_0_2; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_0_3; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_0_4; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_0_5; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_0_6; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_0_7; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_1_0; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_1_1; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_1_2; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_1_3; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_1_4; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_1_5; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_1_6; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_1_7; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_2_0; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_2_1; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_2_2; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_2_3; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_2_4; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_2_5; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_2_6; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_2_7; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_3_0; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_3_1; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_3_2; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_3_3; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_3_4; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_3_5; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_3_6; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_3_7; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_4_0; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_4_1; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_4_2; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_4_3; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_4_4; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_4_5; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_4_6; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_4_7; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_5_0; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_5_1; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_5_2; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_5_3; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_5_4; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_5_5; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_5_6; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_5_7; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_6_0; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_6_1; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_6_2; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_6_3; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_6_4; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_6_5; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_6_6; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_6_7; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_7_0; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_7_1; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_7_2; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_7_3; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_7_4; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_7_5; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_7_6; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_mat_7_7; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_0_0; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_0_1; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_0_2; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_0_3; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_0_4; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_0_5; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_0_6; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_0_7; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_1_0; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_1_1; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_1_2; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_1_3; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_1_4; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_1_5; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_1_6; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_1_7; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_2_0; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_2_1; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_2_2; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_2_3; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_2_4; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_2_5; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_2_6; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_2_7; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_3_0; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_3_1; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_3_2; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_3_3; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_3_4; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_3_5; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_3_6; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_3_7; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_4_0; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_4_1; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_4_2; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_4_3; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_4_4; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_4_5; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_4_6; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_4_7; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_5_0; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_5_1; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_5_2; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_5_3; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_5_4; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_5_5; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_5_6; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_5_7; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_6_0; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_6_1; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_6_2; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_6_3; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_6_4; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_6_5; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_6_6; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_6_7; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_7_0; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_7_1; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_7_2; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_7_3; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_7_4; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_7_5; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_7_6; // @[DIstribution.scala 55:19]
  wire [31:0] part2_io_OutMat_7_7; // @[DIstribution.scala 55:19]
  wire  part2_io_Ovalid; // @[DIstribution.scala 55:19]
  wire  part2_io_ProcessValid; // @[DIstribution.scala 55:19]
  wire  part3_clock; // @[DIstribution.scala 69:23]
  wire  part3_reset; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_0_0; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_0_1; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_0_2; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_0_3; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_0_4; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_0_5; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_0_6; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_0_7; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_1_0; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_1_1; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_1_2; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_1_3; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_1_4; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_1_5; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_1_6; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_1_7; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_2_0; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_2_1; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_2_2; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_2_3; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_2_4; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_2_5; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_2_6; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_2_7; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_3_0; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_3_1; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_3_2; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_3_3; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_3_4; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_3_5; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_3_6; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_3_7; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_4_0; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_4_1; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_4_2; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_4_3; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_4_4; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_4_5; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_4_6; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_4_7; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_5_0; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_5_1; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_5_2; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_5_3; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_5_4; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_5_5; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_5_6; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_5_7; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_6_0; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_6_1; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_6_2; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_6_3; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_6_4; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_6_5; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_6_6; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_6_7; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_7_0; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_7_1; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_7_2; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_7_3; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_7_4; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_7_5; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_7_6; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_PreMat_7_7; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_IDex; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_0_0; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_0_1; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_0_2; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_0_3; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_0_4; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_0_5; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_0_6; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_0_7; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_1_0; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_1_1; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_1_2; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_1_3; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_1_4; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_1_5; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_1_6; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_1_7; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_2_0; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_2_1; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_2_2; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_2_3; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_2_4; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_2_5; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_2_6; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_2_7; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_3_0; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_3_1; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_3_2; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_3_3; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_3_4; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_3_5; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_3_6; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_3_7; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_4_0; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_4_1; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_4_2; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_4_3; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_4_4; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_4_5; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_4_6; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_4_7; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_5_0; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_5_1; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_5_2; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_5_3; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_5_4; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_5_5; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_5_6; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_5_7; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_6_0; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_6_1; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_6_2; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_6_3; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_6_4; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_6_5; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_6_6; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_6_7; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_7_0; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_7_1; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_7_2; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_7_3; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_7_4; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_7_5; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_7_6; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_mat_7_7; // @[DIstribution.scala 69:23]
  wire  part3_io_i_valid; // @[DIstribution.scala 69:23]
  wire  part3_io_valid; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_0_0; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_0_1; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_0_2; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_0_3; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_0_4; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_0_5; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_0_6; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_0_7; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_1_0; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_1_1; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_1_2; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_1_3; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_1_4; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_1_5; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_1_6; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_1_7; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_2_0; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_2_1; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_2_2; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_2_3; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_2_4; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_2_5; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_2_6; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_2_7; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_3_0; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_3_1; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_3_2; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_3_3; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_3_4; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_3_5; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_3_6; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_3_7; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_4_0; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_4_1; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_4_2; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_4_3; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_4_4; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_4_5; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_4_6; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_4_7; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_5_0; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_5_1; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_5_2; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_5_3; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_5_4; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_5_5; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_5_6; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_5_7; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_6_0; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_6_1; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_6_2; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_6_3; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_6_4; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_6_5; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_6_6; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_6_7; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_7_0; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_7_1; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_7_2; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_7_3; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_7_4; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_7_5; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_7_6; // @[DIstribution.scala 69:23]
  wire [31:0] part3_io_Omat_7_7; // @[DIstribution.scala 69:23]
  wire  part3_io_merge; // @[DIstribution.scala 69:23]
  reg [31:0] i; // @[DIstribution.scala 19:20]
  reg [31:0] j; // @[DIstribution.scala 20:20]
  reg [31:0] count; // @[DIstribution.scala 21:24]
  reg [31:0] Idex_0; // @[DIstribution.scala 22:23]
  reg [31:0] Idex_1; // @[DIstribution.scala 22:23]
  reg [31:0] Idex_2; // @[DIstribution.scala 22:23]
  reg [31:0] Idex_3; // @[DIstribution.scala 22:23]
  reg [31:0] Idex_4; // @[DIstribution.scala 22:23]
  reg [31:0] Idex_5; // @[DIstribution.scala 22:23]
  reg [31:0] Idex_6; // @[DIstribution.scala 22:23]
  reg [31:0] Idex_7; // @[DIstribution.scala 22:23]
  reg [31:0] Jdex_0; // @[DIstribution.scala 23:23]
  reg [31:0] Jdex_1; // @[DIstribution.scala 23:23]
  reg [31:0] Jdex_2; // @[DIstribution.scala 23:23]
  reg [31:0] Jdex_3; // @[DIstribution.scala 23:23]
  reg [31:0] Jdex_4; // @[DIstribution.scala 23:23]
  reg [31:0] Jdex_5; // @[DIstribution.scala 23:23]
  reg [31:0] Jdex_6; // @[DIstribution.scala 23:23]
  reg [31:0] Jdex_7; // @[DIstribution.scala 23:23]
  reg [31:0] iterationNo; // @[DIstribution.scala 25:30]
  wire  _io_validIteration_T = i == 32'h7; // @[DIstribution.scala 30:29]
  wire  _io_validIteration_T_1 = j == 32'h7; // @[DIstribution.scala 30:62]
  wire  _io_validIteration_T_2 = i == 32'h7 & j == 32'h7; // @[DIstribution.scala 30:56]
  wire [31:0] _GEN_1 = 3'h0 == i[2:0] & 3'h1 == j[2:0] ? io_matrix_0_1 : io_matrix_0_0; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_2 = 3'h0 == i[2:0] & 3'h2 == j[2:0] ? io_matrix_0_2 : _GEN_1; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_3 = 3'h0 == i[2:0] & 3'h3 == j[2:0] ? io_matrix_0_3 : _GEN_2; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_4 = 3'h0 == i[2:0] & 3'h4 == j[2:0] ? io_matrix_0_4 : _GEN_3; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_5 = 3'h0 == i[2:0] & 3'h5 == j[2:0] ? io_matrix_0_5 : _GEN_4; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_6 = 3'h0 == i[2:0] & 3'h6 == j[2:0] ? io_matrix_0_6 : _GEN_5; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_7 = 3'h0 == i[2:0] & 3'h7 == j[2:0] ? io_matrix_0_7 : _GEN_6; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_8 = 3'h1 == i[2:0] & 3'h0 == j[2:0] ? io_matrix_1_0 : _GEN_7; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_9 = 3'h1 == i[2:0] & 3'h1 == j[2:0] ? io_matrix_1_1 : _GEN_8; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_10 = 3'h1 == i[2:0] & 3'h2 == j[2:0] ? io_matrix_1_2 : _GEN_9; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_11 = 3'h1 == i[2:0] & 3'h3 == j[2:0] ? io_matrix_1_3 : _GEN_10; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_12 = 3'h1 == i[2:0] & 3'h4 == j[2:0] ? io_matrix_1_4 : _GEN_11; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_13 = 3'h1 == i[2:0] & 3'h5 == j[2:0] ? io_matrix_1_5 : _GEN_12; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_14 = 3'h1 == i[2:0] & 3'h6 == j[2:0] ? io_matrix_1_6 : _GEN_13; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_15 = 3'h1 == i[2:0] & 3'h7 == j[2:0] ? io_matrix_1_7 : _GEN_14; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_16 = 3'h2 == i[2:0] & 3'h0 == j[2:0] ? io_matrix_2_0 : _GEN_15; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_17 = 3'h2 == i[2:0] & 3'h1 == j[2:0] ? io_matrix_2_1 : _GEN_16; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_18 = 3'h2 == i[2:0] & 3'h2 == j[2:0] ? io_matrix_2_2 : _GEN_17; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_19 = 3'h2 == i[2:0] & 3'h3 == j[2:0] ? io_matrix_2_3 : _GEN_18; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_20 = 3'h2 == i[2:0] & 3'h4 == j[2:0] ? io_matrix_2_4 : _GEN_19; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_21 = 3'h2 == i[2:0] & 3'h5 == j[2:0] ? io_matrix_2_5 : _GEN_20; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_22 = 3'h2 == i[2:0] & 3'h6 == j[2:0] ? io_matrix_2_6 : _GEN_21; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_23 = 3'h2 == i[2:0] & 3'h7 == j[2:0] ? io_matrix_2_7 : _GEN_22; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_24 = 3'h3 == i[2:0] & 3'h0 == j[2:0] ? io_matrix_3_0 : _GEN_23; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_25 = 3'h3 == i[2:0] & 3'h1 == j[2:0] ? io_matrix_3_1 : _GEN_24; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_26 = 3'h3 == i[2:0] & 3'h2 == j[2:0] ? io_matrix_3_2 : _GEN_25; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_27 = 3'h3 == i[2:0] & 3'h3 == j[2:0] ? io_matrix_3_3 : _GEN_26; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_28 = 3'h3 == i[2:0] & 3'h4 == j[2:0] ? io_matrix_3_4 : _GEN_27; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_29 = 3'h3 == i[2:0] & 3'h5 == j[2:0] ? io_matrix_3_5 : _GEN_28; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_30 = 3'h3 == i[2:0] & 3'h6 == j[2:0] ? io_matrix_3_6 : _GEN_29; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_31 = 3'h3 == i[2:0] & 3'h7 == j[2:0] ? io_matrix_3_7 : _GEN_30; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_32 = 3'h4 == i[2:0] & 3'h0 == j[2:0] ? io_matrix_4_0 : _GEN_31; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_33 = 3'h4 == i[2:0] & 3'h1 == j[2:0] ? io_matrix_4_1 : _GEN_32; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_34 = 3'h4 == i[2:0] & 3'h2 == j[2:0] ? io_matrix_4_2 : _GEN_33; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_35 = 3'h4 == i[2:0] & 3'h3 == j[2:0] ? io_matrix_4_3 : _GEN_34; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_36 = 3'h4 == i[2:0] & 3'h4 == j[2:0] ? io_matrix_4_4 : _GEN_35; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_37 = 3'h4 == i[2:0] & 3'h5 == j[2:0] ? io_matrix_4_5 : _GEN_36; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_38 = 3'h4 == i[2:0] & 3'h6 == j[2:0] ? io_matrix_4_6 : _GEN_37; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_39 = 3'h4 == i[2:0] & 3'h7 == j[2:0] ? io_matrix_4_7 : _GEN_38; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_40 = 3'h5 == i[2:0] & 3'h0 == j[2:0] ? io_matrix_5_0 : _GEN_39; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_41 = 3'h5 == i[2:0] & 3'h1 == j[2:0] ? io_matrix_5_1 : _GEN_40; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_42 = 3'h5 == i[2:0] & 3'h2 == j[2:0] ? io_matrix_5_2 : _GEN_41; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_43 = 3'h5 == i[2:0] & 3'h3 == j[2:0] ? io_matrix_5_3 : _GEN_42; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_44 = 3'h5 == i[2:0] & 3'h4 == j[2:0] ? io_matrix_5_4 : _GEN_43; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_45 = 3'h5 == i[2:0] & 3'h5 == j[2:0] ? io_matrix_5_5 : _GEN_44; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_46 = 3'h5 == i[2:0] & 3'h6 == j[2:0] ? io_matrix_5_6 : _GEN_45; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_47 = 3'h5 == i[2:0] & 3'h7 == j[2:0] ? io_matrix_5_7 : _GEN_46; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_48 = 3'h6 == i[2:0] & 3'h0 == j[2:0] ? io_matrix_6_0 : _GEN_47; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_49 = 3'h6 == i[2:0] & 3'h1 == j[2:0] ? io_matrix_6_1 : _GEN_48; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_50 = 3'h6 == i[2:0] & 3'h2 == j[2:0] ? io_matrix_6_2 : _GEN_49; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_51 = 3'h6 == i[2:0] & 3'h3 == j[2:0] ? io_matrix_6_3 : _GEN_50; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_52 = 3'h6 == i[2:0] & 3'h4 == j[2:0] ? io_matrix_6_4 : _GEN_51; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_53 = 3'h6 == i[2:0] & 3'h5 == j[2:0] ? io_matrix_6_5 : _GEN_52; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_54 = 3'h6 == i[2:0] & 3'h6 == j[2:0] ? io_matrix_6_6 : _GEN_53; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_55 = 3'h6 == i[2:0] & 3'h7 == j[2:0] ? io_matrix_6_7 : _GEN_54; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_56 = 3'h7 == i[2:0] & 3'h0 == j[2:0] ? io_matrix_7_0 : _GEN_55; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_57 = 3'h7 == i[2:0] & 3'h1 == j[2:0] ? io_matrix_7_1 : _GEN_56; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_58 = 3'h7 == i[2:0] & 3'h2 == j[2:0] ? io_matrix_7_2 : _GEN_57; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_59 = 3'h7 == i[2:0] & 3'h3 == j[2:0] ? io_matrix_7_3 : _GEN_58; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_60 = 3'h7 == i[2:0] & 3'h4 == j[2:0] ? io_matrix_7_4 : _GEN_59; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_61 = 3'h7 == i[2:0] & 3'h5 == j[2:0] ? io_matrix_7_5 : _GEN_60; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_62 = 3'h7 == i[2:0] & 3'h6 == j[2:0] ? io_matrix_7_6 : _GEN_61; // @[DIstribution.scala 34:{27,27}]
  wire [31:0] _GEN_63 = 3'h7 == i[2:0] & 3'h7 == j[2:0] ? io_matrix_7_7 : _GEN_62; // @[DIstribution.scala 34:{27,27}]
  wire  _T_2 = _GEN_63 == 32'h1; // @[DIstribution.scala 34:27]
  wire [31:0] _iterationNo_T_1 = iterationNo + 32'h1; // @[DIstribution.scala 35:34]
  wire [31:0] _count_T_1 = count + 32'h1; // @[DIstribution.scala 48:24]
  wire [31:0] _GEN_129 = 3'h0 == count[2:0] ? i : Idex_0; // @[DIstribution.scala 49:{21,21} 22:23]
  wire [31:0] _GEN_130 = 3'h1 == count[2:0] ? i : Idex_1; // @[DIstribution.scala 49:{21,21} 22:23]
  wire [31:0] _GEN_131 = 3'h2 == count[2:0] ? i : Idex_2; // @[DIstribution.scala 49:{21,21} 22:23]
  wire [31:0] _GEN_132 = 3'h3 == count[2:0] ? i : Idex_3; // @[DIstribution.scala 49:{21,21} 22:23]
  wire [31:0] _GEN_133 = 3'h4 == count[2:0] ? i : Idex_4; // @[DIstribution.scala 49:{21,21} 22:23]
  wire [31:0] _GEN_134 = 3'h5 == count[2:0] ? i : Idex_5; // @[DIstribution.scala 49:{21,21} 22:23]
  wire [31:0] _GEN_135 = 3'h6 == count[2:0] ? i : Idex_6; // @[DIstribution.scala 49:{21,21} 22:23]
  wire [31:0] _GEN_136 = 3'h7 == count[2:0] ? i : Idex_7; // @[DIstribution.scala 49:{21,21} 22:23]
  wire [31:0] _GEN_137 = 3'h0 == count[2:0] ? j : Jdex_0; // @[DIstribution.scala 50:{21,21} 23:23]
  wire [31:0] _GEN_138 = 3'h1 == count[2:0] ? j : Jdex_1; // @[DIstribution.scala 50:{21,21} 23:23]
  wire [31:0] _GEN_139 = 3'h2 == count[2:0] ? j : Jdex_2; // @[DIstribution.scala 50:{21,21} 23:23]
  wire [31:0] _GEN_140 = 3'h3 == count[2:0] ? j : Jdex_3; // @[DIstribution.scala 50:{21,21} 23:23]
  wire [31:0] _GEN_141 = 3'h4 == count[2:0] ? j : Jdex_4; // @[DIstribution.scala 50:{21,21} 23:23]
  wire [31:0] _GEN_142 = 3'h5 == count[2:0] ? j : Jdex_5; // @[DIstribution.scala 50:{21,21} 23:23]
  wire [31:0] _GEN_143 = 3'h6 == count[2:0] ? j : Jdex_6; // @[DIstribution.scala 50:{21,21} 23:23]
  wire [31:0] _GEN_144 = 3'h7 == count[2:0] ? j : Jdex_7; // @[DIstribution.scala 50:{21,21} 23:23]
  reg  c; // @[DIstribution.scala 57:20]
  wire [31:0] _GEN_259 = 3'h1 == io_s[2:0] ? Idex_1 : Idex_0; // @[DIstribution.scala 60:{19,19}]
  wire [31:0] _GEN_260 = 3'h2 == io_s[2:0] ? Idex_2 : _GEN_259; // @[DIstribution.scala 60:{19,19}]
  wire [31:0] _GEN_261 = 3'h3 == io_s[2:0] ? Idex_3 : _GEN_260; // @[DIstribution.scala 60:{19,19}]
  wire [31:0] _GEN_262 = 3'h4 == io_s[2:0] ? Idex_4 : _GEN_261; // @[DIstribution.scala 60:{19,19}]
  wire [31:0] _GEN_263 = 3'h5 == io_s[2:0] ? Idex_5 : _GEN_262; // @[DIstribution.scala 60:{19,19}]
  wire [31:0] _GEN_264 = 3'h6 == io_s[2:0] ? Idex_6 : _GEN_263; // @[DIstribution.scala 60:{19,19}]
  wire [31:0] _GEN_265 = 3'h7 == io_s[2:0] ? Idex_7 : _GEN_264; // @[DIstribution.scala 60:{19,19}]
  wire [31:0] _GEN_267 = 3'h1 == io_s[2:0] ? Jdex_1 : Jdex_0; // @[DIstribution.scala 61:{19,19}]
  wire [31:0] _GEN_268 = 3'h2 == io_s[2:0] ? Jdex_2 : _GEN_267; // @[DIstribution.scala 61:{19,19}]
  wire [31:0] _GEN_269 = 3'h3 == io_s[2:0] ? Jdex_3 : _GEN_268; // @[DIstribution.scala 61:{19,19}]
  wire [31:0] _GEN_270 = 3'h4 == io_s[2:0] ? Jdex_4 : _GEN_269; // @[DIstribution.scala 61:{19,19}]
  wire [31:0] _GEN_271 = 3'h5 == io_s[2:0] ? Jdex_5 : _GEN_270; // @[DIstribution.scala 61:{19,19}]
  wire [31:0] _GEN_272 = 3'h6 == io_s[2:0] ? Jdex_6 : _GEN_271; // @[DIstribution.scala 61:{19,19}]
  wire [31:0] _GEN_273 = 3'h7 == io_s[2:0] ? Jdex_7 : _GEN_272; // @[DIstribution.scala 61:{19,19}]
  wire  check = part2_io_Ovalid ? 1'h0 : 1'h1; // @[DIstribution.scala 75:26 76:15 78:15]
  wire [31:0] _e_T_4 = count - 32'h1; // @[DIstribution.scala 80:85]
  wire  e = _io_validIteration_T_2 & _e_T_4 < io_s; // @[DIstribution.scala 80:75]
  reg  part3_io_merge_REG; // @[DIstribution.scala 83:30]
  wire [31:0] _GEN_293 = e ? 32'h0 : part3_io_Omat_0_0; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_294 = e ? 32'h0 : part3_io_Omat_0_1; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_295 = e ? 32'h0 : part3_io_Omat_0_2; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_296 = e ? 32'h0 : part3_io_Omat_0_3; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_297 = e ? 32'h0 : part3_io_Omat_0_4; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_298 = e ? 32'h0 : part3_io_Omat_0_5; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_299 = e ? 32'h0 : part3_io_Omat_0_6; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_300 = e ? 32'h0 : part3_io_Omat_0_7; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_301 = e ? 32'h0 : part3_io_Omat_1_0; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_302 = e ? 32'h0 : part3_io_Omat_1_1; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_303 = e ? 32'h0 : part3_io_Omat_1_2; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_304 = e ? 32'h0 : part3_io_Omat_1_3; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_305 = e ? 32'h0 : part3_io_Omat_1_4; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_306 = e ? 32'h0 : part3_io_Omat_1_5; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_307 = e ? 32'h0 : part3_io_Omat_1_6; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_308 = e ? 32'h0 : part3_io_Omat_1_7; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_309 = e ? 32'h0 : part3_io_Omat_2_0; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_310 = e ? 32'h0 : part3_io_Omat_2_1; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_311 = e ? 32'h0 : part3_io_Omat_2_2; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_312 = e ? 32'h0 : part3_io_Omat_2_3; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_313 = e ? 32'h0 : part3_io_Omat_2_4; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_314 = e ? 32'h0 : part3_io_Omat_2_5; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_315 = e ? 32'h0 : part3_io_Omat_2_6; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_316 = e ? 32'h0 : part3_io_Omat_2_7; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_317 = e ? 32'h0 : part3_io_Omat_3_0; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_318 = e ? 32'h0 : part3_io_Omat_3_1; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_319 = e ? 32'h0 : part3_io_Omat_3_2; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_320 = e ? 32'h0 : part3_io_Omat_3_3; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_321 = e ? 32'h0 : part3_io_Omat_3_4; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_322 = e ? 32'h0 : part3_io_Omat_3_5; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_323 = e ? 32'h0 : part3_io_Omat_3_6; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_324 = e ? 32'h0 : part3_io_Omat_3_7; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_325 = e ? 32'h0 : part3_io_Omat_4_0; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_326 = e ? 32'h0 : part3_io_Omat_4_1; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_327 = e ? 32'h0 : part3_io_Omat_4_2; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_328 = e ? 32'h0 : part3_io_Omat_4_3; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_329 = e ? 32'h0 : part3_io_Omat_4_4; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_330 = e ? 32'h0 : part3_io_Omat_4_5; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_331 = e ? 32'h0 : part3_io_Omat_4_6; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_332 = e ? 32'h0 : part3_io_Omat_4_7; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_333 = e ? 32'h0 : part3_io_Omat_5_0; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_334 = e ? 32'h0 : part3_io_Omat_5_1; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_335 = e ? 32'h0 : part3_io_Omat_5_2; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_336 = e ? 32'h0 : part3_io_Omat_5_3; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_337 = e ? 32'h0 : part3_io_Omat_5_4; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_338 = e ? 32'h0 : part3_io_Omat_5_5; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_339 = e ? 32'h0 : part3_io_Omat_5_6; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_340 = e ? 32'h0 : part3_io_Omat_5_7; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_341 = e ? 32'h0 : part3_io_Omat_6_0; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_342 = e ? 32'h0 : part3_io_Omat_6_1; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_343 = e ? 32'h0 : part3_io_Omat_6_2; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_344 = e ? 32'h0 : part3_io_Omat_6_3; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_345 = e ? 32'h0 : part3_io_Omat_6_4; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_346 = e ? 32'h0 : part3_io_Omat_6_5; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_347 = e ? 32'h0 : part3_io_Omat_6_6; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_348 = e ? 32'h0 : part3_io_Omat_6_7; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_349 = e ? 32'h0 : part3_io_Omat_7_0; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_350 = e ? 32'h0 : part3_io_Omat_7_1; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_351 = e ? 32'h0 : part3_io_Omat_7_2; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_352 = e ? 32'h0 : part3_io_Omat_7_3; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_353 = e ? 32'h0 : part3_io_Omat_7_4; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_354 = e ? 32'h0 : part3_io_Omat_7_5; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_355 = e ? 32'h0 : part3_io_Omat_7_6; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_356 = e ? 32'h0 : part3_io_Omat_7_7; // @[DIstribution.scala 90:96 91:16 93:12]
  wire [31:0] _GEN_357 = e ? 32'h0 : part2_io_OutMat_0_0; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_358 = e ? 32'h0 : part2_io_OutMat_0_1; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_359 = e ? 32'h0 : part2_io_OutMat_0_2; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_360 = e ? 32'h0 : part2_io_OutMat_0_3; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_361 = e ? 32'h0 : part2_io_OutMat_0_4; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_362 = e ? 32'h0 : part2_io_OutMat_0_5; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_363 = e ? 32'h0 : part2_io_OutMat_0_6; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_364 = e ? 32'h0 : part2_io_OutMat_0_7; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_365 = e ? 32'h0 : part2_io_OutMat_1_0; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_366 = e ? 32'h0 : part2_io_OutMat_1_1; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_367 = e ? 32'h0 : part2_io_OutMat_1_2; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_368 = e ? 32'h0 : part2_io_OutMat_1_3; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_369 = e ? 32'h0 : part2_io_OutMat_1_4; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_370 = e ? 32'h0 : part2_io_OutMat_1_5; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_371 = e ? 32'h0 : part2_io_OutMat_1_6; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_372 = e ? 32'h0 : part2_io_OutMat_1_7; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_373 = e ? 32'h0 : part2_io_OutMat_2_0; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_374 = e ? 32'h0 : part2_io_OutMat_2_1; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_375 = e ? 32'h0 : part2_io_OutMat_2_2; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_376 = e ? 32'h0 : part2_io_OutMat_2_3; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_377 = e ? 32'h0 : part2_io_OutMat_2_4; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_378 = e ? 32'h0 : part2_io_OutMat_2_5; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_379 = e ? 32'h0 : part2_io_OutMat_2_6; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_380 = e ? 32'h0 : part2_io_OutMat_2_7; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_381 = e ? 32'h0 : part2_io_OutMat_3_0; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_382 = e ? 32'h0 : part2_io_OutMat_3_1; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_383 = e ? 32'h0 : part2_io_OutMat_3_2; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_384 = e ? 32'h0 : part2_io_OutMat_3_3; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_385 = e ? 32'h0 : part2_io_OutMat_3_4; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_386 = e ? 32'h0 : part2_io_OutMat_3_5; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_387 = e ? 32'h0 : part2_io_OutMat_3_6; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_388 = e ? 32'h0 : part2_io_OutMat_3_7; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_389 = e ? 32'h0 : part2_io_OutMat_4_0; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_390 = e ? 32'h0 : part2_io_OutMat_4_1; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_391 = e ? 32'h0 : part2_io_OutMat_4_2; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_392 = e ? 32'h0 : part2_io_OutMat_4_3; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_393 = e ? 32'h0 : part2_io_OutMat_4_4; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_394 = e ? 32'h0 : part2_io_OutMat_4_5; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_395 = e ? 32'h0 : part2_io_OutMat_4_6; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_396 = e ? 32'h0 : part2_io_OutMat_4_7; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_397 = e ? 32'h0 : part2_io_OutMat_5_0; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_398 = e ? 32'h0 : part2_io_OutMat_5_1; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_399 = e ? 32'h0 : part2_io_OutMat_5_2; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_400 = e ? 32'h0 : part2_io_OutMat_5_3; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_401 = e ? 32'h0 : part2_io_OutMat_5_4; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_402 = e ? 32'h0 : part2_io_OutMat_5_5; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_403 = e ? 32'h0 : part2_io_OutMat_5_6; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_404 = e ? 32'h0 : part2_io_OutMat_5_7; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_405 = e ? 32'h0 : part2_io_OutMat_6_0; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_406 = e ? 32'h0 : part2_io_OutMat_6_1; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_407 = e ? 32'h0 : part2_io_OutMat_6_2; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_408 = e ? 32'h0 : part2_io_OutMat_6_3; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_409 = e ? 32'h0 : part2_io_OutMat_6_4; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_410 = e ? 32'h0 : part2_io_OutMat_6_5; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_411 = e ? 32'h0 : part2_io_OutMat_6_6; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_412 = e ? 32'h0 : part2_io_OutMat_6_7; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_413 = e ? 32'h0 : part2_io_OutMat_7_0; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_414 = e ? 32'h0 : part2_io_OutMat_7_1; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_415 = e ? 32'h0 : part2_io_OutMat_7_2; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_416 = e ? 32'h0 : part2_io_OutMat_7_3; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_417 = e ? 32'h0 : part2_io_OutMat_7_4; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_418 = e ? 32'h0 : part2_io_OutMat_7_5; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_419 = e ? 32'h0 : part2_io_OutMat_7_6; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_420 = e ? 32'h0 : part2_io_OutMat_7_7; // @[DIstribution.scala 102:96 103:16 105:12]
  wire [31:0] _GEN_553 = part2_io_ProcessValid & check ? _GEN_293 : _GEN_357; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_554 = part2_io_ProcessValid & check ? _GEN_294 : _GEN_358; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_555 = part2_io_ProcessValid & check ? _GEN_295 : _GEN_359; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_556 = part2_io_ProcessValid & check ? _GEN_296 : _GEN_360; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_557 = part2_io_ProcessValid & check ? _GEN_297 : _GEN_361; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_558 = part2_io_ProcessValid & check ? _GEN_298 : _GEN_362; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_559 = part2_io_ProcessValid & check ? _GEN_299 : _GEN_363; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_560 = part2_io_ProcessValid & check ? _GEN_300 : _GEN_364; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_561 = part2_io_ProcessValid & check ? _GEN_301 : _GEN_365; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_562 = part2_io_ProcessValid & check ? _GEN_302 : _GEN_366; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_563 = part2_io_ProcessValid & check ? _GEN_303 : _GEN_367; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_564 = part2_io_ProcessValid & check ? _GEN_304 : _GEN_368; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_565 = part2_io_ProcessValid & check ? _GEN_305 : _GEN_369; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_566 = part2_io_ProcessValid & check ? _GEN_306 : _GEN_370; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_567 = part2_io_ProcessValid & check ? _GEN_307 : _GEN_371; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_568 = part2_io_ProcessValid & check ? _GEN_308 : _GEN_372; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_569 = part2_io_ProcessValid & check ? _GEN_309 : _GEN_373; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_570 = part2_io_ProcessValid & check ? _GEN_310 : _GEN_374; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_571 = part2_io_ProcessValid & check ? _GEN_311 : _GEN_375; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_572 = part2_io_ProcessValid & check ? _GEN_312 : _GEN_376; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_573 = part2_io_ProcessValid & check ? _GEN_313 : _GEN_377; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_574 = part2_io_ProcessValid & check ? _GEN_314 : _GEN_378; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_575 = part2_io_ProcessValid & check ? _GEN_315 : _GEN_379; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_576 = part2_io_ProcessValid & check ? _GEN_316 : _GEN_380; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_577 = part2_io_ProcessValid & check ? _GEN_317 : _GEN_381; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_578 = part2_io_ProcessValid & check ? _GEN_318 : _GEN_382; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_579 = part2_io_ProcessValid & check ? _GEN_319 : _GEN_383; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_580 = part2_io_ProcessValid & check ? _GEN_320 : _GEN_384; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_581 = part2_io_ProcessValid & check ? _GEN_321 : _GEN_385; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_582 = part2_io_ProcessValid & check ? _GEN_322 : _GEN_386; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_583 = part2_io_ProcessValid & check ? _GEN_323 : _GEN_387; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_584 = part2_io_ProcessValid & check ? _GEN_324 : _GEN_388; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_585 = part2_io_ProcessValid & check ? _GEN_325 : _GEN_389; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_586 = part2_io_ProcessValid & check ? _GEN_326 : _GEN_390; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_587 = part2_io_ProcessValid & check ? _GEN_327 : _GEN_391; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_588 = part2_io_ProcessValid & check ? _GEN_328 : _GEN_392; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_589 = part2_io_ProcessValid & check ? _GEN_329 : _GEN_393; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_590 = part2_io_ProcessValid & check ? _GEN_330 : _GEN_394; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_591 = part2_io_ProcessValid & check ? _GEN_331 : _GEN_395; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_592 = part2_io_ProcessValid & check ? _GEN_332 : _GEN_396; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_593 = part2_io_ProcessValid & check ? _GEN_333 : _GEN_397; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_594 = part2_io_ProcessValid & check ? _GEN_334 : _GEN_398; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_595 = part2_io_ProcessValid & check ? _GEN_335 : _GEN_399; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_596 = part2_io_ProcessValid & check ? _GEN_336 : _GEN_400; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_597 = part2_io_ProcessValid & check ? _GEN_337 : _GEN_401; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_598 = part2_io_ProcessValid & check ? _GEN_338 : _GEN_402; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_599 = part2_io_ProcessValid & check ? _GEN_339 : _GEN_403; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_600 = part2_io_ProcessValid & check ? _GEN_340 : _GEN_404; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_601 = part2_io_ProcessValid & check ? _GEN_341 : _GEN_405; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_602 = part2_io_ProcessValid & check ? _GEN_342 : _GEN_406; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_603 = part2_io_ProcessValid & check ? _GEN_343 : _GEN_407; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_604 = part2_io_ProcessValid & check ? _GEN_344 : _GEN_408; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_605 = part2_io_ProcessValid & check ? _GEN_345 : _GEN_409; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_606 = part2_io_ProcessValid & check ? _GEN_346 : _GEN_410; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_607 = part2_io_ProcessValid & check ? _GEN_347 : _GEN_411; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_608 = part2_io_ProcessValid & check ? _GEN_348 : _GEN_412; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_609 = part2_io_ProcessValid & check ? _GEN_349 : _GEN_413; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_610 = part2_io_ProcessValid & check ? _GEN_350 : _GEN_414; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_611 = part2_io_ProcessValid & check ? _GEN_351 : _GEN_415; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_612 = part2_io_ProcessValid & check ? _GEN_352 : _GEN_416; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_613 = part2_io_ProcessValid & check ? _GEN_353 : _GEN_417; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_614 = part2_io_ProcessValid & check ? _GEN_354 : _GEN_418; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_615 = part2_io_ProcessValid & check ? _GEN_355 : _GEN_419; // @[DIstribution.scala 82:42]
  wire [31:0] _GEN_616 = part2_io_ProcessValid & check ? _GEN_356 : _GEN_420; // @[DIstribution.scala 82:42]
  wire  _GEN_617 = part2_io_ProcessValid & check ? part3_io_valid : part2_io_Ovalid; // @[DIstribution.scala 106:21 82:42 94:21]
  wire [31:0] _i_T_1 = i + 32'h1; // @[DIstribution.scala 114:16]
  wire  ab = i <= 32'h7 & j < 32'h7; // @[DIstribution.scala 117:42]
  wire [31:0] _j_T_1 = j + 32'h1; // @[DIstribution.scala 120:16]
  abc2 part2 ( // @[DIstribution.scala 55:19]
    .clock(part2_clock),
    .reset(part2_reset),
    .io_IDex(part2_io_IDex),
    .io_JDex(part2_io_JDex),
    .io_valid(part2_io_valid),
    .io_mat_0_0(part2_io_mat_0_0),
    .io_mat_0_1(part2_io_mat_0_1),
    .io_mat_0_2(part2_io_mat_0_2),
    .io_mat_0_3(part2_io_mat_0_3),
    .io_mat_0_4(part2_io_mat_0_4),
    .io_mat_0_5(part2_io_mat_0_5),
    .io_mat_0_6(part2_io_mat_0_6),
    .io_mat_0_7(part2_io_mat_0_7),
    .io_mat_1_0(part2_io_mat_1_0),
    .io_mat_1_1(part2_io_mat_1_1),
    .io_mat_1_2(part2_io_mat_1_2),
    .io_mat_1_3(part2_io_mat_1_3),
    .io_mat_1_4(part2_io_mat_1_4),
    .io_mat_1_5(part2_io_mat_1_5),
    .io_mat_1_6(part2_io_mat_1_6),
    .io_mat_1_7(part2_io_mat_1_7),
    .io_mat_2_0(part2_io_mat_2_0),
    .io_mat_2_1(part2_io_mat_2_1),
    .io_mat_2_2(part2_io_mat_2_2),
    .io_mat_2_3(part2_io_mat_2_3),
    .io_mat_2_4(part2_io_mat_2_4),
    .io_mat_2_5(part2_io_mat_2_5),
    .io_mat_2_6(part2_io_mat_2_6),
    .io_mat_2_7(part2_io_mat_2_7),
    .io_mat_3_0(part2_io_mat_3_0),
    .io_mat_3_1(part2_io_mat_3_1),
    .io_mat_3_2(part2_io_mat_3_2),
    .io_mat_3_3(part2_io_mat_3_3),
    .io_mat_3_4(part2_io_mat_3_4),
    .io_mat_3_5(part2_io_mat_3_5),
    .io_mat_3_6(part2_io_mat_3_6),
    .io_mat_3_7(part2_io_mat_3_7),
    .io_mat_4_0(part2_io_mat_4_0),
    .io_mat_4_1(part2_io_mat_4_1),
    .io_mat_4_2(part2_io_mat_4_2),
    .io_mat_4_3(part2_io_mat_4_3),
    .io_mat_4_4(part2_io_mat_4_4),
    .io_mat_4_5(part2_io_mat_4_5),
    .io_mat_4_6(part2_io_mat_4_6),
    .io_mat_4_7(part2_io_mat_4_7),
    .io_mat_5_0(part2_io_mat_5_0),
    .io_mat_5_1(part2_io_mat_5_1),
    .io_mat_5_2(part2_io_mat_5_2),
    .io_mat_5_3(part2_io_mat_5_3),
    .io_mat_5_4(part2_io_mat_5_4),
    .io_mat_5_5(part2_io_mat_5_5),
    .io_mat_5_6(part2_io_mat_5_6),
    .io_mat_5_7(part2_io_mat_5_7),
    .io_mat_6_0(part2_io_mat_6_0),
    .io_mat_6_1(part2_io_mat_6_1),
    .io_mat_6_2(part2_io_mat_6_2),
    .io_mat_6_3(part2_io_mat_6_3),
    .io_mat_6_4(part2_io_mat_6_4),
    .io_mat_6_5(part2_io_mat_6_5),
    .io_mat_6_6(part2_io_mat_6_6),
    .io_mat_6_7(part2_io_mat_6_7),
    .io_mat_7_0(part2_io_mat_7_0),
    .io_mat_7_1(part2_io_mat_7_1),
    .io_mat_7_2(part2_io_mat_7_2),
    .io_mat_7_3(part2_io_mat_7_3),
    .io_mat_7_4(part2_io_mat_7_4),
    .io_mat_7_5(part2_io_mat_7_5),
    .io_mat_7_6(part2_io_mat_7_6),
    .io_mat_7_7(part2_io_mat_7_7),
    .io_OutMat_0_0(part2_io_OutMat_0_0),
    .io_OutMat_0_1(part2_io_OutMat_0_1),
    .io_OutMat_0_2(part2_io_OutMat_0_2),
    .io_OutMat_0_3(part2_io_OutMat_0_3),
    .io_OutMat_0_4(part2_io_OutMat_0_4),
    .io_OutMat_0_5(part2_io_OutMat_0_5),
    .io_OutMat_0_6(part2_io_OutMat_0_6),
    .io_OutMat_0_7(part2_io_OutMat_0_7),
    .io_OutMat_1_0(part2_io_OutMat_1_0),
    .io_OutMat_1_1(part2_io_OutMat_1_1),
    .io_OutMat_1_2(part2_io_OutMat_1_2),
    .io_OutMat_1_3(part2_io_OutMat_1_3),
    .io_OutMat_1_4(part2_io_OutMat_1_4),
    .io_OutMat_1_5(part2_io_OutMat_1_5),
    .io_OutMat_1_6(part2_io_OutMat_1_6),
    .io_OutMat_1_7(part2_io_OutMat_1_7),
    .io_OutMat_2_0(part2_io_OutMat_2_0),
    .io_OutMat_2_1(part2_io_OutMat_2_1),
    .io_OutMat_2_2(part2_io_OutMat_2_2),
    .io_OutMat_2_3(part2_io_OutMat_2_3),
    .io_OutMat_2_4(part2_io_OutMat_2_4),
    .io_OutMat_2_5(part2_io_OutMat_2_5),
    .io_OutMat_2_6(part2_io_OutMat_2_6),
    .io_OutMat_2_7(part2_io_OutMat_2_7),
    .io_OutMat_3_0(part2_io_OutMat_3_0),
    .io_OutMat_3_1(part2_io_OutMat_3_1),
    .io_OutMat_3_2(part2_io_OutMat_3_2),
    .io_OutMat_3_3(part2_io_OutMat_3_3),
    .io_OutMat_3_4(part2_io_OutMat_3_4),
    .io_OutMat_3_5(part2_io_OutMat_3_5),
    .io_OutMat_3_6(part2_io_OutMat_3_6),
    .io_OutMat_3_7(part2_io_OutMat_3_7),
    .io_OutMat_4_0(part2_io_OutMat_4_0),
    .io_OutMat_4_1(part2_io_OutMat_4_1),
    .io_OutMat_4_2(part2_io_OutMat_4_2),
    .io_OutMat_4_3(part2_io_OutMat_4_3),
    .io_OutMat_4_4(part2_io_OutMat_4_4),
    .io_OutMat_4_5(part2_io_OutMat_4_5),
    .io_OutMat_4_6(part2_io_OutMat_4_6),
    .io_OutMat_4_7(part2_io_OutMat_4_7),
    .io_OutMat_5_0(part2_io_OutMat_5_0),
    .io_OutMat_5_1(part2_io_OutMat_5_1),
    .io_OutMat_5_2(part2_io_OutMat_5_2),
    .io_OutMat_5_3(part2_io_OutMat_5_3),
    .io_OutMat_5_4(part2_io_OutMat_5_4),
    .io_OutMat_5_5(part2_io_OutMat_5_5),
    .io_OutMat_5_6(part2_io_OutMat_5_6),
    .io_OutMat_5_7(part2_io_OutMat_5_7),
    .io_OutMat_6_0(part2_io_OutMat_6_0),
    .io_OutMat_6_1(part2_io_OutMat_6_1),
    .io_OutMat_6_2(part2_io_OutMat_6_2),
    .io_OutMat_6_3(part2_io_OutMat_6_3),
    .io_OutMat_6_4(part2_io_OutMat_6_4),
    .io_OutMat_6_5(part2_io_OutMat_6_5),
    .io_OutMat_6_6(part2_io_OutMat_6_6),
    .io_OutMat_6_7(part2_io_OutMat_6_7),
    .io_OutMat_7_0(part2_io_OutMat_7_0),
    .io_OutMat_7_1(part2_io_OutMat_7_1),
    .io_OutMat_7_2(part2_io_OutMat_7_2),
    .io_OutMat_7_3(part2_io_OutMat_7_3),
    .io_OutMat_7_4(part2_io_OutMat_7_4),
    .io_OutMat_7_5(part2_io_OutMat_7_5),
    .io_OutMat_7_6(part2_io_OutMat_7_6),
    .io_OutMat_7_7(part2_io_OutMat_7_7),
    .io_Ovalid(part2_io_Ovalid),
    .io_ProcessValid(part2_io_ProcessValid)
  );
  abc3 part3 ( // @[DIstribution.scala 69:23]
    .clock(part3_clock),
    .reset(part3_reset),
    .io_PreMat_0_0(part3_io_PreMat_0_0),
    .io_PreMat_0_1(part3_io_PreMat_0_1),
    .io_PreMat_0_2(part3_io_PreMat_0_2),
    .io_PreMat_0_3(part3_io_PreMat_0_3),
    .io_PreMat_0_4(part3_io_PreMat_0_4),
    .io_PreMat_0_5(part3_io_PreMat_0_5),
    .io_PreMat_0_6(part3_io_PreMat_0_6),
    .io_PreMat_0_7(part3_io_PreMat_0_7),
    .io_PreMat_1_0(part3_io_PreMat_1_0),
    .io_PreMat_1_1(part3_io_PreMat_1_1),
    .io_PreMat_1_2(part3_io_PreMat_1_2),
    .io_PreMat_1_3(part3_io_PreMat_1_3),
    .io_PreMat_1_4(part3_io_PreMat_1_4),
    .io_PreMat_1_5(part3_io_PreMat_1_5),
    .io_PreMat_1_6(part3_io_PreMat_1_6),
    .io_PreMat_1_7(part3_io_PreMat_1_7),
    .io_PreMat_2_0(part3_io_PreMat_2_0),
    .io_PreMat_2_1(part3_io_PreMat_2_1),
    .io_PreMat_2_2(part3_io_PreMat_2_2),
    .io_PreMat_2_3(part3_io_PreMat_2_3),
    .io_PreMat_2_4(part3_io_PreMat_2_4),
    .io_PreMat_2_5(part3_io_PreMat_2_5),
    .io_PreMat_2_6(part3_io_PreMat_2_6),
    .io_PreMat_2_7(part3_io_PreMat_2_7),
    .io_PreMat_3_0(part3_io_PreMat_3_0),
    .io_PreMat_3_1(part3_io_PreMat_3_1),
    .io_PreMat_3_2(part3_io_PreMat_3_2),
    .io_PreMat_3_3(part3_io_PreMat_3_3),
    .io_PreMat_3_4(part3_io_PreMat_3_4),
    .io_PreMat_3_5(part3_io_PreMat_3_5),
    .io_PreMat_3_6(part3_io_PreMat_3_6),
    .io_PreMat_3_7(part3_io_PreMat_3_7),
    .io_PreMat_4_0(part3_io_PreMat_4_0),
    .io_PreMat_4_1(part3_io_PreMat_4_1),
    .io_PreMat_4_2(part3_io_PreMat_4_2),
    .io_PreMat_4_3(part3_io_PreMat_4_3),
    .io_PreMat_4_4(part3_io_PreMat_4_4),
    .io_PreMat_4_5(part3_io_PreMat_4_5),
    .io_PreMat_4_6(part3_io_PreMat_4_6),
    .io_PreMat_4_7(part3_io_PreMat_4_7),
    .io_PreMat_5_0(part3_io_PreMat_5_0),
    .io_PreMat_5_1(part3_io_PreMat_5_1),
    .io_PreMat_5_2(part3_io_PreMat_5_2),
    .io_PreMat_5_3(part3_io_PreMat_5_3),
    .io_PreMat_5_4(part3_io_PreMat_5_4),
    .io_PreMat_5_5(part3_io_PreMat_5_5),
    .io_PreMat_5_6(part3_io_PreMat_5_6),
    .io_PreMat_5_7(part3_io_PreMat_5_7),
    .io_PreMat_6_0(part3_io_PreMat_6_0),
    .io_PreMat_6_1(part3_io_PreMat_6_1),
    .io_PreMat_6_2(part3_io_PreMat_6_2),
    .io_PreMat_6_3(part3_io_PreMat_6_3),
    .io_PreMat_6_4(part3_io_PreMat_6_4),
    .io_PreMat_6_5(part3_io_PreMat_6_5),
    .io_PreMat_6_6(part3_io_PreMat_6_6),
    .io_PreMat_6_7(part3_io_PreMat_6_7),
    .io_PreMat_7_0(part3_io_PreMat_7_0),
    .io_PreMat_7_1(part3_io_PreMat_7_1),
    .io_PreMat_7_2(part3_io_PreMat_7_2),
    .io_PreMat_7_3(part3_io_PreMat_7_3),
    .io_PreMat_7_4(part3_io_PreMat_7_4),
    .io_PreMat_7_5(part3_io_PreMat_7_5),
    .io_PreMat_7_6(part3_io_PreMat_7_6),
    .io_PreMat_7_7(part3_io_PreMat_7_7),
    .io_IDex(part3_io_IDex),
    .io_mat_0_0(part3_io_mat_0_0),
    .io_mat_0_1(part3_io_mat_0_1),
    .io_mat_0_2(part3_io_mat_0_2),
    .io_mat_0_3(part3_io_mat_0_3),
    .io_mat_0_4(part3_io_mat_0_4),
    .io_mat_0_5(part3_io_mat_0_5),
    .io_mat_0_6(part3_io_mat_0_6),
    .io_mat_0_7(part3_io_mat_0_7),
    .io_mat_1_0(part3_io_mat_1_0),
    .io_mat_1_1(part3_io_mat_1_1),
    .io_mat_1_2(part3_io_mat_1_2),
    .io_mat_1_3(part3_io_mat_1_3),
    .io_mat_1_4(part3_io_mat_1_4),
    .io_mat_1_5(part3_io_mat_1_5),
    .io_mat_1_6(part3_io_mat_1_6),
    .io_mat_1_7(part3_io_mat_1_7),
    .io_mat_2_0(part3_io_mat_2_0),
    .io_mat_2_1(part3_io_mat_2_1),
    .io_mat_2_2(part3_io_mat_2_2),
    .io_mat_2_3(part3_io_mat_2_3),
    .io_mat_2_4(part3_io_mat_2_4),
    .io_mat_2_5(part3_io_mat_2_5),
    .io_mat_2_6(part3_io_mat_2_6),
    .io_mat_2_7(part3_io_mat_2_7),
    .io_mat_3_0(part3_io_mat_3_0),
    .io_mat_3_1(part3_io_mat_3_1),
    .io_mat_3_2(part3_io_mat_3_2),
    .io_mat_3_3(part3_io_mat_3_3),
    .io_mat_3_4(part3_io_mat_3_4),
    .io_mat_3_5(part3_io_mat_3_5),
    .io_mat_3_6(part3_io_mat_3_6),
    .io_mat_3_7(part3_io_mat_3_7),
    .io_mat_4_0(part3_io_mat_4_0),
    .io_mat_4_1(part3_io_mat_4_1),
    .io_mat_4_2(part3_io_mat_4_2),
    .io_mat_4_3(part3_io_mat_4_3),
    .io_mat_4_4(part3_io_mat_4_4),
    .io_mat_4_5(part3_io_mat_4_5),
    .io_mat_4_6(part3_io_mat_4_6),
    .io_mat_4_7(part3_io_mat_4_7),
    .io_mat_5_0(part3_io_mat_5_0),
    .io_mat_5_1(part3_io_mat_5_1),
    .io_mat_5_2(part3_io_mat_5_2),
    .io_mat_5_3(part3_io_mat_5_3),
    .io_mat_5_4(part3_io_mat_5_4),
    .io_mat_5_5(part3_io_mat_5_5),
    .io_mat_5_6(part3_io_mat_5_6),
    .io_mat_5_7(part3_io_mat_5_7),
    .io_mat_6_0(part3_io_mat_6_0),
    .io_mat_6_1(part3_io_mat_6_1),
    .io_mat_6_2(part3_io_mat_6_2),
    .io_mat_6_3(part3_io_mat_6_3),
    .io_mat_6_4(part3_io_mat_6_4),
    .io_mat_6_5(part3_io_mat_6_5),
    .io_mat_6_6(part3_io_mat_6_6),
    .io_mat_6_7(part3_io_mat_6_7),
    .io_mat_7_0(part3_io_mat_7_0),
    .io_mat_7_1(part3_io_mat_7_1),
    .io_mat_7_2(part3_io_mat_7_2),
    .io_mat_7_3(part3_io_mat_7_3),
    .io_mat_7_4(part3_io_mat_7_4),
    .io_mat_7_5(part3_io_mat_7_5),
    .io_mat_7_6(part3_io_mat_7_6),
    .io_mat_7_7(part3_io_mat_7_7),
    .io_i_valid(part3_io_i_valid),
    .io_valid(part3_io_valid),
    .io_Omat_0_0(part3_io_Omat_0_0),
    .io_Omat_0_1(part3_io_Omat_0_1),
    .io_Omat_0_2(part3_io_Omat_0_2),
    .io_Omat_0_3(part3_io_Omat_0_3),
    .io_Omat_0_4(part3_io_Omat_0_4),
    .io_Omat_0_5(part3_io_Omat_0_5),
    .io_Omat_0_6(part3_io_Omat_0_6),
    .io_Omat_0_7(part3_io_Omat_0_7),
    .io_Omat_1_0(part3_io_Omat_1_0),
    .io_Omat_1_1(part3_io_Omat_1_1),
    .io_Omat_1_2(part3_io_Omat_1_2),
    .io_Omat_1_3(part3_io_Omat_1_3),
    .io_Omat_1_4(part3_io_Omat_1_4),
    .io_Omat_1_5(part3_io_Omat_1_5),
    .io_Omat_1_6(part3_io_Omat_1_6),
    .io_Omat_1_7(part3_io_Omat_1_7),
    .io_Omat_2_0(part3_io_Omat_2_0),
    .io_Omat_2_1(part3_io_Omat_2_1),
    .io_Omat_2_2(part3_io_Omat_2_2),
    .io_Omat_2_3(part3_io_Omat_2_3),
    .io_Omat_2_4(part3_io_Omat_2_4),
    .io_Omat_2_5(part3_io_Omat_2_5),
    .io_Omat_2_6(part3_io_Omat_2_6),
    .io_Omat_2_7(part3_io_Omat_2_7),
    .io_Omat_3_0(part3_io_Omat_3_0),
    .io_Omat_3_1(part3_io_Omat_3_1),
    .io_Omat_3_2(part3_io_Omat_3_2),
    .io_Omat_3_3(part3_io_Omat_3_3),
    .io_Omat_3_4(part3_io_Omat_3_4),
    .io_Omat_3_5(part3_io_Omat_3_5),
    .io_Omat_3_6(part3_io_Omat_3_6),
    .io_Omat_3_7(part3_io_Omat_3_7),
    .io_Omat_4_0(part3_io_Omat_4_0),
    .io_Omat_4_1(part3_io_Omat_4_1),
    .io_Omat_4_2(part3_io_Omat_4_2),
    .io_Omat_4_3(part3_io_Omat_4_3),
    .io_Omat_4_4(part3_io_Omat_4_4),
    .io_Omat_4_5(part3_io_Omat_4_5),
    .io_Omat_4_6(part3_io_Omat_4_6),
    .io_Omat_4_7(part3_io_Omat_4_7),
    .io_Omat_5_0(part3_io_Omat_5_0),
    .io_Omat_5_1(part3_io_Omat_5_1),
    .io_Omat_5_2(part3_io_Omat_5_2),
    .io_Omat_5_3(part3_io_Omat_5_3),
    .io_Omat_5_4(part3_io_Omat_5_4),
    .io_Omat_5_5(part3_io_Omat_5_5),
    .io_Omat_5_6(part3_io_Omat_5_6),
    .io_Omat_5_7(part3_io_Omat_5_7),
    .io_Omat_6_0(part3_io_Omat_6_0),
    .io_Omat_6_1(part3_io_Omat_6_1),
    .io_Omat_6_2(part3_io_Omat_6_2),
    .io_Omat_6_3(part3_io_Omat_6_3),
    .io_Omat_6_4(part3_io_Omat_6_4),
    .io_Omat_6_5(part3_io_Omat_6_5),
    .io_Omat_6_6(part3_io_Omat_6_6),
    .io_Omat_6_7(part3_io_Omat_6_7),
    .io_Omat_7_0(part3_io_Omat_7_0),
    .io_Omat_7_1(part3_io_Omat_7_1),
    .io_Omat_7_2(part3_io_Omat_7_2),
    .io_Omat_7_3(part3_io_Omat_7_3),
    .io_Omat_7_4(part3_io_Omat_7_4),
    .io_Omat_7_5(part3_io_Omat_7_5),
    .io_Omat_7_6(part3_io_Omat_7_6),
    .io_Omat_7_7(part3_io_Omat_7_7),
    .io_merge(part3_io_merge)
  );
  assign io_out_0_0 = io_valid ? _GEN_553 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_0_1 = io_valid ? _GEN_554 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_0_2 = io_valid ? _GEN_555 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_0_3 = io_valid ? _GEN_556 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_0_4 = io_valid ? _GEN_557 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_0_5 = io_valid ? _GEN_558 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_0_6 = io_valid ? _GEN_559 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_0_7 = io_valid ? _GEN_560 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_1_0 = io_valid ? _GEN_561 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_1_1 = io_valid ? _GEN_562 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_1_2 = io_valid ? _GEN_563 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_1_3 = io_valid ? _GEN_564 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_1_4 = io_valid ? _GEN_565 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_1_5 = io_valid ? _GEN_566 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_1_6 = io_valid ? _GEN_567 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_1_7 = io_valid ? _GEN_568 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_2_0 = io_valid ? _GEN_569 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_2_1 = io_valid ? _GEN_570 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_2_2 = io_valid ? _GEN_571 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_2_3 = io_valid ? _GEN_572 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_2_4 = io_valid ? _GEN_573 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_2_5 = io_valid ? _GEN_574 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_2_6 = io_valid ? _GEN_575 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_2_7 = io_valid ? _GEN_576 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_3_0 = io_valid ? _GEN_577 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_3_1 = io_valid ? _GEN_578 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_3_2 = io_valid ? _GEN_579 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_3_3 = io_valid ? _GEN_580 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_3_4 = io_valid ? _GEN_581 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_3_5 = io_valid ? _GEN_582 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_3_6 = io_valid ? _GEN_583 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_3_7 = io_valid ? _GEN_584 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_4_0 = io_valid ? _GEN_585 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_4_1 = io_valid ? _GEN_586 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_4_2 = io_valid ? _GEN_587 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_4_3 = io_valid ? _GEN_588 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_4_4 = io_valid ? _GEN_589 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_4_5 = io_valid ? _GEN_590 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_4_6 = io_valid ? _GEN_591 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_4_7 = io_valid ? _GEN_592 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_5_0 = io_valid ? _GEN_593 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_5_1 = io_valid ? _GEN_594 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_5_2 = io_valid ? _GEN_595 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_5_3 = io_valid ? _GEN_596 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_5_4 = io_valid ? _GEN_597 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_5_5 = io_valid ? _GEN_598 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_5_6 = io_valid ? _GEN_599 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_5_7 = io_valid ? _GEN_600 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_6_0 = io_valid ? _GEN_601 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_6_1 = io_valid ? _GEN_602 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_6_2 = io_valid ? _GEN_603 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_6_3 = io_valid ? _GEN_604 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_6_4 = io_valid ? _GEN_605 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_6_5 = io_valid ? _GEN_606 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_6_6 = io_valid ? _GEN_607 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_6_7 = io_valid ? _GEN_608 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_7_0 = io_valid ? _GEN_609 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_7_1 = io_valid ? _GEN_610 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_7_2 = io_valid ? _GEN_611 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_7_3 = io_valid ? _GEN_612 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_7_4 = io_valid ? _GEN_613 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_7_5 = io_valid ? _GEN_614 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_7_6 = io_valid ? _GEN_615 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_out_7_7 = io_valid ? _GEN_616 : 32'h0; // @[DIstribution.scala 131:16 27:21]
  assign io_ProcessValid = io_valid & _GEN_617; // @[DIstribution.scala 27:21 132:25]
  assign part2_clock = clock;
  assign part2_reset = reset;
  assign part2_io_IDex = c ? _GEN_265 : 32'h0; // @[DIstribution.scala 59:13 60:19 63:19]
  assign part2_io_JDex = c ? _GEN_273 : 32'h0; // @[DIstribution.scala 59:13 61:19 64:19]
  assign part2_io_valid = c; // @[DIstribution.scala 58:20]
  assign part2_io_mat_0_0 = io_matrix_0_0; // @[DIstribution.scala 56:14]
  assign part2_io_mat_0_1 = io_matrix_0_1; // @[DIstribution.scala 56:14]
  assign part2_io_mat_0_2 = io_matrix_0_2; // @[DIstribution.scala 56:14]
  assign part2_io_mat_0_3 = io_matrix_0_3; // @[DIstribution.scala 56:14]
  assign part2_io_mat_0_4 = io_matrix_0_4; // @[DIstribution.scala 56:14]
  assign part2_io_mat_0_5 = io_matrix_0_5; // @[DIstribution.scala 56:14]
  assign part2_io_mat_0_6 = io_matrix_0_6; // @[DIstribution.scala 56:14]
  assign part2_io_mat_0_7 = io_matrix_0_7; // @[DIstribution.scala 56:14]
  assign part2_io_mat_1_0 = io_matrix_1_0; // @[DIstribution.scala 56:14]
  assign part2_io_mat_1_1 = io_matrix_1_1; // @[DIstribution.scala 56:14]
  assign part2_io_mat_1_2 = io_matrix_1_2; // @[DIstribution.scala 56:14]
  assign part2_io_mat_1_3 = io_matrix_1_3; // @[DIstribution.scala 56:14]
  assign part2_io_mat_1_4 = io_matrix_1_4; // @[DIstribution.scala 56:14]
  assign part2_io_mat_1_5 = io_matrix_1_5; // @[DIstribution.scala 56:14]
  assign part2_io_mat_1_6 = io_matrix_1_6; // @[DIstribution.scala 56:14]
  assign part2_io_mat_1_7 = io_matrix_1_7; // @[DIstribution.scala 56:14]
  assign part2_io_mat_2_0 = io_matrix_2_0; // @[DIstribution.scala 56:14]
  assign part2_io_mat_2_1 = io_matrix_2_1; // @[DIstribution.scala 56:14]
  assign part2_io_mat_2_2 = io_matrix_2_2; // @[DIstribution.scala 56:14]
  assign part2_io_mat_2_3 = io_matrix_2_3; // @[DIstribution.scala 56:14]
  assign part2_io_mat_2_4 = io_matrix_2_4; // @[DIstribution.scala 56:14]
  assign part2_io_mat_2_5 = io_matrix_2_5; // @[DIstribution.scala 56:14]
  assign part2_io_mat_2_6 = io_matrix_2_6; // @[DIstribution.scala 56:14]
  assign part2_io_mat_2_7 = io_matrix_2_7; // @[DIstribution.scala 56:14]
  assign part2_io_mat_3_0 = io_matrix_3_0; // @[DIstribution.scala 56:14]
  assign part2_io_mat_3_1 = io_matrix_3_1; // @[DIstribution.scala 56:14]
  assign part2_io_mat_3_2 = io_matrix_3_2; // @[DIstribution.scala 56:14]
  assign part2_io_mat_3_3 = io_matrix_3_3; // @[DIstribution.scala 56:14]
  assign part2_io_mat_3_4 = io_matrix_3_4; // @[DIstribution.scala 56:14]
  assign part2_io_mat_3_5 = io_matrix_3_5; // @[DIstribution.scala 56:14]
  assign part2_io_mat_3_6 = io_matrix_3_6; // @[DIstribution.scala 56:14]
  assign part2_io_mat_3_7 = io_matrix_3_7; // @[DIstribution.scala 56:14]
  assign part2_io_mat_4_0 = io_matrix_4_0; // @[DIstribution.scala 56:14]
  assign part2_io_mat_4_1 = io_matrix_4_1; // @[DIstribution.scala 56:14]
  assign part2_io_mat_4_2 = io_matrix_4_2; // @[DIstribution.scala 56:14]
  assign part2_io_mat_4_3 = io_matrix_4_3; // @[DIstribution.scala 56:14]
  assign part2_io_mat_4_4 = io_matrix_4_4; // @[DIstribution.scala 56:14]
  assign part2_io_mat_4_5 = io_matrix_4_5; // @[DIstribution.scala 56:14]
  assign part2_io_mat_4_6 = io_matrix_4_6; // @[DIstribution.scala 56:14]
  assign part2_io_mat_4_7 = io_matrix_4_7; // @[DIstribution.scala 56:14]
  assign part2_io_mat_5_0 = io_matrix_5_0; // @[DIstribution.scala 56:14]
  assign part2_io_mat_5_1 = io_matrix_5_1; // @[DIstribution.scala 56:14]
  assign part2_io_mat_5_2 = io_matrix_5_2; // @[DIstribution.scala 56:14]
  assign part2_io_mat_5_3 = io_matrix_5_3; // @[DIstribution.scala 56:14]
  assign part2_io_mat_5_4 = io_matrix_5_4; // @[DIstribution.scala 56:14]
  assign part2_io_mat_5_5 = io_matrix_5_5; // @[DIstribution.scala 56:14]
  assign part2_io_mat_5_6 = io_matrix_5_6; // @[DIstribution.scala 56:14]
  assign part2_io_mat_5_7 = io_matrix_5_7; // @[DIstribution.scala 56:14]
  assign part2_io_mat_6_0 = io_matrix_6_0; // @[DIstribution.scala 56:14]
  assign part2_io_mat_6_1 = io_matrix_6_1; // @[DIstribution.scala 56:14]
  assign part2_io_mat_6_2 = io_matrix_6_2; // @[DIstribution.scala 56:14]
  assign part2_io_mat_6_3 = io_matrix_6_3; // @[DIstribution.scala 56:14]
  assign part2_io_mat_6_4 = io_matrix_6_4; // @[DIstribution.scala 56:14]
  assign part2_io_mat_6_5 = io_matrix_6_5; // @[DIstribution.scala 56:14]
  assign part2_io_mat_6_6 = io_matrix_6_6; // @[DIstribution.scala 56:14]
  assign part2_io_mat_6_7 = io_matrix_6_7; // @[DIstribution.scala 56:14]
  assign part2_io_mat_7_0 = io_matrix_7_0; // @[DIstribution.scala 56:14]
  assign part2_io_mat_7_1 = io_matrix_7_1; // @[DIstribution.scala 56:14]
  assign part2_io_mat_7_2 = io_matrix_7_2; // @[DIstribution.scala 56:14]
  assign part2_io_mat_7_3 = io_matrix_7_3; // @[DIstribution.scala 56:14]
  assign part2_io_mat_7_4 = io_matrix_7_4; // @[DIstribution.scala 56:14]
  assign part2_io_mat_7_5 = io_matrix_7_5; // @[DIstribution.scala 56:14]
  assign part2_io_mat_7_6 = io_matrix_7_6; // @[DIstribution.scala 56:14]
  assign part2_io_mat_7_7 = io_matrix_7_7; // @[DIstribution.scala 56:14]
  assign part3_clock = clock;
  assign part3_reset = reset;
  assign part3_io_PreMat_0_0 = part2_io_ProcessValid & check ? part2_io_OutMat_0_0 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_0_1 = part2_io_ProcessValid & check ? part2_io_OutMat_0_1 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_0_2 = part2_io_ProcessValid & check ? part2_io_OutMat_0_2 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_0_3 = part2_io_ProcessValid & check ? part2_io_OutMat_0_3 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_0_4 = part2_io_ProcessValid & check ? part2_io_OutMat_0_4 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_0_5 = part2_io_ProcessValid & check ? part2_io_OutMat_0_5 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_0_6 = part2_io_ProcessValid & check ? part2_io_OutMat_0_6 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_0_7 = part2_io_ProcessValid & check ? part2_io_OutMat_0_7 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_1_0 = part2_io_ProcessValid & check ? part2_io_OutMat_1_0 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_1_1 = part2_io_ProcessValid & check ? part2_io_OutMat_1_1 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_1_2 = part2_io_ProcessValid & check ? part2_io_OutMat_1_2 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_1_3 = part2_io_ProcessValid & check ? part2_io_OutMat_1_3 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_1_4 = part2_io_ProcessValid & check ? part2_io_OutMat_1_4 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_1_5 = part2_io_ProcessValid & check ? part2_io_OutMat_1_5 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_1_6 = part2_io_ProcessValid & check ? part2_io_OutMat_1_6 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_1_7 = part2_io_ProcessValid & check ? part2_io_OutMat_1_7 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_2_0 = part2_io_ProcessValid & check ? part2_io_OutMat_2_0 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_2_1 = part2_io_ProcessValid & check ? part2_io_OutMat_2_1 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_2_2 = part2_io_ProcessValid & check ? part2_io_OutMat_2_2 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_2_3 = part2_io_ProcessValid & check ? part2_io_OutMat_2_3 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_2_4 = part2_io_ProcessValid & check ? part2_io_OutMat_2_4 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_2_5 = part2_io_ProcessValid & check ? part2_io_OutMat_2_5 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_2_6 = part2_io_ProcessValid & check ? part2_io_OutMat_2_6 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_2_7 = part2_io_ProcessValid & check ? part2_io_OutMat_2_7 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_3_0 = part2_io_ProcessValid & check ? part2_io_OutMat_3_0 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_3_1 = part2_io_ProcessValid & check ? part2_io_OutMat_3_1 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_3_2 = part2_io_ProcessValid & check ? part2_io_OutMat_3_2 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_3_3 = part2_io_ProcessValid & check ? part2_io_OutMat_3_3 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_3_4 = part2_io_ProcessValid & check ? part2_io_OutMat_3_4 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_3_5 = part2_io_ProcessValid & check ? part2_io_OutMat_3_5 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_3_6 = part2_io_ProcessValid & check ? part2_io_OutMat_3_6 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_3_7 = part2_io_ProcessValid & check ? part2_io_OutMat_3_7 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_4_0 = part2_io_ProcessValid & check ? part2_io_OutMat_4_0 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_4_1 = part2_io_ProcessValid & check ? part2_io_OutMat_4_1 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_4_2 = part2_io_ProcessValid & check ? part2_io_OutMat_4_2 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_4_3 = part2_io_ProcessValid & check ? part2_io_OutMat_4_3 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_4_4 = part2_io_ProcessValid & check ? part2_io_OutMat_4_4 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_4_5 = part2_io_ProcessValid & check ? part2_io_OutMat_4_5 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_4_6 = part2_io_ProcessValid & check ? part2_io_OutMat_4_6 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_4_7 = part2_io_ProcessValid & check ? part2_io_OutMat_4_7 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_5_0 = part2_io_ProcessValid & check ? part2_io_OutMat_5_0 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_5_1 = part2_io_ProcessValid & check ? part2_io_OutMat_5_1 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_5_2 = part2_io_ProcessValid & check ? part2_io_OutMat_5_2 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_5_3 = part2_io_ProcessValid & check ? part2_io_OutMat_5_3 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_5_4 = part2_io_ProcessValid & check ? part2_io_OutMat_5_4 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_5_5 = part2_io_ProcessValid & check ? part2_io_OutMat_5_5 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_5_6 = part2_io_ProcessValid & check ? part2_io_OutMat_5_6 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_5_7 = part2_io_ProcessValid & check ? part2_io_OutMat_5_7 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_6_0 = part2_io_ProcessValid & check ? part2_io_OutMat_6_0 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_6_1 = part2_io_ProcessValid & check ? part2_io_OutMat_6_1 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_6_2 = part2_io_ProcessValid & check ? part2_io_OutMat_6_2 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_6_3 = part2_io_ProcessValid & check ? part2_io_OutMat_6_3 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_6_4 = part2_io_ProcessValid & check ? part2_io_OutMat_6_4 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_6_5 = part2_io_ProcessValid & check ? part2_io_OutMat_6_5 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_6_6 = part2_io_ProcessValid & check ? part2_io_OutMat_6_6 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_6_7 = part2_io_ProcessValid & check ? part2_io_OutMat_6_7 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_7_0 = part2_io_ProcessValid & check ? part2_io_OutMat_7_0 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_7_1 = part2_io_ProcessValid & check ? part2_io_OutMat_7_1 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_7_2 = part2_io_ProcessValid & check ? part2_io_OutMat_7_2 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_7_3 = part2_io_ProcessValid & check ? part2_io_OutMat_7_3 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_7_4 = part2_io_ProcessValid & check ? part2_io_OutMat_7_4 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_7_5 = part2_io_ProcessValid & check ? part2_io_OutMat_7_5 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_7_6 = part2_io_ProcessValid & check ? part2_io_OutMat_7_6 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_PreMat_7_7 = part2_io_ProcessValid & check ? part2_io_OutMat_7_7 : 32'h0; // @[DIstribution.scala 82:42 86:21 99:21]
  assign part3_io_IDex = part2_io_ProcessValid & check ? _GEN_265 : 32'h0; // @[DIstribution.scala 100:19 82:42 88:19]
  assign part3_io_mat_0_0 = part2_io_ProcessValid & check ? io_matrix_0_0 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_0_1 = part2_io_ProcessValid & check ? io_matrix_0_1 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_0_2 = part2_io_ProcessValid & check ? io_matrix_0_2 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_0_3 = part2_io_ProcessValid & check ? io_matrix_0_3 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_0_4 = part2_io_ProcessValid & check ? io_matrix_0_4 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_0_5 = part2_io_ProcessValid & check ? io_matrix_0_5 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_0_6 = part2_io_ProcessValid & check ? io_matrix_0_6 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_0_7 = part2_io_ProcessValid & check ? io_matrix_0_7 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_1_0 = part2_io_ProcessValid & check ? io_matrix_1_0 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_1_1 = part2_io_ProcessValid & check ? io_matrix_1_1 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_1_2 = part2_io_ProcessValid & check ? io_matrix_1_2 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_1_3 = part2_io_ProcessValid & check ? io_matrix_1_3 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_1_4 = part2_io_ProcessValid & check ? io_matrix_1_4 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_1_5 = part2_io_ProcessValid & check ? io_matrix_1_5 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_1_6 = part2_io_ProcessValid & check ? io_matrix_1_6 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_1_7 = part2_io_ProcessValid & check ? io_matrix_1_7 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_2_0 = part2_io_ProcessValid & check ? io_matrix_2_0 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_2_1 = part2_io_ProcessValid & check ? io_matrix_2_1 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_2_2 = part2_io_ProcessValid & check ? io_matrix_2_2 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_2_3 = part2_io_ProcessValid & check ? io_matrix_2_3 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_2_4 = part2_io_ProcessValid & check ? io_matrix_2_4 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_2_5 = part2_io_ProcessValid & check ? io_matrix_2_5 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_2_6 = part2_io_ProcessValid & check ? io_matrix_2_6 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_2_7 = part2_io_ProcessValid & check ? io_matrix_2_7 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_3_0 = part2_io_ProcessValid & check ? io_matrix_3_0 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_3_1 = part2_io_ProcessValid & check ? io_matrix_3_1 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_3_2 = part2_io_ProcessValid & check ? io_matrix_3_2 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_3_3 = part2_io_ProcessValid & check ? io_matrix_3_3 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_3_4 = part2_io_ProcessValid & check ? io_matrix_3_4 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_3_5 = part2_io_ProcessValid & check ? io_matrix_3_5 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_3_6 = part2_io_ProcessValid & check ? io_matrix_3_6 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_3_7 = part2_io_ProcessValid & check ? io_matrix_3_7 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_4_0 = part2_io_ProcessValid & check ? io_matrix_4_0 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_4_1 = part2_io_ProcessValid & check ? io_matrix_4_1 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_4_2 = part2_io_ProcessValid & check ? io_matrix_4_2 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_4_3 = part2_io_ProcessValid & check ? io_matrix_4_3 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_4_4 = part2_io_ProcessValid & check ? io_matrix_4_4 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_4_5 = part2_io_ProcessValid & check ? io_matrix_4_5 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_4_6 = part2_io_ProcessValid & check ? io_matrix_4_6 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_4_7 = part2_io_ProcessValid & check ? io_matrix_4_7 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_5_0 = part2_io_ProcessValid & check ? io_matrix_5_0 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_5_1 = part2_io_ProcessValid & check ? io_matrix_5_1 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_5_2 = part2_io_ProcessValid & check ? io_matrix_5_2 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_5_3 = part2_io_ProcessValid & check ? io_matrix_5_3 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_5_4 = part2_io_ProcessValid & check ? io_matrix_5_4 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_5_5 = part2_io_ProcessValid & check ? io_matrix_5_5 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_5_6 = part2_io_ProcessValid & check ? io_matrix_5_6 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_5_7 = part2_io_ProcessValid & check ? io_matrix_5_7 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_6_0 = part2_io_ProcessValid & check ? io_matrix_6_0 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_6_1 = part2_io_ProcessValid & check ? io_matrix_6_1 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_6_2 = part2_io_ProcessValid & check ? io_matrix_6_2 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_6_3 = part2_io_ProcessValid & check ? io_matrix_6_3 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_6_4 = part2_io_ProcessValid & check ? io_matrix_6_4 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_6_5 = part2_io_ProcessValid & check ? io_matrix_6_5 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_6_6 = part2_io_ProcessValid & check ? io_matrix_6_6 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_6_7 = part2_io_ProcessValid & check ? io_matrix_6_7 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_7_0 = part2_io_ProcessValid & check ? io_matrix_7_0 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_7_1 = part2_io_ProcessValid & check ? io_matrix_7_1 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_7_2 = part2_io_ProcessValid & check ? io_matrix_7_2 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_7_3 = part2_io_ProcessValid & check ? io_matrix_7_3 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_7_4 = part2_io_ProcessValid & check ? io_matrix_7_4 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_7_5 = part2_io_ProcessValid & check ? io_matrix_7_5 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_7_6 = part2_io_ProcessValid & check ? io_matrix_7_6 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_mat_7_7 = part2_io_ProcessValid & check ? io_matrix_7_7 : 32'h0; // @[DIstribution.scala 82:42 87:18 97:22]
  assign part3_io_i_valid = part2_io_ProcessValid & check & part2_io_ProcessValid; // @[DIstribution.scala 82:42 85:22 98:26]
  assign part3_io_merge = part2_io_ProcessValid & check & part3_io_merge_REG; // @[DIstribution.scala 82:42 83:20 96:24]
  always @(posedge clock) begin
    if (reset) begin // @[DIstribution.scala 19:20]
      i <= 32'h0; // @[DIstribution.scala 19:20]
    end else if (io_valid) begin // @[DIstribution.scala 27:21]
      if (i < 32'h7 & _io_validIteration_T_1) begin // @[DIstribution.scala 113:69]
        i <= _i_T_1; // @[DIstribution.scala 114:11]
      end
    end
    if (reset) begin // @[DIstribution.scala 20:20]
      j <= 32'h0; // @[DIstribution.scala 20:20]
    end else if (io_valid) begin // @[DIstribution.scala 27:21]
      if (ab) begin // @[DIstribution.scala 119:68]
        j <= _j_T_1; // @[DIstribution.scala 120:11]
      end else if (!(_io_validIteration_T_2)) begin // @[DIstribution.scala 121:75]
        j <= 32'h0; // @[DIstribution.scala 124:11]
      end
    end
    if (reset) begin // @[DIstribution.scala 21:24]
      count <= 32'h0; // @[DIstribution.scala 21:24]
    end else if (io_valid) begin // @[DIstribution.scala 27:21]
      if (_T_2) begin // @[DIstribution.scala 47:38]
        count <= _count_T_1; // @[DIstribution.scala 48:15]
      end
    end
    if (reset) begin // @[DIstribution.scala 22:23]
      Idex_0 <= 32'h0; // @[DIstribution.scala 22:23]
    end else if (io_valid) begin // @[DIstribution.scala 27:21]
      if (_T_2) begin // @[DIstribution.scala 47:38]
        Idex_0 <= _GEN_129;
      end else if (_T_2 & _io_validIteration_T & _io_validIteration_T_1) begin // @[DIstribution.scala 51:106]
        Idex_0 <= _GEN_129;
      end
    end
    if (reset) begin // @[DIstribution.scala 22:23]
      Idex_1 <= 32'h0; // @[DIstribution.scala 22:23]
    end else if (io_valid) begin // @[DIstribution.scala 27:21]
      if (_T_2) begin // @[DIstribution.scala 47:38]
        Idex_1 <= _GEN_130;
      end else if (_T_2 & _io_validIteration_T & _io_validIteration_T_1) begin // @[DIstribution.scala 51:106]
        Idex_1 <= _GEN_130;
      end
    end
    if (reset) begin // @[DIstribution.scala 22:23]
      Idex_2 <= 32'h0; // @[DIstribution.scala 22:23]
    end else if (io_valid) begin // @[DIstribution.scala 27:21]
      if (_T_2) begin // @[DIstribution.scala 47:38]
        Idex_2 <= _GEN_131;
      end else if (_T_2 & _io_validIteration_T & _io_validIteration_T_1) begin // @[DIstribution.scala 51:106]
        Idex_2 <= _GEN_131;
      end
    end
    if (reset) begin // @[DIstribution.scala 22:23]
      Idex_3 <= 32'h0; // @[DIstribution.scala 22:23]
    end else if (io_valid) begin // @[DIstribution.scala 27:21]
      if (_T_2) begin // @[DIstribution.scala 47:38]
        Idex_3 <= _GEN_132;
      end else if (_T_2 & _io_validIteration_T & _io_validIteration_T_1) begin // @[DIstribution.scala 51:106]
        Idex_3 <= _GEN_132;
      end
    end
    if (reset) begin // @[DIstribution.scala 22:23]
      Idex_4 <= 32'h0; // @[DIstribution.scala 22:23]
    end else if (io_valid) begin // @[DIstribution.scala 27:21]
      if (_T_2) begin // @[DIstribution.scala 47:38]
        Idex_4 <= _GEN_133;
      end else if (_T_2 & _io_validIteration_T & _io_validIteration_T_1) begin // @[DIstribution.scala 51:106]
        Idex_4 <= _GEN_133;
      end
    end
    if (reset) begin // @[DIstribution.scala 22:23]
      Idex_5 <= 32'h0; // @[DIstribution.scala 22:23]
    end else if (io_valid) begin // @[DIstribution.scala 27:21]
      if (_T_2) begin // @[DIstribution.scala 47:38]
        Idex_5 <= _GEN_134;
      end else if (_T_2 & _io_validIteration_T & _io_validIteration_T_1) begin // @[DIstribution.scala 51:106]
        Idex_5 <= _GEN_134;
      end
    end
    if (reset) begin // @[DIstribution.scala 22:23]
      Idex_6 <= 32'h0; // @[DIstribution.scala 22:23]
    end else if (io_valid) begin // @[DIstribution.scala 27:21]
      if (_T_2) begin // @[DIstribution.scala 47:38]
        Idex_6 <= _GEN_135;
      end else if (_T_2 & _io_validIteration_T & _io_validIteration_T_1) begin // @[DIstribution.scala 51:106]
        Idex_6 <= _GEN_135;
      end
    end
    if (reset) begin // @[DIstribution.scala 22:23]
      Idex_7 <= 32'h0; // @[DIstribution.scala 22:23]
    end else if (io_valid) begin // @[DIstribution.scala 27:21]
      if (_T_2) begin // @[DIstribution.scala 47:38]
        Idex_7 <= _GEN_136;
      end else if (_T_2 & _io_validIteration_T & _io_validIteration_T_1) begin // @[DIstribution.scala 51:106]
        Idex_7 <= _GEN_136;
      end
    end
    if (reset) begin // @[DIstribution.scala 23:23]
      Jdex_0 <= 32'h0; // @[DIstribution.scala 23:23]
    end else if (io_valid) begin // @[DIstribution.scala 27:21]
      if (_T_2) begin // @[DIstribution.scala 47:38]
        Jdex_0 <= _GEN_137;
      end else if (_T_2 & _io_validIteration_T & _io_validIteration_T_1) begin // @[DIstribution.scala 51:106]
        Jdex_0 <= _GEN_137;
      end
    end
    if (reset) begin // @[DIstribution.scala 23:23]
      Jdex_1 <= 32'h0; // @[DIstribution.scala 23:23]
    end else if (io_valid) begin // @[DIstribution.scala 27:21]
      if (_T_2) begin // @[DIstribution.scala 47:38]
        Jdex_1 <= _GEN_138;
      end else if (_T_2 & _io_validIteration_T & _io_validIteration_T_1) begin // @[DIstribution.scala 51:106]
        Jdex_1 <= _GEN_138;
      end
    end
    if (reset) begin // @[DIstribution.scala 23:23]
      Jdex_2 <= 32'h0; // @[DIstribution.scala 23:23]
    end else if (io_valid) begin // @[DIstribution.scala 27:21]
      if (_T_2) begin // @[DIstribution.scala 47:38]
        Jdex_2 <= _GEN_139;
      end else if (_T_2 & _io_validIteration_T & _io_validIteration_T_1) begin // @[DIstribution.scala 51:106]
        Jdex_2 <= _GEN_139;
      end
    end
    if (reset) begin // @[DIstribution.scala 23:23]
      Jdex_3 <= 32'h0; // @[DIstribution.scala 23:23]
    end else if (io_valid) begin // @[DIstribution.scala 27:21]
      if (_T_2) begin // @[DIstribution.scala 47:38]
        Jdex_3 <= _GEN_140;
      end else if (_T_2 & _io_validIteration_T & _io_validIteration_T_1) begin // @[DIstribution.scala 51:106]
        Jdex_3 <= _GEN_140;
      end
    end
    if (reset) begin // @[DIstribution.scala 23:23]
      Jdex_4 <= 32'h0; // @[DIstribution.scala 23:23]
    end else if (io_valid) begin // @[DIstribution.scala 27:21]
      if (_T_2) begin // @[DIstribution.scala 47:38]
        Jdex_4 <= _GEN_141;
      end else if (_T_2 & _io_validIteration_T & _io_validIteration_T_1) begin // @[DIstribution.scala 51:106]
        Jdex_4 <= _GEN_141;
      end
    end
    if (reset) begin // @[DIstribution.scala 23:23]
      Jdex_5 <= 32'h0; // @[DIstribution.scala 23:23]
    end else if (io_valid) begin // @[DIstribution.scala 27:21]
      if (_T_2) begin // @[DIstribution.scala 47:38]
        Jdex_5 <= _GEN_142;
      end else if (_T_2 & _io_validIteration_T & _io_validIteration_T_1) begin // @[DIstribution.scala 51:106]
        Jdex_5 <= _GEN_142;
      end
    end
    if (reset) begin // @[DIstribution.scala 23:23]
      Jdex_6 <= 32'h0; // @[DIstribution.scala 23:23]
    end else if (io_valid) begin // @[DIstribution.scala 27:21]
      if (_T_2) begin // @[DIstribution.scala 47:38]
        Jdex_6 <= _GEN_143;
      end else if (_T_2 & _io_validIteration_T & _io_validIteration_T_1) begin // @[DIstribution.scala 51:106]
        Jdex_6 <= _GEN_143;
      end
    end
    if (reset) begin // @[DIstribution.scala 23:23]
      Jdex_7 <= 32'h0; // @[DIstribution.scala 23:23]
    end else if (io_valid) begin // @[DIstribution.scala 27:21]
      if (_T_2) begin // @[DIstribution.scala 47:38]
        Jdex_7 <= _GEN_144;
      end else if (_T_2 & _io_validIteration_T & _io_validIteration_T_1) begin // @[DIstribution.scala 51:106]
        Jdex_7 <= _GEN_144;
      end
    end
    if (reset) begin // @[DIstribution.scala 25:30]
      iterationNo <= 32'h0; // @[DIstribution.scala 25:30]
    end else if (io_valid) begin // @[DIstribution.scala 27:21]
      if (_GEN_63 == 32'h1) begin // @[DIstribution.scala 34:35]
        iterationNo <= _iterationNo_T_1; // @[DIstribution.scala 35:19]
      end
    end
    c <= _io_validIteration_T & _io_validIteration_T_1; // @[DIstribution.scala 57:48]
    part3_io_merge_REG <= c; // @[DIstribution.scala 83:30]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  i = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  j = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  count = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  Idex_0 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  Idex_1 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  Idex_2 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  Idex_3 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  Idex_4 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  Idex_5 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  Idex_6 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  Idex_7 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  Jdex_0 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  Jdex_1 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  Jdex_2 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  Jdex_3 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  Jdex_4 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  Jdex_5 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  Jdex_6 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  Jdex_7 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  iterationNo = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  c = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  part3_io_merge_REG = _RAND_21[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PathFinder(
  input         clock,
  input         reset,
  input  [15:0] io_Stationary_matrix_0_0,
  input  [15:0] io_Stationary_matrix_0_1,
  input  [15:0] io_Stationary_matrix_0_2,
  input  [15:0] io_Stationary_matrix_0_3,
  input  [15:0] io_Stationary_matrix_0_4,
  input  [15:0] io_Stationary_matrix_0_5,
  input  [15:0] io_Stationary_matrix_0_6,
  input  [15:0] io_Stationary_matrix_0_7,
  input  [15:0] io_Stationary_matrix_1_0,
  input  [15:0] io_Stationary_matrix_1_1,
  input  [15:0] io_Stationary_matrix_1_2,
  input  [15:0] io_Stationary_matrix_1_3,
  input  [15:0] io_Stationary_matrix_1_4,
  input  [15:0] io_Stationary_matrix_1_5,
  input  [15:0] io_Stationary_matrix_1_6,
  input  [15:0] io_Stationary_matrix_1_7,
  input  [15:0] io_Stationary_matrix_2_0,
  input  [15:0] io_Stationary_matrix_2_1,
  input  [15:0] io_Stationary_matrix_2_2,
  input  [15:0] io_Stationary_matrix_2_3,
  input  [15:0] io_Stationary_matrix_2_4,
  input  [15:0] io_Stationary_matrix_2_5,
  input  [15:0] io_Stationary_matrix_2_6,
  input  [15:0] io_Stationary_matrix_2_7,
  input  [15:0] io_Stationary_matrix_3_0,
  input  [15:0] io_Stationary_matrix_3_1,
  input  [15:0] io_Stationary_matrix_3_2,
  input  [15:0] io_Stationary_matrix_3_3,
  input  [15:0] io_Stationary_matrix_3_4,
  input  [15:0] io_Stationary_matrix_3_5,
  input  [15:0] io_Stationary_matrix_3_6,
  input  [15:0] io_Stationary_matrix_3_7,
  input  [15:0] io_Stationary_matrix_4_0,
  input  [15:0] io_Stationary_matrix_4_1,
  input  [15:0] io_Stationary_matrix_4_2,
  input  [15:0] io_Stationary_matrix_4_3,
  input  [15:0] io_Stationary_matrix_4_4,
  input  [15:0] io_Stationary_matrix_4_5,
  input  [15:0] io_Stationary_matrix_4_6,
  input  [15:0] io_Stationary_matrix_4_7,
  input  [15:0] io_Stationary_matrix_5_0,
  input  [15:0] io_Stationary_matrix_5_1,
  input  [15:0] io_Stationary_matrix_5_2,
  input  [15:0] io_Stationary_matrix_5_3,
  input  [15:0] io_Stationary_matrix_5_4,
  input  [15:0] io_Stationary_matrix_5_5,
  input  [15:0] io_Stationary_matrix_5_6,
  input  [15:0] io_Stationary_matrix_5_7,
  input  [15:0] io_Stationary_matrix_6_0,
  input  [15:0] io_Stationary_matrix_6_1,
  input  [15:0] io_Stationary_matrix_6_2,
  input  [15:0] io_Stationary_matrix_6_3,
  input  [15:0] io_Stationary_matrix_6_4,
  input  [15:0] io_Stationary_matrix_6_5,
  input  [15:0] io_Stationary_matrix_6_6,
  input  [15:0] io_Stationary_matrix_6_7,
  input  [15:0] io_Stationary_matrix_7_0,
  input  [15:0] io_Stationary_matrix_7_1,
  input  [15:0] io_Stationary_matrix_7_2,
  input  [15:0] io_Stationary_matrix_7_3,
  input  [15:0] io_Stationary_matrix_7_4,
  input  [15:0] io_Stationary_matrix_7_5,
  input  [15:0] io_Stationary_matrix_7_6,
  input  [15:0] io_Stationary_matrix_7_7,
  input  [15:0] io_Streaming_matrix_0,
  input  [15:0] io_Streaming_matrix_1,
  input  [15:0] io_Streaming_matrix_2,
  input  [15:0] io_Streaming_matrix_3,
  input  [15:0] io_Streaming_matrix_4,
  input  [15:0] io_Streaming_matrix_5,
  input  [15:0] io_Streaming_matrix_6,
  input  [15:0] io_Streaming_matrix_7,
  output [3:0]  io_i_mux_bus_0,
  output [3:0]  io_i_mux_bus_1,
  output [3:0]  io_i_mux_bus_2,
  output [3:0]  io_i_mux_bus_3,
  output [15:0] io_Source_0,
  output [15:0] io_Source_1,
  output [15:0] io_Source_2,
  output [15:0] io_Source_3,
  output [15:0] io_destination_0,
  output [15:0] io_destination_1,
  output [15:0] io_destination_2,
  output [15:0] io_destination_3,
  output        io_PF_Valid,
  input  [31:0] io_NoDPE,
  input         io_DataValid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  myMuxes_clock; // @[PathFinder.scala 26:23]
  wire  myMuxes_reset; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_0_0; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_0_1; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_0_2; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_0_3; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_0_4; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_0_5; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_0_6; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_0_7; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_1_0; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_1_1; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_1_2; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_1_3; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_1_4; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_1_5; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_1_6; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_1_7; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_2_0; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_2_1; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_2_2; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_2_3; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_2_4; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_2_5; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_2_6; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_2_7; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_3_0; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_3_1; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_3_2; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_3_3; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_3_4; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_3_5; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_3_6; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_3_7; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_4_0; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_4_1; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_4_2; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_4_3; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_4_4; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_4_5; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_4_6; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_4_7; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_5_0; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_5_1; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_5_2; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_5_3; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_5_4; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_5_5; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_5_6; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_5_7; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_6_0; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_6_1; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_6_2; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_6_3; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_6_4; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_6_5; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_6_6; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_6_7; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_7_0; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_7_1; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_7_2; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_7_3; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_7_4; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_7_5; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_7_6; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat1_7_7; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat2_0; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat2_1; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat2_2; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat2_3; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat2_4; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat2_5; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat2_6; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_mat2_7; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_0_0; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_0_1; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_0_2; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_0_3; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_0_4; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_0_5; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_0_6; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_0_7; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_1_0; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_1_1; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_1_2; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_1_3; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_1_4; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_1_5; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_1_6; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_1_7; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_2_0; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_2_1; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_2_2; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_2_3; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_2_4; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_2_5; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_2_6; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_2_7; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_3_0; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_3_1; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_3_2; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_3_3; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_3_4; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_3_5; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_3_6; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_3_7; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_4_0; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_4_1; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_4_2; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_4_3; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_4_4; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_4_5; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_4_6; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_4_7; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_5_0; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_5_1; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_5_2; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_5_3; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_5_4; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_5_5; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_5_6; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_5_7; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_6_0; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_6_1; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_6_2; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_6_3; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_6_4; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_6_5; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_6_6; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_6_7; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_7_0; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_7_1; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_7_2; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_7_3; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_7_4; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_7_5; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_7_6; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix1_7_7; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix2_0; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix2_1; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix2_2; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix2_3; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix2_4; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix2_5; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix2_6; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_counterMatrix2_7; // @[PathFinder.scala 26:23]
  wire [3:0] myMuxes_io_i_mux_bus_0; // @[PathFinder.scala 26:23]
  wire [3:0] myMuxes_io_i_mux_bus_1; // @[PathFinder.scala 26:23]
  wire [3:0] myMuxes_io_i_mux_bus_2; // @[PathFinder.scala 26:23]
  wire [3:0] myMuxes_io_i_mux_bus_3; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_Source_0; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_Source_1; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_Source_2; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_Source_3; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_destination_0; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_destination_1; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_destination_2; // @[PathFinder.scala 26:23]
  wire [15:0] myMuxes_io_destination_3; // @[PathFinder.scala 26:23]
  wire  myMuxes_io_valid; // @[PathFinder.scala 26:23]
  wire  myCounter_clock; // @[PathFinder.scala 32:25]
  wire  myCounter_reset; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_0_0; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_0_1; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_0_2; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_0_3; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_0_4; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_0_5; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_0_6; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_0_7; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_1_0; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_1_1; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_1_2; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_1_3; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_1_4; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_1_5; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_1_6; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_1_7; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_2_0; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_2_1; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_2_2; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_2_3; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_2_4; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_2_5; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_2_6; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_2_7; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_3_0; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_3_1; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_3_2; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_3_3; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_3_4; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_3_5; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_3_6; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_3_7; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_4_0; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_4_1; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_4_2; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_4_3; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_4_4; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_4_5; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_4_6; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_4_7; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_5_0; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_5_1; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_5_2; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_5_3; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_5_4; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_5_5; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_5_6; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_5_7; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_6_0; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_6_1; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_6_2; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_6_3; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_6_4; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_6_5; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_6_6; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_6_7; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_7_0; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_7_1; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_7_2; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_7_3; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_7_4; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_7_5; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_7_6; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Stationary_matrix_7_7; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Streaming_matrix_0; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Streaming_matrix_1; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Streaming_matrix_2; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Streaming_matrix_3; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Streaming_matrix_4; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Streaming_matrix_5; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Streaming_matrix_6; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_Streaming_matrix_7; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_0_0; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_0_1; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_0_2; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_0_3; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_0_4; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_0_5; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_0_6; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_0_7; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_1_0; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_1_1; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_1_2; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_1_3; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_1_4; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_1_5; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_1_6; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_1_7; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_2_0; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_2_1; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_2_2; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_2_3; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_2_4; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_2_5; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_2_6; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_2_7; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_3_0; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_3_1; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_3_2; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_3_3; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_3_4; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_3_5; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_3_6; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_3_7; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_4_0; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_4_1; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_4_2; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_4_3; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_4_4; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_4_5; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_4_6; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_4_7; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_5_0; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_5_1; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_5_2; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_5_3; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_5_4; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_5_5; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_5_6; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_5_7; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_6_0; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_6_1; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_6_2; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_6_3; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_6_4; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_6_5; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_6_6; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_6_7; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_7_0; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_7_1; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_7_2; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_7_3; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_7_4; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_7_5; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_7_6; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_7_7; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix2_bits_0; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix2_bits_1; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix2_bits_2; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix2_bits_3; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix2_bits_4; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix2_bits_5; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix2_bits_6; // @[PathFinder.scala 32:25]
  wire [15:0] myCounter_io_counterMatrix2_bits_7; // @[PathFinder.scala 32:25]
  wire  myCounter_io_valid; // @[PathFinder.scala 32:25]
  wire  myCounter_io_start; // @[PathFinder.scala 32:25]
  wire  Distribution_clock; // @[PathFinder.scala 37:28]
  wire  Distribution_reset; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_0_0; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_0_1; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_0_2; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_0_3; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_0_4; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_0_5; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_0_6; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_0_7; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_1_0; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_1_1; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_1_2; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_1_3; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_1_4; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_1_5; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_1_6; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_1_7; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_2_0; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_2_1; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_2_2; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_2_3; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_2_4; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_2_5; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_2_6; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_2_7; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_3_0; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_3_1; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_3_2; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_3_3; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_3_4; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_3_5; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_3_6; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_3_7; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_4_0; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_4_1; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_4_2; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_4_3; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_4_4; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_4_5; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_4_6; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_4_7; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_5_0; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_5_1; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_5_2; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_5_3; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_5_4; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_5_5; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_5_6; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_5_7; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_6_0; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_6_1; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_6_2; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_6_3; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_6_4; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_6_5; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_6_6; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_6_7; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_7_0; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_7_1; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_7_2; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_7_3; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_7_4; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_7_5; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_7_6; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_matrix_7_7; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_s; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_0_0; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_0_1; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_0_2; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_0_3; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_0_4; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_0_5; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_0_6; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_0_7; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_1_0; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_1_1; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_1_2; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_1_3; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_1_4; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_1_5; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_1_6; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_1_7; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_2_0; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_2_1; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_2_2; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_2_3; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_2_4; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_2_5; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_2_6; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_2_7; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_3_0; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_3_1; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_3_2; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_3_3; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_3_4; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_3_5; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_3_6; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_3_7; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_4_0; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_4_1; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_4_2; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_4_3; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_4_4; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_4_5; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_4_6; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_4_7; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_5_0; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_5_1; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_5_2; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_5_3; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_5_4; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_5_5; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_5_6; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_5_7; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_6_0; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_6_1; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_6_2; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_6_3; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_6_4; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_6_5; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_6_6; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_6_7; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_7_0; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_7_1; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_7_2; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_7_3; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_7_4; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_7_5; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_7_6; // @[PathFinder.scala 37:28]
  wire [31:0] Distribution_io_out_7_7; // @[PathFinder.scala 37:28]
  wire  Distribution_io_ProcessValid; // @[PathFinder.scala 37:28]
  wire  Distribution_io_valid; // @[PathFinder.scala 37:28]
  reg  myCounter_io_start_REG; // @[PathFinder.scala 33:32]
  wire [31:0] _GEN_73 = Distribution_io_ProcessValid ? Distribution_io_out_0_0 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_74 = Distribution_io_ProcessValid ? Distribution_io_out_0_1 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_75 = Distribution_io_ProcessValid ? Distribution_io_out_0_2 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_76 = Distribution_io_ProcessValid ? Distribution_io_out_0_3 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_77 = Distribution_io_ProcessValid ? Distribution_io_out_0_4 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_78 = Distribution_io_ProcessValid ? Distribution_io_out_0_5 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_79 = Distribution_io_ProcessValid ? Distribution_io_out_0_6 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_80 = Distribution_io_ProcessValid ? Distribution_io_out_0_7 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_81 = Distribution_io_ProcessValid ? Distribution_io_out_1_0 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_82 = Distribution_io_ProcessValid ? Distribution_io_out_1_1 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_83 = Distribution_io_ProcessValid ? Distribution_io_out_1_2 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_84 = Distribution_io_ProcessValid ? Distribution_io_out_1_3 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_85 = Distribution_io_ProcessValid ? Distribution_io_out_1_4 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_86 = Distribution_io_ProcessValid ? Distribution_io_out_1_5 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_87 = Distribution_io_ProcessValid ? Distribution_io_out_1_6 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_88 = Distribution_io_ProcessValid ? Distribution_io_out_1_7 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_89 = Distribution_io_ProcessValid ? Distribution_io_out_2_0 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_90 = Distribution_io_ProcessValid ? Distribution_io_out_2_1 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_91 = Distribution_io_ProcessValid ? Distribution_io_out_2_2 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_92 = Distribution_io_ProcessValid ? Distribution_io_out_2_3 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_93 = Distribution_io_ProcessValid ? Distribution_io_out_2_4 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_94 = Distribution_io_ProcessValid ? Distribution_io_out_2_5 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_95 = Distribution_io_ProcessValid ? Distribution_io_out_2_6 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_96 = Distribution_io_ProcessValid ? Distribution_io_out_2_7 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_97 = Distribution_io_ProcessValid ? Distribution_io_out_3_0 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_98 = Distribution_io_ProcessValid ? Distribution_io_out_3_1 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_99 = Distribution_io_ProcessValid ? Distribution_io_out_3_2 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_100 = Distribution_io_ProcessValid ? Distribution_io_out_3_3 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_101 = Distribution_io_ProcessValid ? Distribution_io_out_3_4 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_102 = Distribution_io_ProcessValid ? Distribution_io_out_3_5 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_103 = Distribution_io_ProcessValid ? Distribution_io_out_3_6 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_104 = Distribution_io_ProcessValid ? Distribution_io_out_3_7 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_105 = Distribution_io_ProcessValid ? Distribution_io_out_4_0 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_106 = Distribution_io_ProcessValid ? Distribution_io_out_4_1 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_107 = Distribution_io_ProcessValid ? Distribution_io_out_4_2 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_108 = Distribution_io_ProcessValid ? Distribution_io_out_4_3 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_109 = Distribution_io_ProcessValid ? Distribution_io_out_4_4 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_110 = Distribution_io_ProcessValid ? Distribution_io_out_4_5 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_111 = Distribution_io_ProcessValid ? Distribution_io_out_4_6 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_112 = Distribution_io_ProcessValid ? Distribution_io_out_4_7 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_113 = Distribution_io_ProcessValid ? Distribution_io_out_5_0 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_114 = Distribution_io_ProcessValid ? Distribution_io_out_5_1 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_115 = Distribution_io_ProcessValid ? Distribution_io_out_5_2 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_116 = Distribution_io_ProcessValid ? Distribution_io_out_5_3 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_117 = Distribution_io_ProcessValid ? Distribution_io_out_5_4 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_118 = Distribution_io_ProcessValid ? Distribution_io_out_5_5 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_119 = Distribution_io_ProcessValid ? Distribution_io_out_5_6 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_120 = Distribution_io_ProcessValid ? Distribution_io_out_5_7 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_121 = Distribution_io_ProcessValid ? Distribution_io_out_6_0 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_122 = Distribution_io_ProcessValid ? Distribution_io_out_6_1 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_123 = Distribution_io_ProcessValid ? Distribution_io_out_6_2 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_124 = Distribution_io_ProcessValid ? Distribution_io_out_6_3 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_125 = Distribution_io_ProcessValid ? Distribution_io_out_6_4 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_126 = Distribution_io_ProcessValid ? Distribution_io_out_6_5 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_127 = Distribution_io_ProcessValid ? Distribution_io_out_6_6 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_128 = Distribution_io_ProcessValid ? Distribution_io_out_6_7 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_129 = Distribution_io_ProcessValid ? Distribution_io_out_7_0 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_130 = Distribution_io_ProcessValid ? Distribution_io_out_7_1 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_131 = Distribution_io_ProcessValid ? Distribution_io_out_7_2 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_132 = Distribution_io_ProcessValid ? Distribution_io_out_7_3 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_133 = Distribution_io_ProcessValid ? Distribution_io_out_7_4 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_134 = Distribution_io_ProcessValid ? Distribution_io_out_7_5 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_135 = Distribution_io_ProcessValid ? Distribution_io_out_7_6 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_136 = Distribution_io_ProcessValid ? Distribution_io_out_7_7 : 32'h0; // @[PathFinder.scala 52:40 58:31 67:31]
  wire [31:0] _GEN_148 = io_DataValid ? {{28'd0}, myMuxes_io_i_mux_bus_0} : 32'h0; // @[PathFinder.scala 20:20 75:16 82:16]
  wire [31:0] _GEN_149 = io_DataValid ? {{28'd0}, myMuxes_io_i_mux_bus_1} : 32'h0; // @[PathFinder.scala 20:20 75:16 82:16]
  wire [31:0] _GEN_150 = io_DataValid ? {{28'd0}, myMuxes_io_i_mux_bus_2} : 32'h0; // @[PathFinder.scala 20:20 75:16 82:16]
  wire [31:0] _GEN_151 = io_DataValid ? {{28'd0}, myMuxes_io_i_mux_bus_3} : 32'h0; // @[PathFinder.scala 20:20 75:16 82:16]
  wire [31:0] _GEN_212 = io_DataValid ? {{16'd0}, myMuxes_io_Source_0} : 32'h0; // @[PathFinder.scala 20:20 76:13 83:13]
  wire [31:0] _GEN_213 = io_DataValid ? {{16'd0}, myMuxes_io_Source_1} : 32'h0; // @[PathFinder.scala 20:20 76:13 83:13]
  wire [31:0] _GEN_214 = io_DataValid ? {{16'd0}, myMuxes_io_Source_2} : 32'h0; // @[PathFinder.scala 20:20 76:13 83:13]
  wire [31:0] _GEN_215 = io_DataValid ? {{16'd0}, myMuxes_io_Source_3} : 32'h0; // @[PathFinder.scala 20:20 76:13 83:13]
  wire [31:0] _GEN_276 = io_DataValid ? {{16'd0}, myMuxes_io_destination_0} : 32'h0; // @[PathFinder.scala 20:20 77:18 84:18]
  wire [31:0] _GEN_277 = io_DataValid ? {{16'd0}, myMuxes_io_destination_1} : 32'h0; // @[PathFinder.scala 20:20 77:18 84:18]
  wire [31:0] _GEN_278 = io_DataValid ? {{16'd0}, myMuxes_io_destination_2} : 32'h0; // @[PathFinder.scala 20:20 77:18 84:18]
  wire [31:0] _GEN_279 = io_DataValid ? {{16'd0}, myMuxes_io_destination_3} : 32'h0; // @[PathFinder.scala 20:20 77:18 84:18]
  Muxes myMuxes ( // @[PathFinder.scala 26:23]
    .clock(myMuxes_clock),
    .reset(myMuxes_reset),
    .io_mat1_0_0(myMuxes_io_mat1_0_0),
    .io_mat1_0_1(myMuxes_io_mat1_0_1),
    .io_mat1_0_2(myMuxes_io_mat1_0_2),
    .io_mat1_0_3(myMuxes_io_mat1_0_3),
    .io_mat1_0_4(myMuxes_io_mat1_0_4),
    .io_mat1_0_5(myMuxes_io_mat1_0_5),
    .io_mat1_0_6(myMuxes_io_mat1_0_6),
    .io_mat1_0_7(myMuxes_io_mat1_0_7),
    .io_mat1_1_0(myMuxes_io_mat1_1_0),
    .io_mat1_1_1(myMuxes_io_mat1_1_1),
    .io_mat1_1_2(myMuxes_io_mat1_1_2),
    .io_mat1_1_3(myMuxes_io_mat1_1_3),
    .io_mat1_1_4(myMuxes_io_mat1_1_4),
    .io_mat1_1_5(myMuxes_io_mat1_1_5),
    .io_mat1_1_6(myMuxes_io_mat1_1_6),
    .io_mat1_1_7(myMuxes_io_mat1_1_7),
    .io_mat1_2_0(myMuxes_io_mat1_2_0),
    .io_mat1_2_1(myMuxes_io_mat1_2_1),
    .io_mat1_2_2(myMuxes_io_mat1_2_2),
    .io_mat1_2_3(myMuxes_io_mat1_2_3),
    .io_mat1_2_4(myMuxes_io_mat1_2_4),
    .io_mat1_2_5(myMuxes_io_mat1_2_5),
    .io_mat1_2_6(myMuxes_io_mat1_2_6),
    .io_mat1_2_7(myMuxes_io_mat1_2_7),
    .io_mat1_3_0(myMuxes_io_mat1_3_0),
    .io_mat1_3_1(myMuxes_io_mat1_3_1),
    .io_mat1_3_2(myMuxes_io_mat1_3_2),
    .io_mat1_3_3(myMuxes_io_mat1_3_3),
    .io_mat1_3_4(myMuxes_io_mat1_3_4),
    .io_mat1_3_5(myMuxes_io_mat1_3_5),
    .io_mat1_3_6(myMuxes_io_mat1_3_6),
    .io_mat1_3_7(myMuxes_io_mat1_3_7),
    .io_mat1_4_0(myMuxes_io_mat1_4_0),
    .io_mat1_4_1(myMuxes_io_mat1_4_1),
    .io_mat1_4_2(myMuxes_io_mat1_4_2),
    .io_mat1_4_3(myMuxes_io_mat1_4_3),
    .io_mat1_4_4(myMuxes_io_mat1_4_4),
    .io_mat1_4_5(myMuxes_io_mat1_4_5),
    .io_mat1_4_6(myMuxes_io_mat1_4_6),
    .io_mat1_4_7(myMuxes_io_mat1_4_7),
    .io_mat1_5_0(myMuxes_io_mat1_5_0),
    .io_mat1_5_1(myMuxes_io_mat1_5_1),
    .io_mat1_5_2(myMuxes_io_mat1_5_2),
    .io_mat1_5_3(myMuxes_io_mat1_5_3),
    .io_mat1_5_4(myMuxes_io_mat1_5_4),
    .io_mat1_5_5(myMuxes_io_mat1_5_5),
    .io_mat1_5_6(myMuxes_io_mat1_5_6),
    .io_mat1_5_7(myMuxes_io_mat1_5_7),
    .io_mat1_6_0(myMuxes_io_mat1_6_0),
    .io_mat1_6_1(myMuxes_io_mat1_6_1),
    .io_mat1_6_2(myMuxes_io_mat1_6_2),
    .io_mat1_6_3(myMuxes_io_mat1_6_3),
    .io_mat1_6_4(myMuxes_io_mat1_6_4),
    .io_mat1_6_5(myMuxes_io_mat1_6_5),
    .io_mat1_6_6(myMuxes_io_mat1_6_6),
    .io_mat1_6_7(myMuxes_io_mat1_6_7),
    .io_mat1_7_0(myMuxes_io_mat1_7_0),
    .io_mat1_7_1(myMuxes_io_mat1_7_1),
    .io_mat1_7_2(myMuxes_io_mat1_7_2),
    .io_mat1_7_3(myMuxes_io_mat1_7_3),
    .io_mat1_7_4(myMuxes_io_mat1_7_4),
    .io_mat1_7_5(myMuxes_io_mat1_7_5),
    .io_mat1_7_6(myMuxes_io_mat1_7_6),
    .io_mat1_7_7(myMuxes_io_mat1_7_7),
    .io_mat2_0(myMuxes_io_mat2_0),
    .io_mat2_1(myMuxes_io_mat2_1),
    .io_mat2_2(myMuxes_io_mat2_2),
    .io_mat2_3(myMuxes_io_mat2_3),
    .io_mat2_4(myMuxes_io_mat2_4),
    .io_mat2_5(myMuxes_io_mat2_5),
    .io_mat2_6(myMuxes_io_mat2_6),
    .io_mat2_7(myMuxes_io_mat2_7),
    .io_counterMatrix1_0_0(myMuxes_io_counterMatrix1_0_0),
    .io_counterMatrix1_0_1(myMuxes_io_counterMatrix1_0_1),
    .io_counterMatrix1_0_2(myMuxes_io_counterMatrix1_0_2),
    .io_counterMatrix1_0_3(myMuxes_io_counterMatrix1_0_3),
    .io_counterMatrix1_0_4(myMuxes_io_counterMatrix1_0_4),
    .io_counterMatrix1_0_5(myMuxes_io_counterMatrix1_0_5),
    .io_counterMatrix1_0_6(myMuxes_io_counterMatrix1_0_6),
    .io_counterMatrix1_0_7(myMuxes_io_counterMatrix1_0_7),
    .io_counterMatrix1_1_0(myMuxes_io_counterMatrix1_1_0),
    .io_counterMatrix1_1_1(myMuxes_io_counterMatrix1_1_1),
    .io_counterMatrix1_1_2(myMuxes_io_counterMatrix1_1_2),
    .io_counterMatrix1_1_3(myMuxes_io_counterMatrix1_1_3),
    .io_counterMatrix1_1_4(myMuxes_io_counterMatrix1_1_4),
    .io_counterMatrix1_1_5(myMuxes_io_counterMatrix1_1_5),
    .io_counterMatrix1_1_6(myMuxes_io_counterMatrix1_1_6),
    .io_counterMatrix1_1_7(myMuxes_io_counterMatrix1_1_7),
    .io_counterMatrix1_2_0(myMuxes_io_counterMatrix1_2_0),
    .io_counterMatrix1_2_1(myMuxes_io_counterMatrix1_2_1),
    .io_counterMatrix1_2_2(myMuxes_io_counterMatrix1_2_2),
    .io_counterMatrix1_2_3(myMuxes_io_counterMatrix1_2_3),
    .io_counterMatrix1_2_4(myMuxes_io_counterMatrix1_2_4),
    .io_counterMatrix1_2_5(myMuxes_io_counterMatrix1_2_5),
    .io_counterMatrix1_2_6(myMuxes_io_counterMatrix1_2_6),
    .io_counterMatrix1_2_7(myMuxes_io_counterMatrix1_2_7),
    .io_counterMatrix1_3_0(myMuxes_io_counterMatrix1_3_0),
    .io_counterMatrix1_3_1(myMuxes_io_counterMatrix1_3_1),
    .io_counterMatrix1_3_2(myMuxes_io_counterMatrix1_3_2),
    .io_counterMatrix1_3_3(myMuxes_io_counterMatrix1_3_3),
    .io_counterMatrix1_3_4(myMuxes_io_counterMatrix1_3_4),
    .io_counterMatrix1_3_5(myMuxes_io_counterMatrix1_3_5),
    .io_counterMatrix1_3_6(myMuxes_io_counterMatrix1_3_6),
    .io_counterMatrix1_3_7(myMuxes_io_counterMatrix1_3_7),
    .io_counterMatrix1_4_0(myMuxes_io_counterMatrix1_4_0),
    .io_counterMatrix1_4_1(myMuxes_io_counterMatrix1_4_1),
    .io_counterMatrix1_4_2(myMuxes_io_counterMatrix1_4_2),
    .io_counterMatrix1_4_3(myMuxes_io_counterMatrix1_4_3),
    .io_counterMatrix1_4_4(myMuxes_io_counterMatrix1_4_4),
    .io_counterMatrix1_4_5(myMuxes_io_counterMatrix1_4_5),
    .io_counterMatrix1_4_6(myMuxes_io_counterMatrix1_4_6),
    .io_counterMatrix1_4_7(myMuxes_io_counterMatrix1_4_7),
    .io_counterMatrix1_5_0(myMuxes_io_counterMatrix1_5_0),
    .io_counterMatrix1_5_1(myMuxes_io_counterMatrix1_5_1),
    .io_counterMatrix1_5_2(myMuxes_io_counterMatrix1_5_2),
    .io_counterMatrix1_5_3(myMuxes_io_counterMatrix1_5_3),
    .io_counterMatrix1_5_4(myMuxes_io_counterMatrix1_5_4),
    .io_counterMatrix1_5_5(myMuxes_io_counterMatrix1_5_5),
    .io_counterMatrix1_5_6(myMuxes_io_counterMatrix1_5_6),
    .io_counterMatrix1_5_7(myMuxes_io_counterMatrix1_5_7),
    .io_counterMatrix1_6_0(myMuxes_io_counterMatrix1_6_0),
    .io_counterMatrix1_6_1(myMuxes_io_counterMatrix1_6_1),
    .io_counterMatrix1_6_2(myMuxes_io_counterMatrix1_6_2),
    .io_counterMatrix1_6_3(myMuxes_io_counterMatrix1_6_3),
    .io_counterMatrix1_6_4(myMuxes_io_counterMatrix1_6_4),
    .io_counterMatrix1_6_5(myMuxes_io_counterMatrix1_6_5),
    .io_counterMatrix1_6_6(myMuxes_io_counterMatrix1_6_6),
    .io_counterMatrix1_6_7(myMuxes_io_counterMatrix1_6_7),
    .io_counterMatrix1_7_0(myMuxes_io_counterMatrix1_7_0),
    .io_counterMatrix1_7_1(myMuxes_io_counterMatrix1_7_1),
    .io_counterMatrix1_7_2(myMuxes_io_counterMatrix1_7_2),
    .io_counterMatrix1_7_3(myMuxes_io_counterMatrix1_7_3),
    .io_counterMatrix1_7_4(myMuxes_io_counterMatrix1_7_4),
    .io_counterMatrix1_7_5(myMuxes_io_counterMatrix1_7_5),
    .io_counterMatrix1_7_6(myMuxes_io_counterMatrix1_7_6),
    .io_counterMatrix1_7_7(myMuxes_io_counterMatrix1_7_7),
    .io_counterMatrix2_0(myMuxes_io_counterMatrix2_0),
    .io_counterMatrix2_1(myMuxes_io_counterMatrix2_1),
    .io_counterMatrix2_2(myMuxes_io_counterMatrix2_2),
    .io_counterMatrix2_3(myMuxes_io_counterMatrix2_3),
    .io_counterMatrix2_4(myMuxes_io_counterMatrix2_4),
    .io_counterMatrix2_5(myMuxes_io_counterMatrix2_5),
    .io_counterMatrix2_6(myMuxes_io_counterMatrix2_6),
    .io_counterMatrix2_7(myMuxes_io_counterMatrix2_7),
    .io_i_mux_bus_0(myMuxes_io_i_mux_bus_0),
    .io_i_mux_bus_1(myMuxes_io_i_mux_bus_1),
    .io_i_mux_bus_2(myMuxes_io_i_mux_bus_2),
    .io_i_mux_bus_3(myMuxes_io_i_mux_bus_3),
    .io_Source_0(myMuxes_io_Source_0),
    .io_Source_1(myMuxes_io_Source_1),
    .io_Source_2(myMuxes_io_Source_2),
    .io_Source_3(myMuxes_io_Source_3),
    .io_destination_0(myMuxes_io_destination_0),
    .io_destination_1(myMuxes_io_destination_1),
    .io_destination_2(myMuxes_io_destination_2),
    .io_destination_3(myMuxes_io_destination_3),
    .io_valid(myMuxes_io_valid)
  );
  SourceDestination myCounter ( // @[PathFinder.scala 32:25]
    .clock(myCounter_clock),
    .reset(myCounter_reset),
    .io_Stationary_matrix_0_0(myCounter_io_Stationary_matrix_0_0),
    .io_Stationary_matrix_0_1(myCounter_io_Stationary_matrix_0_1),
    .io_Stationary_matrix_0_2(myCounter_io_Stationary_matrix_0_2),
    .io_Stationary_matrix_0_3(myCounter_io_Stationary_matrix_0_3),
    .io_Stationary_matrix_0_4(myCounter_io_Stationary_matrix_0_4),
    .io_Stationary_matrix_0_5(myCounter_io_Stationary_matrix_0_5),
    .io_Stationary_matrix_0_6(myCounter_io_Stationary_matrix_0_6),
    .io_Stationary_matrix_0_7(myCounter_io_Stationary_matrix_0_7),
    .io_Stationary_matrix_1_0(myCounter_io_Stationary_matrix_1_0),
    .io_Stationary_matrix_1_1(myCounter_io_Stationary_matrix_1_1),
    .io_Stationary_matrix_1_2(myCounter_io_Stationary_matrix_1_2),
    .io_Stationary_matrix_1_3(myCounter_io_Stationary_matrix_1_3),
    .io_Stationary_matrix_1_4(myCounter_io_Stationary_matrix_1_4),
    .io_Stationary_matrix_1_5(myCounter_io_Stationary_matrix_1_5),
    .io_Stationary_matrix_1_6(myCounter_io_Stationary_matrix_1_6),
    .io_Stationary_matrix_1_7(myCounter_io_Stationary_matrix_1_7),
    .io_Stationary_matrix_2_0(myCounter_io_Stationary_matrix_2_0),
    .io_Stationary_matrix_2_1(myCounter_io_Stationary_matrix_2_1),
    .io_Stationary_matrix_2_2(myCounter_io_Stationary_matrix_2_2),
    .io_Stationary_matrix_2_3(myCounter_io_Stationary_matrix_2_3),
    .io_Stationary_matrix_2_4(myCounter_io_Stationary_matrix_2_4),
    .io_Stationary_matrix_2_5(myCounter_io_Stationary_matrix_2_5),
    .io_Stationary_matrix_2_6(myCounter_io_Stationary_matrix_2_6),
    .io_Stationary_matrix_2_7(myCounter_io_Stationary_matrix_2_7),
    .io_Stationary_matrix_3_0(myCounter_io_Stationary_matrix_3_0),
    .io_Stationary_matrix_3_1(myCounter_io_Stationary_matrix_3_1),
    .io_Stationary_matrix_3_2(myCounter_io_Stationary_matrix_3_2),
    .io_Stationary_matrix_3_3(myCounter_io_Stationary_matrix_3_3),
    .io_Stationary_matrix_3_4(myCounter_io_Stationary_matrix_3_4),
    .io_Stationary_matrix_3_5(myCounter_io_Stationary_matrix_3_5),
    .io_Stationary_matrix_3_6(myCounter_io_Stationary_matrix_3_6),
    .io_Stationary_matrix_3_7(myCounter_io_Stationary_matrix_3_7),
    .io_Stationary_matrix_4_0(myCounter_io_Stationary_matrix_4_0),
    .io_Stationary_matrix_4_1(myCounter_io_Stationary_matrix_4_1),
    .io_Stationary_matrix_4_2(myCounter_io_Stationary_matrix_4_2),
    .io_Stationary_matrix_4_3(myCounter_io_Stationary_matrix_4_3),
    .io_Stationary_matrix_4_4(myCounter_io_Stationary_matrix_4_4),
    .io_Stationary_matrix_4_5(myCounter_io_Stationary_matrix_4_5),
    .io_Stationary_matrix_4_6(myCounter_io_Stationary_matrix_4_6),
    .io_Stationary_matrix_4_7(myCounter_io_Stationary_matrix_4_7),
    .io_Stationary_matrix_5_0(myCounter_io_Stationary_matrix_5_0),
    .io_Stationary_matrix_5_1(myCounter_io_Stationary_matrix_5_1),
    .io_Stationary_matrix_5_2(myCounter_io_Stationary_matrix_5_2),
    .io_Stationary_matrix_5_3(myCounter_io_Stationary_matrix_5_3),
    .io_Stationary_matrix_5_4(myCounter_io_Stationary_matrix_5_4),
    .io_Stationary_matrix_5_5(myCounter_io_Stationary_matrix_5_5),
    .io_Stationary_matrix_5_6(myCounter_io_Stationary_matrix_5_6),
    .io_Stationary_matrix_5_7(myCounter_io_Stationary_matrix_5_7),
    .io_Stationary_matrix_6_0(myCounter_io_Stationary_matrix_6_0),
    .io_Stationary_matrix_6_1(myCounter_io_Stationary_matrix_6_1),
    .io_Stationary_matrix_6_2(myCounter_io_Stationary_matrix_6_2),
    .io_Stationary_matrix_6_3(myCounter_io_Stationary_matrix_6_3),
    .io_Stationary_matrix_6_4(myCounter_io_Stationary_matrix_6_4),
    .io_Stationary_matrix_6_5(myCounter_io_Stationary_matrix_6_5),
    .io_Stationary_matrix_6_6(myCounter_io_Stationary_matrix_6_6),
    .io_Stationary_matrix_6_7(myCounter_io_Stationary_matrix_6_7),
    .io_Stationary_matrix_7_0(myCounter_io_Stationary_matrix_7_0),
    .io_Stationary_matrix_7_1(myCounter_io_Stationary_matrix_7_1),
    .io_Stationary_matrix_7_2(myCounter_io_Stationary_matrix_7_2),
    .io_Stationary_matrix_7_3(myCounter_io_Stationary_matrix_7_3),
    .io_Stationary_matrix_7_4(myCounter_io_Stationary_matrix_7_4),
    .io_Stationary_matrix_7_5(myCounter_io_Stationary_matrix_7_5),
    .io_Stationary_matrix_7_6(myCounter_io_Stationary_matrix_7_6),
    .io_Stationary_matrix_7_7(myCounter_io_Stationary_matrix_7_7),
    .io_Streaming_matrix_0(myCounter_io_Streaming_matrix_0),
    .io_Streaming_matrix_1(myCounter_io_Streaming_matrix_1),
    .io_Streaming_matrix_2(myCounter_io_Streaming_matrix_2),
    .io_Streaming_matrix_3(myCounter_io_Streaming_matrix_3),
    .io_Streaming_matrix_4(myCounter_io_Streaming_matrix_4),
    .io_Streaming_matrix_5(myCounter_io_Streaming_matrix_5),
    .io_Streaming_matrix_6(myCounter_io_Streaming_matrix_6),
    .io_Streaming_matrix_7(myCounter_io_Streaming_matrix_7),
    .io_counterMatrix1_bits_0_0(myCounter_io_counterMatrix1_bits_0_0),
    .io_counterMatrix1_bits_0_1(myCounter_io_counterMatrix1_bits_0_1),
    .io_counterMatrix1_bits_0_2(myCounter_io_counterMatrix1_bits_0_2),
    .io_counterMatrix1_bits_0_3(myCounter_io_counterMatrix1_bits_0_3),
    .io_counterMatrix1_bits_0_4(myCounter_io_counterMatrix1_bits_0_4),
    .io_counterMatrix1_bits_0_5(myCounter_io_counterMatrix1_bits_0_5),
    .io_counterMatrix1_bits_0_6(myCounter_io_counterMatrix1_bits_0_6),
    .io_counterMatrix1_bits_0_7(myCounter_io_counterMatrix1_bits_0_7),
    .io_counterMatrix1_bits_1_0(myCounter_io_counterMatrix1_bits_1_0),
    .io_counterMatrix1_bits_1_1(myCounter_io_counterMatrix1_bits_1_1),
    .io_counterMatrix1_bits_1_2(myCounter_io_counterMatrix1_bits_1_2),
    .io_counterMatrix1_bits_1_3(myCounter_io_counterMatrix1_bits_1_3),
    .io_counterMatrix1_bits_1_4(myCounter_io_counterMatrix1_bits_1_4),
    .io_counterMatrix1_bits_1_5(myCounter_io_counterMatrix1_bits_1_5),
    .io_counterMatrix1_bits_1_6(myCounter_io_counterMatrix1_bits_1_6),
    .io_counterMatrix1_bits_1_7(myCounter_io_counterMatrix1_bits_1_7),
    .io_counterMatrix1_bits_2_0(myCounter_io_counterMatrix1_bits_2_0),
    .io_counterMatrix1_bits_2_1(myCounter_io_counterMatrix1_bits_2_1),
    .io_counterMatrix1_bits_2_2(myCounter_io_counterMatrix1_bits_2_2),
    .io_counterMatrix1_bits_2_3(myCounter_io_counterMatrix1_bits_2_3),
    .io_counterMatrix1_bits_2_4(myCounter_io_counterMatrix1_bits_2_4),
    .io_counterMatrix1_bits_2_5(myCounter_io_counterMatrix1_bits_2_5),
    .io_counterMatrix1_bits_2_6(myCounter_io_counterMatrix1_bits_2_6),
    .io_counterMatrix1_bits_2_7(myCounter_io_counterMatrix1_bits_2_7),
    .io_counterMatrix1_bits_3_0(myCounter_io_counterMatrix1_bits_3_0),
    .io_counterMatrix1_bits_3_1(myCounter_io_counterMatrix1_bits_3_1),
    .io_counterMatrix1_bits_3_2(myCounter_io_counterMatrix1_bits_3_2),
    .io_counterMatrix1_bits_3_3(myCounter_io_counterMatrix1_bits_3_3),
    .io_counterMatrix1_bits_3_4(myCounter_io_counterMatrix1_bits_3_4),
    .io_counterMatrix1_bits_3_5(myCounter_io_counterMatrix1_bits_3_5),
    .io_counterMatrix1_bits_3_6(myCounter_io_counterMatrix1_bits_3_6),
    .io_counterMatrix1_bits_3_7(myCounter_io_counterMatrix1_bits_3_7),
    .io_counterMatrix1_bits_4_0(myCounter_io_counterMatrix1_bits_4_0),
    .io_counterMatrix1_bits_4_1(myCounter_io_counterMatrix1_bits_4_1),
    .io_counterMatrix1_bits_4_2(myCounter_io_counterMatrix1_bits_4_2),
    .io_counterMatrix1_bits_4_3(myCounter_io_counterMatrix1_bits_4_3),
    .io_counterMatrix1_bits_4_4(myCounter_io_counterMatrix1_bits_4_4),
    .io_counterMatrix1_bits_4_5(myCounter_io_counterMatrix1_bits_4_5),
    .io_counterMatrix1_bits_4_6(myCounter_io_counterMatrix1_bits_4_6),
    .io_counterMatrix1_bits_4_7(myCounter_io_counterMatrix1_bits_4_7),
    .io_counterMatrix1_bits_5_0(myCounter_io_counterMatrix1_bits_5_0),
    .io_counterMatrix1_bits_5_1(myCounter_io_counterMatrix1_bits_5_1),
    .io_counterMatrix1_bits_5_2(myCounter_io_counterMatrix1_bits_5_2),
    .io_counterMatrix1_bits_5_3(myCounter_io_counterMatrix1_bits_5_3),
    .io_counterMatrix1_bits_5_4(myCounter_io_counterMatrix1_bits_5_4),
    .io_counterMatrix1_bits_5_5(myCounter_io_counterMatrix1_bits_5_5),
    .io_counterMatrix1_bits_5_6(myCounter_io_counterMatrix1_bits_5_6),
    .io_counterMatrix1_bits_5_7(myCounter_io_counterMatrix1_bits_5_7),
    .io_counterMatrix1_bits_6_0(myCounter_io_counterMatrix1_bits_6_0),
    .io_counterMatrix1_bits_6_1(myCounter_io_counterMatrix1_bits_6_1),
    .io_counterMatrix1_bits_6_2(myCounter_io_counterMatrix1_bits_6_2),
    .io_counterMatrix1_bits_6_3(myCounter_io_counterMatrix1_bits_6_3),
    .io_counterMatrix1_bits_6_4(myCounter_io_counterMatrix1_bits_6_4),
    .io_counterMatrix1_bits_6_5(myCounter_io_counterMatrix1_bits_6_5),
    .io_counterMatrix1_bits_6_6(myCounter_io_counterMatrix1_bits_6_6),
    .io_counterMatrix1_bits_6_7(myCounter_io_counterMatrix1_bits_6_7),
    .io_counterMatrix1_bits_7_0(myCounter_io_counterMatrix1_bits_7_0),
    .io_counterMatrix1_bits_7_1(myCounter_io_counterMatrix1_bits_7_1),
    .io_counterMatrix1_bits_7_2(myCounter_io_counterMatrix1_bits_7_2),
    .io_counterMatrix1_bits_7_3(myCounter_io_counterMatrix1_bits_7_3),
    .io_counterMatrix1_bits_7_4(myCounter_io_counterMatrix1_bits_7_4),
    .io_counterMatrix1_bits_7_5(myCounter_io_counterMatrix1_bits_7_5),
    .io_counterMatrix1_bits_7_6(myCounter_io_counterMatrix1_bits_7_6),
    .io_counterMatrix1_bits_7_7(myCounter_io_counterMatrix1_bits_7_7),
    .io_counterMatrix2_bits_0(myCounter_io_counterMatrix2_bits_0),
    .io_counterMatrix2_bits_1(myCounter_io_counterMatrix2_bits_1),
    .io_counterMatrix2_bits_2(myCounter_io_counterMatrix2_bits_2),
    .io_counterMatrix2_bits_3(myCounter_io_counterMatrix2_bits_3),
    .io_counterMatrix2_bits_4(myCounter_io_counterMatrix2_bits_4),
    .io_counterMatrix2_bits_5(myCounter_io_counterMatrix2_bits_5),
    .io_counterMatrix2_bits_6(myCounter_io_counterMatrix2_bits_6),
    .io_counterMatrix2_bits_7(myCounter_io_counterMatrix2_bits_7),
    .io_valid(myCounter_io_valid),
    .io_start(myCounter_io_start)
  );
  Distribution Distribution ( // @[PathFinder.scala 37:28]
    .clock(Distribution_clock),
    .reset(Distribution_reset),
    .io_matrix_0_0(Distribution_io_matrix_0_0),
    .io_matrix_0_1(Distribution_io_matrix_0_1),
    .io_matrix_0_2(Distribution_io_matrix_0_2),
    .io_matrix_0_3(Distribution_io_matrix_0_3),
    .io_matrix_0_4(Distribution_io_matrix_0_4),
    .io_matrix_0_5(Distribution_io_matrix_0_5),
    .io_matrix_0_6(Distribution_io_matrix_0_6),
    .io_matrix_0_7(Distribution_io_matrix_0_7),
    .io_matrix_1_0(Distribution_io_matrix_1_0),
    .io_matrix_1_1(Distribution_io_matrix_1_1),
    .io_matrix_1_2(Distribution_io_matrix_1_2),
    .io_matrix_1_3(Distribution_io_matrix_1_3),
    .io_matrix_1_4(Distribution_io_matrix_1_4),
    .io_matrix_1_5(Distribution_io_matrix_1_5),
    .io_matrix_1_6(Distribution_io_matrix_1_6),
    .io_matrix_1_7(Distribution_io_matrix_1_7),
    .io_matrix_2_0(Distribution_io_matrix_2_0),
    .io_matrix_2_1(Distribution_io_matrix_2_1),
    .io_matrix_2_2(Distribution_io_matrix_2_2),
    .io_matrix_2_3(Distribution_io_matrix_2_3),
    .io_matrix_2_4(Distribution_io_matrix_2_4),
    .io_matrix_2_5(Distribution_io_matrix_2_5),
    .io_matrix_2_6(Distribution_io_matrix_2_6),
    .io_matrix_2_7(Distribution_io_matrix_2_7),
    .io_matrix_3_0(Distribution_io_matrix_3_0),
    .io_matrix_3_1(Distribution_io_matrix_3_1),
    .io_matrix_3_2(Distribution_io_matrix_3_2),
    .io_matrix_3_3(Distribution_io_matrix_3_3),
    .io_matrix_3_4(Distribution_io_matrix_3_4),
    .io_matrix_3_5(Distribution_io_matrix_3_5),
    .io_matrix_3_6(Distribution_io_matrix_3_6),
    .io_matrix_3_7(Distribution_io_matrix_3_7),
    .io_matrix_4_0(Distribution_io_matrix_4_0),
    .io_matrix_4_1(Distribution_io_matrix_4_1),
    .io_matrix_4_2(Distribution_io_matrix_4_2),
    .io_matrix_4_3(Distribution_io_matrix_4_3),
    .io_matrix_4_4(Distribution_io_matrix_4_4),
    .io_matrix_4_5(Distribution_io_matrix_4_5),
    .io_matrix_4_6(Distribution_io_matrix_4_6),
    .io_matrix_4_7(Distribution_io_matrix_4_7),
    .io_matrix_5_0(Distribution_io_matrix_5_0),
    .io_matrix_5_1(Distribution_io_matrix_5_1),
    .io_matrix_5_2(Distribution_io_matrix_5_2),
    .io_matrix_5_3(Distribution_io_matrix_5_3),
    .io_matrix_5_4(Distribution_io_matrix_5_4),
    .io_matrix_5_5(Distribution_io_matrix_5_5),
    .io_matrix_5_6(Distribution_io_matrix_5_6),
    .io_matrix_5_7(Distribution_io_matrix_5_7),
    .io_matrix_6_0(Distribution_io_matrix_6_0),
    .io_matrix_6_1(Distribution_io_matrix_6_1),
    .io_matrix_6_2(Distribution_io_matrix_6_2),
    .io_matrix_6_3(Distribution_io_matrix_6_3),
    .io_matrix_6_4(Distribution_io_matrix_6_4),
    .io_matrix_6_5(Distribution_io_matrix_6_5),
    .io_matrix_6_6(Distribution_io_matrix_6_6),
    .io_matrix_6_7(Distribution_io_matrix_6_7),
    .io_matrix_7_0(Distribution_io_matrix_7_0),
    .io_matrix_7_1(Distribution_io_matrix_7_1),
    .io_matrix_7_2(Distribution_io_matrix_7_2),
    .io_matrix_7_3(Distribution_io_matrix_7_3),
    .io_matrix_7_4(Distribution_io_matrix_7_4),
    .io_matrix_7_5(Distribution_io_matrix_7_5),
    .io_matrix_7_6(Distribution_io_matrix_7_6),
    .io_matrix_7_7(Distribution_io_matrix_7_7),
    .io_s(Distribution_io_s),
    .io_out_0_0(Distribution_io_out_0_0),
    .io_out_0_1(Distribution_io_out_0_1),
    .io_out_0_2(Distribution_io_out_0_2),
    .io_out_0_3(Distribution_io_out_0_3),
    .io_out_0_4(Distribution_io_out_0_4),
    .io_out_0_5(Distribution_io_out_0_5),
    .io_out_0_6(Distribution_io_out_0_6),
    .io_out_0_7(Distribution_io_out_0_7),
    .io_out_1_0(Distribution_io_out_1_0),
    .io_out_1_1(Distribution_io_out_1_1),
    .io_out_1_2(Distribution_io_out_1_2),
    .io_out_1_3(Distribution_io_out_1_3),
    .io_out_1_4(Distribution_io_out_1_4),
    .io_out_1_5(Distribution_io_out_1_5),
    .io_out_1_6(Distribution_io_out_1_6),
    .io_out_1_7(Distribution_io_out_1_7),
    .io_out_2_0(Distribution_io_out_2_0),
    .io_out_2_1(Distribution_io_out_2_1),
    .io_out_2_2(Distribution_io_out_2_2),
    .io_out_2_3(Distribution_io_out_2_3),
    .io_out_2_4(Distribution_io_out_2_4),
    .io_out_2_5(Distribution_io_out_2_5),
    .io_out_2_6(Distribution_io_out_2_6),
    .io_out_2_7(Distribution_io_out_2_7),
    .io_out_3_0(Distribution_io_out_3_0),
    .io_out_3_1(Distribution_io_out_3_1),
    .io_out_3_2(Distribution_io_out_3_2),
    .io_out_3_3(Distribution_io_out_3_3),
    .io_out_3_4(Distribution_io_out_3_4),
    .io_out_3_5(Distribution_io_out_3_5),
    .io_out_3_6(Distribution_io_out_3_6),
    .io_out_3_7(Distribution_io_out_3_7),
    .io_out_4_0(Distribution_io_out_4_0),
    .io_out_4_1(Distribution_io_out_4_1),
    .io_out_4_2(Distribution_io_out_4_2),
    .io_out_4_3(Distribution_io_out_4_3),
    .io_out_4_4(Distribution_io_out_4_4),
    .io_out_4_5(Distribution_io_out_4_5),
    .io_out_4_6(Distribution_io_out_4_6),
    .io_out_4_7(Distribution_io_out_4_7),
    .io_out_5_0(Distribution_io_out_5_0),
    .io_out_5_1(Distribution_io_out_5_1),
    .io_out_5_2(Distribution_io_out_5_2),
    .io_out_5_3(Distribution_io_out_5_3),
    .io_out_5_4(Distribution_io_out_5_4),
    .io_out_5_5(Distribution_io_out_5_5),
    .io_out_5_6(Distribution_io_out_5_6),
    .io_out_5_7(Distribution_io_out_5_7),
    .io_out_6_0(Distribution_io_out_6_0),
    .io_out_6_1(Distribution_io_out_6_1),
    .io_out_6_2(Distribution_io_out_6_2),
    .io_out_6_3(Distribution_io_out_6_3),
    .io_out_6_4(Distribution_io_out_6_4),
    .io_out_6_5(Distribution_io_out_6_5),
    .io_out_6_6(Distribution_io_out_6_6),
    .io_out_6_7(Distribution_io_out_6_7),
    .io_out_7_0(Distribution_io_out_7_0),
    .io_out_7_1(Distribution_io_out_7_1),
    .io_out_7_2(Distribution_io_out_7_2),
    .io_out_7_3(Distribution_io_out_7_3),
    .io_out_7_4(Distribution_io_out_7_4),
    .io_out_7_5(Distribution_io_out_7_5),
    .io_out_7_6(Distribution_io_out_7_6),
    .io_out_7_7(Distribution_io_out_7_7),
    .io_ProcessValid(Distribution_io_ProcessValid),
    .io_valid(Distribution_io_valid)
  );
  assign io_i_mux_bus_0 = _GEN_148[3:0];
  assign io_i_mux_bus_1 = _GEN_149[3:0];
  assign io_i_mux_bus_2 = _GEN_150[3:0];
  assign io_i_mux_bus_3 = _GEN_151[3:0];
  assign io_Source_0 = _GEN_212[15:0];
  assign io_Source_1 = _GEN_213[15:0];
  assign io_Source_2 = _GEN_214[15:0];
  assign io_Source_3 = _GEN_215[15:0];
  assign io_destination_0 = _GEN_276[15:0];
  assign io_destination_1 = _GEN_277[15:0];
  assign io_destination_2 = _GEN_278[15:0];
  assign io_destination_3 = _GEN_279[15:0];
  assign io_PF_Valid = io_DataValid & myMuxes_io_valid; // @[PathFinder.scala 20:20 74:15 81:15]
  assign myMuxes_clock = clock;
  assign myMuxes_reset = reset;
  assign myMuxes_io_mat1_0_0 = Distribution_io_ProcessValid ? io_Stationary_matrix_0_0 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_0_1 = Distribution_io_ProcessValid ? io_Stationary_matrix_0_1 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_0_2 = Distribution_io_ProcessValid ? io_Stationary_matrix_0_2 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_0_3 = Distribution_io_ProcessValid ? io_Stationary_matrix_0_3 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_0_4 = Distribution_io_ProcessValid ? io_Stationary_matrix_0_4 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_0_5 = Distribution_io_ProcessValid ? io_Stationary_matrix_0_5 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_0_6 = Distribution_io_ProcessValid ? io_Stationary_matrix_0_6 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_0_7 = Distribution_io_ProcessValid ? io_Stationary_matrix_0_7 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_1_0 = Distribution_io_ProcessValid ? io_Stationary_matrix_1_0 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_1_1 = Distribution_io_ProcessValid ? io_Stationary_matrix_1_1 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_1_2 = Distribution_io_ProcessValid ? io_Stationary_matrix_1_2 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_1_3 = Distribution_io_ProcessValid ? io_Stationary_matrix_1_3 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_1_4 = Distribution_io_ProcessValid ? io_Stationary_matrix_1_4 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_1_5 = Distribution_io_ProcessValid ? io_Stationary_matrix_1_5 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_1_6 = Distribution_io_ProcessValid ? io_Stationary_matrix_1_6 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_1_7 = Distribution_io_ProcessValid ? io_Stationary_matrix_1_7 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_2_0 = Distribution_io_ProcessValid ? io_Stationary_matrix_2_0 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_2_1 = Distribution_io_ProcessValid ? io_Stationary_matrix_2_1 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_2_2 = Distribution_io_ProcessValid ? io_Stationary_matrix_2_2 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_2_3 = Distribution_io_ProcessValid ? io_Stationary_matrix_2_3 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_2_4 = Distribution_io_ProcessValid ? io_Stationary_matrix_2_4 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_2_5 = Distribution_io_ProcessValid ? io_Stationary_matrix_2_5 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_2_6 = Distribution_io_ProcessValid ? io_Stationary_matrix_2_6 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_2_7 = Distribution_io_ProcessValid ? io_Stationary_matrix_2_7 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_3_0 = Distribution_io_ProcessValid ? io_Stationary_matrix_3_0 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_3_1 = Distribution_io_ProcessValid ? io_Stationary_matrix_3_1 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_3_2 = Distribution_io_ProcessValid ? io_Stationary_matrix_3_2 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_3_3 = Distribution_io_ProcessValid ? io_Stationary_matrix_3_3 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_3_4 = Distribution_io_ProcessValid ? io_Stationary_matrix_3_4 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_3_5 = Distribution_io_ProcessValid ? io_Stationary_matrix_3_5 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_3_6 = Distribution_io_ProcessValid ? io_Stationary_matrix_3_6 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_3_7 = Distribution_io_ProcessValid ? io_Stationary_matrix_3_7 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_4_0 = Distribution_io_ProcessValid ? io_Stationary_matrix_4_0 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_4_1 = Distribution_io_ProcessValid ? io_Stationary_matrix_4_1 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_4_2 = Distribution_io_ProcessValid ? io_Stationary_matrix_4_2 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_4_3 = Distribution_io_ProcessValid ? io_Stationary_matrix_4_3 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_4_4 = Distribution_io_ProcessValid ? io_Stationary_matrix_4_4 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_4_5 = Distribution_io_ProcessValid ? io_Stationary_matrix_4_5 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_4_6 = Distribution_io_ProcessValid ? io_Stationary_matrix_4_6 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_4_7 = Distribution_io_ProcessValid ? io_Stationary_matrix_4_7 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_5_0 = Distribution_io_ProcessValid ? io_Stationary_matrix_5_0 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_5_1 = Distribution_io_ProcessValid ? io_Stationary_matrix_5_1 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_5_2 = Distribution_io_ProcessValid ? io_Stationary_matrix_5_2 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_5_3 = Distribution_io_ProcessValid ? io_Stationary_matrix_5_3 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_5_4 = Distribution_io_ProcessValid ? io_Stationary_matrix_5_4 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_5_5 = Distribution_io_ProcessValid ? io_Stationary_matrix_5_5 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_5_6 = Distribution_io_ProcessValid ? io_Stationary_matrix_5_6 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_5_7 = Distribution_io_ProcessValid ? io_Stationary_matrix_5_7 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_6_0 = Distribution_io_ProcessValid ? io_Stationary_matrix_6_0 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_6_1 = Distribution_io_ProcessValid ? io_Stationary_matrix_6_1 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_6_2 = Distribution_io_ProcessValid ? io_Stationary_matrix_6_2 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_6_3 = Distribution_io_ProcessValid ? io_Stationary_matrix_6_3 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_6_4 = Distribution_io_ProcessValid ? io_Stationary_matrix_6_4 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_6_5 = Distribution_io_ProcessValid ? io_Stationary_matrix_6_5 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_6_6 = Distribution_io_ProcessValid ? io_Stationary_matrix_6_6 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_6_7 = Distribution_io_ProcessValid ? io_Stationary_matrix_6_7 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_7_0 = Distribution_io_ProcessValid ? io_Stationary_matrix_7_0 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_7_1 = Distribution_io_ProcessValid ? io_Stationary_matrix_7_1 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_7_2 = Distribution_io_ProcessValid ? io_Stationary_matrix_7_2 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_7_3 = Distribution_io_ProcessValid ? io_Stationary_matrix_7_3 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_7_4 = Distribution_io_ProcessValid ? io_Stationary_matrix_7_4 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_7_5 = Distribution_io_ProcessValid ? io_Stationary_matrix_7_5 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_7_6 = Distribution_io_ProcessValid ? io_Stationary_matrix_7_6 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat1_7_7 = Distribution_io_ProcessValid ? io_Stationary_matrix_7_7 : 16'h0; // @[PathFinder.scala 52:40 55:21 65:21]
  assign myMuxes_io_mat2_0 = Distribution_io_ProcessValid ? io_Streaming_matrix_0 : 16'h0; // @[PathFinder.scala 52:40 57:21 66:21]
  assign myMuxes_io_mat2_1 = Distribution_io_ProcessValid ? io_Streaming_matrix_1 : 16'h0; // @[PathFinder.scala 52:40 57:21 66:21]
  assign myMuxes_io_mat2_2 = Distribution_io_ProcessValid ? io_Streaming_matrix_2 : 16'h0; // @[PathFinder.scala 52:40 57:21 66:21]
  assign myMuxes_io_mat2_3 = Distribution_io_ProcessValid ? io_Streaming_matrix_3 : 16'h0; // @[PathFinder.scala 52:40 57:21 66:21]
  assign myMuxes_io_mat2_4 = Distribution_io_ProcessValid ? io_Streaming_matrix_4 : 16'h0; // @[PathFinder.scala 52:40 57:21 66:21]
  assign myMuxes_io_mat2_5 = Distribution_io_ProcessValid ? io_Streaming_matrix_5 : 16'h0; // @[PathFinder.scala 52:40 57:21 66:21]
  assign myMuxes_io_mat2_6 = Distribution_io_ProcessValid ? io_Streaming_matrix_6 : 16'h0; // @[PathFinder.scala 52:40 57:21 66:21]
  assign myMuxes_io_mat2_7 = Distribution_io_ProcessValid ? io_Streaming_matrix_7 : 16'h0; // @[PathFinder.scala 52:40 57:21 66:21]
  assign myMuxes_io_counterMatrix1_0_0 = _GEN_73[15:0];
  assign myMuxes_io_counterMatrix1_0_1 = _GEN_74[15:0];
  assign myMuxes_io_counterMatrix1_0_2 = _GEN_75[15:0];
  assign myMuxes_io_counterMatrix1_0_3 = _GEN_76[15:0];
  assign myMuxes_io_counterMatrix1_0_4 = _GEN_77[15:0];
  assign myMuxes_io_counterMatrix1_0_5 = _GEN_78[15:0];
  assign myMuxes_io_counterMatrix1_0_6 = _GEN_79[15:0];
  assign myMuxes_io_counterMatrix1_0_7 = _GEN_80[15:0];
  assign myMuxes_io_counterMatrix1_1_0 = _GEN_81[15:0];
  assign myMuxes_io_counterMatrix1_1_1 = _GEN_82[15:0];
  assign myMuxes_io_counterMatrix1_1_2 = _GEN_83[15:0];
  assign myMuxes_io_counterMatrix1_1_3 = _GEN_84[15:0];
  assign myMuxes_io_counterMatrix1_1_4 = _GEN_85[15:0];
  assign myMuxes_io_counterMatrix1_1_5 = _GEN_86[15:0];
  assign myMuxes_io_counterMatrix1_1_6 = _GEN_87[15:0];
  assign myMuxes_io_counterMatrix1_1_7 = _GEN_88[15:0];
  assign myMuxes_io_counterMatrix1_2_0 = _GEN_89[15:0];
  assign myMuxes_io_counterMatrix1_2_1 = _GEN_90[15:0];
  assign myMuxes_io_counterMatrix1_2_2 = _GEN_91[15:0];
  assign myMuxes_io_counterMatrix1_2_3 = _GEN_92[15:0];
  assign myMuxes_io_counterMatrix1_2_4 = _GEN_93[15:0];
  assign myMuxes_io_counterMatrix1_2_5 = _GEN_94[15:0];
  assign myMuxes_io_counterMatrix1_2_6 = _GEN_95[15:0];
  assign myMuxes_io_counterMatrix1_2_7 = _GEN_96[15:0];
  assign myMuxes_io_counterMatrix1_3_0 = _GEN_97[15:0];
  assign myMuxes_io_counterMatrix1_3_1 = _GEN_98[15:0];
  assign myMuxes_io_counterMatrix1_3_2 = _GEN_99[15:0];
  assign myMuxes_io_counterMatrix1_3_3 = _GEN_100[15:0];
  assign myMuxes_io_counterMatrix1_3_4 = _GEN_101[15:0];
  assign myMuxes_io_counterMatrix1_3_5 = _GEN_102[15:0];
  assign myMuxes_io_counterMatrix1_3_6 = _GEN_103[15:0];
  assign myMuxes_io_counterMatrix1_3_7 = _GEN_104[15:0];
  assign myMuxes_io_counterMatrix1_4_0 = _GEN_105[15:0];
  assign myMuxes_io_counterMatrix1_4_1 = _GEN_106[15:0];
  assign myMuxes_io_counterMatrix1_4_2 = _GEN_107[15:0];
  assign myMuxes_io_counterMatrix1_4_3 = _GEN_108[15:0];
  assign myMuxes_io_counterMatrix1_4_4 = _GEN_109[15:0];
  assign myMuxes_io_counterMatrix1_4_5 = _GEN_110[15:0];
  assign myMuxes_io_counterMatrix1_4_6 = _GEN_111[15:0];
  assign myMuxes_io_counterMatrix1_4_7 = _GEN_112[15:0];
  assign myMuxes_io_counterMatrix1_5_0 = _GEN_113[15:0];
  assign myMuxes_io_counterMatrix1_5_1 = _GEN_114[15:0];
  assign myMuxes_io_counterMatrix1_5_2 = _GEN_115[15:0];
  assign myMuxes_io_counterMatrix1_5_3 = _GEN_116[15:0];
  assign myMuxes_io_counterMatrix1_5_4 = _GEN_117[15:0];
  assign myMuxes_io_counterMatrix1_5_5 = _GEN_118[15:0];
  assign myMuxes_io_counterMatrix1_5_6 = _GEN_119[15:0];
  assign myMuxes_io_counterMatrix1_5_7 = _GEN_120[15:0];
  assign myMuxes_io_counterMatrix1_6_0 = _GEN_121[15:0];
  assign myMuxes_io_counterMatrix1_6_1 = _GEN_122[15:0];
  assign myMuxes_io_counterMatrix1_6_2 = _GEN_123[15:0];
  assign myMuxes_io_counterMatrix1_6_3 = _GEN_124[15:0];
  assign myMuxes_io_counterMatrix1_6_4 = _GEN_125[15:0];
  assign myMuxes_io_counterMatrix1_6_5 = _GEN_126[15:0];
  assign myMuxes_io_counterMatrix1_6_6 = _GEN_127[15:0];
  assign myMuxes_io_counterMatrix1_6_7 = _GEN_128[15:0];
  assign myMuxes_io_counterMatrix1_7_0 = _GEN_129[15:0];
  assign myMuxes_io_counterMatrix1_7_1 = _GEN_130[15:0];
  assign myMuxes_io_counterMatrix1_7_2 = _GEN_131[15:0];
  assign myMuxes_io_counterMatrix1_7_3 = _GEN_132[15:0];
  assign myMuxes_io_counterMatrix1_7_4 = _GEN_133[15:0];
  assign myMuxes_io_counterMatrix1_7_5 = _GEN_134[15:0];
  assign myMuxes_io_counterMatrix1_7_6 = _GEN_135[15:0];
  assign myMuxes_io_counterMatrix1_7_7 = _GEN_136[15:0];
  assign myMuxes_io_counterMatrix2_0 = Distribution_io_ProcessValid ? myCounter_io_counterMatrix2_bits_0 : 16'h0; // @[PathFinder.scala 52:40 59:31 68:31]
  assign myMuxes_io_counterMatrix2_1 = Distribution_io_ProcessValid ? myCounter_io_counterMatrix2_bits_1 : 16'h0; // @[PathFinder.scala 52:40 59:31 68:31]
  assign myMuxes_io_counterMatrix2_2 = Distribution_io_ProcessValid ? myCounter_io_counterMatrix2_bits_2 : 16'h0; // @[PathFinder.scala 52:40 59:31 68:31]
  assign myMuxes_io_counterMatrix2_3 = Distribution_io_ProcessValid ? myCounter_io_counterMatrix2_bits_3 : 16'h0; // @[PathFinder.scala 52:40 59:31 68:31]
  assign myMuxes_io_counterMatrix2_4 = Distribution_io_ProcessValid ? myCounter_io_counterMatrix2_bits_4 : 16'h0; // @[PathFinder.scala 52:40 59:31 68:31]
  assign myMuxes_io_counterMatrix2_5 = Distribution_io_ProcessValid ? myCounter_io_counterMatrix2_bits_5 : 16'h0; // @[PathFinder.scala 52:40 59:31 68:31]
  assign myMuxes_io_counterMatrix2_6 = Distribution_io_ProcessValid ? myCounter_io_counterMatrix2_bits_6 : 16'h0; // @[PathFinder.scala 52:40 59:31 68:31]
  assign myMuxes_io_counterMatrix2_7 = Distribution_io_ProcessValid ? myCounter_io_counterMatrix2_bits_7 : 16'h0; // @[PathFinder.scala 52:40 59:31 68:31]
  assign myCounter_clock = clock;
  assign myCounter_reset = reset;
  assign myCounter_io_Stationary_matrix_0_0 = io_Stationary_matrix_0_0; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_0_1 = io_Stationary_matrix_0_1; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_0_2 = io_Stationary_matrix_0_2; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_0_3 = io_Stationary_matrix_0_3; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_0_4 = io_Stationary_matrix_0_4; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_0_5 = io_Stationary_matrix_0_5; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_0_6 = io_Stationary_matrix_0_6; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_0_7 = io_Stationary_matrix_0_7; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_1_0 = io_Stationary_matrix_1_0; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_1_1 = io_Stationary_matrix_1_1; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_1_2 = io_Stationary_matrix_1_2; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_1_3 = io_Stationary_matrix_1_3; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_1_4 = io_Stationary_matrix_1_4; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_1_5 = io_Stationary_matrix_1_5; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_1_6 = io_Stationary_matrix_1_6; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_1_7 = io_Stationary_matrix_1_7; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_2_0 = io_Stationary_matrix_2_0; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_2_1 = io_Stationary_matrix_2_1; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_2_2 = io_Stationary_matrix_2_2; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_2_3 = io_Stationary_matrix_2_3; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_2_4 = io_Stationary_matrix_2_4; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_2_5 = io_Stationary_matrix_2_5; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_2_6 = io_Stationary_matrix_2_6; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_2_7 = io_Stationary_matrix_2_7; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_3_0 = io_Stationary_matrix_3_0; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_3_1 = io_Stationary_matrix_3_1; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_3_2 = io_Stationary_matrix_3_2; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_3_3 = io_Stationary_matrix_3_3; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_3_4 = io_Stationary_matrix_3_4; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_3_5 = io_Stationary_matrix_3_5; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_3_6 = io_Stationary_matrix_3_6; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_3_7 = io_Stationary_matrix_3_7; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_4_0 = io_Stationary_matrix_4_0; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_4_1 = io_Stationary_matrix_4_1; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_4_2 = io_Stationary_matrix_4_2; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_4_3 = io_Stationary_matrix_4_3; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_4_4 = io_Stationary_matrix_4_4; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_4_5 = io_Stationary_matrix_4_5; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_4_6 = io_Stationary_matrix_4_6; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_4_7 = io_Stationary_matrix_4_7; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_5_0 = io_Stationary_matrix_5_0; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_5_1 = io_Stationary_matrix_5_1; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_5_2 = io_Stationary_matrix_5_2; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_5_3 = io_Stationary_matrix_5_3; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_5_4 = io_Stationary_matrix_5_4; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_5_5 = io_Stationary_matrix_5_5; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_5_6 = io_Stationary_matrix_5_6; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_5_7 = io_Stationary_matrix_5_7; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_6_0 = io_Stationary_matrix_6_0; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_6_1 = io_Stationary_matrix_6_1; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_6_2 = io_Stationary_matrix_6_2; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_6_3 = io_Stationary_matrix_6_3; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_6_4 = io_Stationary_matrix_6_4; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_6_5 = io_Stationary_matrix_6_5; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_6_6 = io_Stationary_matrix_6_6; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_6_7 = io_Stationary_matrix_6_7; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_7_0 = io_Stationary_matrix_7_0; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_7_1 = io_Stationary_matrix_7_1; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_7_2 = io_Stationary_matrix_7_2; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_7_3 = io_Stationary_matrix_7_3; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_7_4 = io_Stationary_matrix_7_4; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_7_5 = io_Stationary_matrix_7_5; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_7_6 = io_Stationary_matrix_7_6; // @[PathFinder.scala 34:34]
  assign myCounter_io_Stationary_matrix_7_7 = io_Stationary_matrix_7_7; // @[PathFinder.scala 34:34]
  assign myCounter_io_Streaming_matrix_0 = io_Streaming_matrix_0; // @[PathFinder.scala 35:33]
  assign myCounter_io_Streaming_matrix_1 = io_Streaming_matrix_1; // @[PathFinder.scala 35:33]
  assign myCounter_io_Streaming_matrix_2 = io_Streaming_matrix_2; // @[PathFinder.scala 35:33]
  assign myCounter_io_Streaming_matrix_3 = io_Streaming_matrix_3; // @[PathFinder.scala 35:33]
  assign myCounter_io_Streaming_matrix_4 = io_Streaming_matrix_4; // @[PathFinder.scala 35:33]
  assign myCounter_io_Streaming_matrix_5 = io_Streaming_matrix_5; // @[PathFinder.scala 35:33]
  assign myCounter_io_Streaming_matrix_6 = io_Streaming_matrix_6; // @[PathFinder.scala 35:33]
  assign myCounter_io_Streaming_matrix_7 = io_Streaming_matrix_7; // @[PathFinder.scala 35:33]
  assign myCounter_io_start = myCounter_io_start_REG; // @[PathFinder.scala 33:22]
  assign Distribution_clock = clock;
  assign Distribution_reset = reset;
  assign Distribution_io_matrix_0_0 = {{16'd0}, myCounter_io_counterMatrix1_bits_0_0}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_0_1 = {{16'd0}, myCounter_io_counterMatrix1_bits_0_1}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_0_2 = {{16'd0}, myCounter_io_counterMatrix1_bits_0_2}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_0_3 = {{16'd0}, myCounter_io_counterMatrix1_bits_0_3}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_0_4 = {{16'd0}, myCounter_io_counterMatrix1_bits_0_4}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_0_5 = {{16'd0}, myCounter_io_counterMatrix1_bits_0_5}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_0_6 = {{16'd0}, myCounter_io_counterMatrix1_bits_0_6}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_0_7 = {{16'd0}, myCounter_io_counterMatrix1_bits_0_7}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_1_0 = {{16'd0}, myCounter_io_counterMatrix1_bits_1_0}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_1_1 = {{16'd0}, myCounter_io_counterMatrix1_bits_1_1}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_1_2 = {{16'd0}, myCounter_io_counterMatrix1_bits_1_2}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_1_3 = {{16'd0}, myCounter_io_counterMatrix1_bits_1_3}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_1_4 = {{16'd0}, myCounter_io_counterMatrix1_bits_1_4}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_1_5 = {{16'd0}, myCounter_io_counterMatrix1_bits_1_5}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_1_6 = {{16'd0}, myCounter_io_counterMatrix1_bits_1_6}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_1_7 = {{16'd0}, myCounter_io_counterMatrix1_bits_1_7}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_2_0 = {{16'd0}, myCounter_io_counterMatrix1_bits_2_0}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_2_1 = {{16'd0}, myCounter_io_counterMatrix1_bits_2_1}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_2_2 = {{16'd0}, myCounter_io_counterMatrix1_bits_2_2}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_2_3 = {{16'd0}, myCounter_io_counterMatrix1_bits_2_3}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_2_4 = {{16'd0}, myCounter_io_counterMatrix1_bits_2_4}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_2_5 = {{16'd0}, myCounter_io_counterMatrix1_bits_2_5}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_2_6 = {{16'd0}, myCounter_io_counterMatrix1_bits_2_6}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_2_7 = {{16'd0}, myCounter_io_counterMatrix1_bits_2_7}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_3_0 = {{16'd0}, myCounter_io_counterMatrix1_bits_3_0}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_3_1 = {{16'd0}, myCounter_io_counterMatrix1_bits_3_1}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_3_2 = {{16'd0}, myCounter_io_counterMatrix1_bits_3_2}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_3_3 = {{16'd0}, myCounter_io_counterMatrix1_bits_3_3}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_3_4 = {{16'd0}, myCounter_io_counterMatrix1_bits_3_4}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_3_5 = {{16'd0}, myCounter_io_counterMatrix1_bits_3_5}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_3_6 = {{16'd0}, myCounter_io_counterMatrix1_bits_3_6}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_3_7 = {{16'd0}, myCounter_io_counterMatrix1_bits_3_7}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_4_0 = {{16'd0}, myCounter_io_counterMatrix1_bits_4_0}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_4_1 = {{16'd0}, myCounter_io_counterMatrix1_bits_4_1}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_4_2 = {{16'd0}, myCounter_io_counterMatrix1_bits_4_2}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_4_3 = {{16'd0}, myCounter_io_counterMatrix1_bits_4_3}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_4_4 = {{16'd0}, myCounter_io_counterMatrix1_bits_4_4}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_4_5 = {{16'd0}, myCounter_io_counterMatrix1_bits_4_5}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_4_6 = {{16'd0}, myCounter_io_counterMatrix1_bits_4_6}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_4_7 = {{16'd0}, myCounter_io_counterMatrix1_bits_4_7}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_5_0 = {{16'd0}, myCounter_io_counterMatrix1_bits_5_0}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_5_1 = {{16'd0}, myCounter_io_counterMatrix1_bits_5_1}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_5_2 = {{16'd0}, myCounter_io_counterMatrix1_bits_5_2}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_5_3 = {{16'd0}, myCounter_io_counterMatrix1_bits_5_3}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_5_4 = {{16'd0}, myCounter_io_counterMatrix1_bits_5_4}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_5_5 = {{16'd0}, myCounter_io_counterMatrix1_bits_5_5}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_5_6 = {{16'd0}, myCounter_io_counterMatrix1_bits_5_6}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_5_7 = {{16'd0}, myCounter_io_counterMatrix1_bits_5_7}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_6_0 = {{16'd0}, myCounter_io_counterMatrix1_bits_6_0}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_6_1 = {{16'd0}, myCounter_io_counterMatrix1_bits_6_1}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_6_2 = {{16'd0}, myCounter_io_counterMatrix1_bits_6_2}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_6_3 = {{16'd0}, myCounter_io_counterMatrix1_bits_6_3}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_6_4 = {{16'd0}, myCounter_io_counterMatrix1_bits_6_4}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_6_5 = {{16'd0}, myCounter_io_counterMatrix1_bits_6_5}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_6_6 = {{16'd0}, myCounter_io_counterMatrix1_bits_6_6}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_6_7 = {{16'd0}, myCounter_io_counterMatrix1_bits_6_7}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_7_0 = {{16'd0}, myCounter_io_counterMatrix1_bits_7_0}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_7_1 = {{16'd0}, myCounter_io_counterMatrix1_bits_7_1}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_7_2 = {{16'd0}, myCounter_io_counterMatrix1_bits_7_2}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_7_3 = {{16'd0}, myCounter_io_counterMatrix1_bits_7_3}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_7_4 = {{16'd0}, myCounter_io_counterMatrix1_bits_7_4}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_7_5 = {{16'd0}, myCounter_io_counterMatrix1_bits_7_5}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_7_6 = {{16'd0}, myCounter_io_counterMatrix1_bits_7_6}; // @[PathFinder.scala 43:26]
  assign Distribution_io_matrix_7_7 = {{16'd0}, myCounter_io_counterMatrix1_bits_7_7}; // @[PathFinder.scala 43:26]
  assign Distribution_io_s = io_NoDPE; // @[PathFinder.scala 40:21]
  assign Distribution_io_valid = myCounter_io_valid; // @[PathFinder.scala 39:25]
  always @(posedge clock) begin
    myCounter_io_start_REG <= io_DataValid; // @[PathFinder.scala 33:32]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  myCounter_io_start_REG = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module fancontrol4(
  input        clock,
  input        reset,
  input        io_i_data_valid,
  output       io_o_reduction_add_0,
  output       io_o_reduction_add_1,
  output       io_o_reduction_add_2,
  output [2:0] io_o_reduction_cmd_0,
  output [2:0] io_o_reduction_cmd_1,
  output [2:0] io_o_reduction_cmd_2,
  output       io_o_reduction_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
`endif // RANDOMIZE_REG_INIT
  reg  r_reduction_add_0; // @[FanCtrl.scala 19:34]
  reg  r_reduction_add_1; // @[FanCtrl.scala 19:34]
  reg  r_reduction_add_2; // @[FanCtrl.scala 19:34]
  reg [2:0] r_reduction_cmd_0; // @[FanCtrl.scala 20:34]
  reg [2:0] r_reduction_cmd_1; // @[FanCtrl.scala 20:34]
  reg [2:0] r_reduction_cmd_2; // @[FanCtrl.scala 20:34]
  reg  r_add_lvl_0Reg_6; // @[FanCtrl.scala 23:33]
  reg  r_add_lvl_0Reg_7; // @[FanCtrl.scala 23:33]
  reg  r_add_lvl_1Reg_4; // @[FanCtrl.scala 24:33]
  reg [2:0] r_cmd_lvl_0Reg_6; // @[FanCtrl.scala 27:33]
  reg [2:0] r_cmd_lvl_0Reg_7; // @[FanCtrl.scala 27:33]
  reg [2:0] r_cmd_lvl_1Reg_4; // @[FanCtrl.scala 28:33]
  reg [4:0] w_vn_0; // @[FanCtrl.scala 34:23]
  reg [4:0] w_vn_1; // @[FanCtrl.scala 34:23]
  reg [4:0] w_vn_2; // @[FanCtrl.scala 34:23]
  reg [4:0] w_vn_3; // @[FanCtrl.scala 34:23]
  reg  r_valid_0; // @[FanCtrl.scala 35:26]
  reg  r_valid_1; // @[FanCtrl.scala 35:26]
  reg  r_valid_2; // @[FanCtrl.scala 35:26]
  reg  r_valid_3; // @[FanCtrl.scala 35:26]
  wire [2:0] _T_2 = 2'h2 * 1'h0; // @[FanCtrl.scala 42:25]
  wire [3:0] _T_3 = {{1'd0}, _T_2}; // @[FanCtrl.scala 42:31]
  wire [2:0] _T_8 = _T_2 + 3'h1; // @[FanCtrl.scala 42:58]
  wire [4:0] _GEN_1 = 2'h1 == _T_3[1:0] ? w_vn_1 : w_vn_0; // @[FanCtrl.scala 42:{39,39}]
  wire [4:0] _GEN_2 = 2'h2 == _T_3[1:0] ? w_vn_2 : _GEN_1; // @[FanCtrl.scala 42:{39,39}]
  wire [4:0] _GEN_3 = 2'h3 == _T_3[1:0] ? w_vn_3 : _GEN_2; // @[FanCtrl.scala 42:{39,39}]
  wire [4:0] _GEN_5 = 2'h1 == _T_8[1:0] ? w_vn_1 : w_vn_0; // @[FanCtrl.scala 42:{39,39}]
  wire [4:0] _GEN_6 = 2'h2 == _T_8[1:0] ? w_vn_2 : _GEN_5; // @[FanCtrl.scala 42:{39,39}]
  wire [4:0] _GEN_7 = 2'h3 == _T_8[1:0] ? w_vn_3 : _GEN_6; // @[FanCtrl.scala 42:{39,39}]
  wire  _T_10 = _GEN_3 == _GEN_7; // @[FanCtrl.scala 42:39]
  wire [2:0] _T_21 = _T_2 + 3'h2; // @[FanCtrl.scala 49:32]
  wire [4:0] _GEN_22 = 2'h1 == _T_21[1:0] ? w_vn_1 : w_vn_0; // @[FanCtrl.scala 48:{41,41}]
  wire [4:0] _GEN_23 = 2'h2 == _T_21[1:0] ? w_vn_2 : _GEN_22; // @[FanCtrl.scala 48:{41,41}]
  wire [4:0] _GEN_24 = 2'h3 == _T_21[1:0] ? w_vn_3 : _GEN_23; // @[FanCtrl.scala 48:{41,41}]
  wire  _T_23 = _GEN_7 != _GEN_24; // @[FanCtrl.scala 48:41]
  wire  _T_32 = _GEN_3 != _GEN_7; // @[FanCtrl.scala 50:41]
  wire  _T_33 = _T_23 & _T_32; // @[FanCtrl.scala 49:41]
  wire  _T_42 = _GEN_7 == _GEN_24; // @[FanCtrl.scala 55:48]
  wire  _T_52 = _T_42 & _T_32; // @[FanCtrl.scala 56:46]
  wire [1:0] _GEN_49 = _T_52 ? 2'h3 : 2'h0; // @[FanCtrl.scala 58:48 60:40 63:38]
  wire  _GEN_54 = r_valid_1 & _T_10; // @[FanCtrl.scala 41:34]
  wire [2:0] _T_113 = 2'h2 * 1'h1; // @[FanCtrl.scala 42:25]
  wire [3:0] _T_114 = {{1'd0}, _T_113}; // @[FanCtrl.scala 42:31]
  wire [2:0] _T_119 = _T_113 + 3'h1; // @[FanCtrl.scala 42:58]
  wire [4:0] _GEN_124 = 2'h1 == _T_114[1:0] ? w_vn_1 : w_vn_0; // @[FanCtrl.scala 42:{39,39}]
  wire [4:0] _GEN_125 = 2'h2 == _T_114[1:0] ? w_vn_2 : _GEN_124; // @[FanCtrl.scala 42:{39,39}]
  wire [4:0] _GEN_126 = 2'h3 == _T_114[1:0] ? w_vn_3 : _GEN_125; // @[FanCtrl.scala 42:{39,39}]
  wire [4:0] _GEN_128 = 2'h1 == _T_119[1:0] ? w_vn_1 : w_vn_0; // @[FanCtrl.scala 42:{39,39}]
  wire [4:0] _GEN_129 = 2'h2 == _T_119[1:0] ? w_vn_2 : _GEN_128; // @[FanCtrl.scala 42:{39,39}]
  wire [4:0] _GEN_130 = 2'h3 == _T_119[1:0] ? w_vn_3 : _GEN_129; // @[FanCtrl.scala 42:{39,39}]
  wire  _T_121 = _GEN_126 == _GEN_130; // @[FanCtrl.scala 42:39]
  wire  _T_143 = _GEN_126 != _GEN_130; // @[FanCtrl.scala 50:41]
  wire  _GEN_178 = r_valid_1 & _T_121; // @[FanCtrl.scala 41:34]
  wire [2:0] _T_188 = _T_113 - 3'h1; // @[FanCtrl.scala 88:58]
  wire [4:0] _GEN_206 = 2'h1 == _T_188[1:0] ? w_vn_1 : w_vn_0; // @[FanCtrl.scala 88:{39,39}]
  wire [4:0] _GEN_207 = 2'h2 == _T_188[1:0] ? w_vn_2 : _GEN_206; // @[FanCtrl.scala 88:{39,39}]
  wire [4:0] _GEN_208 = 2'h3 == _T_188[1:0] ? w_vn_3 : _GEN_207; // @[FanCtrl.scala 88:{39,39}]
  wire  _T_200 = _GEN_126 != _GEN_208 & _T_143; // @[FanCtrl.scala 88:67]
  wire  _T_219 = _GEN_126 == _GEN_208 & _T_143; // @[FanCtrl.scala 93:73]
  wire [3:0] _T_228 = 3'h4 * 1'h0; // @[FanCtrl.scala 117:23]
  wire [3:0] _T_230 = _T_228 + 4'h1; // @[FanCtrl.scala 117:29]
  wire [3:0] _T_234 = _T_228 + 4'h2; // @[FanCtrl.scala 117:56]
  wire [4:0] _GEN_254 = 2'h1 == _T_230[1:0] ? w_vn_1 : w_vn_0; // @[FanCtrl.scala 117:{37,37}]
  wire [4:0] _GEN_255 = 2'h2 == _T_230[1:0] ? w_vn_2 : _GEN_254; // @[FanCtrl.scala 117:{37,37}]
  wire [4:0] _GEN_256 = 2'h3 == _T_230[1:0] ? w_vn_3 : _GEN_255; // @[FanCtrl.scala 117:{37,37}]
  wire [4:0] _GEN_258 = 2'h1 == _T_234[1:0] ? w_vn_1 : w_vn_0; // @[FanCtrl.scala 117:{37,37}]
  wire [4:0] _GEN_259 = 2'h2 == _T_234[1:0] ? w_vn_2 : _GEN_258; // @[FanCtrl.scala 117:{37,37}]
  wire [4:0] _GEN_260 = 2'h3 == _T_234[1:0] ? w_vn_3 : _GEN_259; // @[FanCtrl.scala 117:{37,37}]
  wire  _T_236 = _GEN_256 == _GEN_260; // @[FanCtrl.scala 117:37]
  wire [4:0] _T_242 = {{1'd0}, _T_228}; // @[FanCtrl.scala 123:30]
  wire [4:0] _GEN_271 = 2'h1 == _T_242[1:0] ? w_vn_1 : w_vn_0; // @[FanCtrl.scala 123:{38,38}]
  wire [4:0] _GEN_272 = 2'h2 == _T_242[1:0] ? w_vn_2 : _GEN_271; // @[FanCtrl.scala 123:{38,38}]
  wire [4:0] _GEN_273 = 2'h3 == _T_242[1:0] ? w_vn_3 : _GEN_272; // @[FanCtrl.scala 123:{38,38}]
  wire  _T_249 = _GEN_273 == _GEN_256; // @[FanCtrl.scala 123:38]
  wire [3:0] _T_256 = _T_228 + 4'h3; // @[FanCtrl.scala 124:55]
  wire [4:0] _GEN_283 = 2'h1 == _T_256[1:0] ? w_vn_1 : w_vn_0; // @[FanCtrl.scala 124:{36,36}]
  wire [4:0] _GEN_284 = 2'h2 == _T_256[1:0] ? w_vn_2 : _GEN_283; // @[FanCtrl.scala 124:{36,36}]
  wire [4:0] _GEN_285 = 2'h3 == _T_256[1:0] ? w_vn_3 : _GEN_284; // @[FanCtrl.scala 124:{36,36}]
  wire  _T_258 = _GEN_260 == _GEN_285; // @[FanCtrl.scala 124:36]
  wire  _T_259 = _GEN_273 == _GEN_256 & _T_258; // @[FanCtrl.scala 123:65]
  wire [3:0] _T_262 = _T_228 + 4'h4; // @[FanCtrl.scala 125:29]
  wire [4:0] _GEN_287 = 2'h1 == _T_262[1:0] ? w_vn_1 : w_vn_0; // @[FanCtrl.scala 125:{37,37}]
  wire [4:0] _GEN_288 = 2'h2 == _T_262[1:0] ? w_vn_2 : _GEN_287; // @[FanCtrl.scala 125:{37,37}]
  wire [4:0] _GEN_289 = 2'h3 == _T_262[1:0] ? w_vn_3 : _GEN_288; // @[FanCtrl.scala 125:{37,37}]
  wire  _T_268 = _GEN_289 != _GEN_285; // @[FanCtrl.scala 125:37]
  wire  _T_269 = _T_259 & _T_268; // @[FanCtrl.scala 124:64]
  wire  _T_278 = _GEN_256 != _GEN_260; // @[FanCtrl.scala 126:37]
  wire  _T_279 = _T_269 & _T_278; // @[FanCtrl.scala 125:64]
  wire  _T_300 = _T_258 & _T_268; // @[FanCtrl.scala 130:71]
  wire  _T_310 = _T_300 & _T_278; // @[FanCtrl.scala 131:71]
  wire  _T_331 = _T_249 & _T_278; // @[FanCtrl.scala 136:71]
  wire [2:0] _GEN_356 = _T_331 ? 3'h3 : 3'h0; // @[FanCtrl.scala 137:72]
  wire  _GEN_371 = r_valid_1 & _T_236; // @[FanCtrl.scala 116:32]
  assign io_o_reduction_add_0 = r_add_lvl_0Reg_6; // @[FanCtrl.scala 227:{35,35}]
  assign io_o_reduction_add_1 = r_add_lvl_0Reg_7; // @[FanCtrl.scala 227:{35,35}]
  assign io_o_reduction_add_2 = r_add_lvl_1Reg_4; // @[FanCtrl.scala 227:{35,35}]
  assign io_o_reduction_cmd_0 = r_cmd_lvl_0Reg_6; // @[FanCtrl.scala 236:{34,34}]
  assign io_o_reduction_cmd_1 = r_cmd_lvl_0Reg_7; // @[FanCtrl.scala 236:{34,34}]
  assign io_o_reduction_cmd_2 = r_cmd_lvl_1Reg_4; // @[FanCtrl.scala 236:{34,34}]
  assign io_o_reduction_valid = r_valid_3; // @[FanCtrl.scala 226:26]
  always @(posedge clock) begin
    if (reset) begin // @[FanCtrl.scala 19:34]
      r_reduction_add_0 <= 1'h0; // @[FanCtrl.scala 19:34]
    end else begin
      r_reduction_add_0 <= _GEN_54;
    end
    if (reset) begin // @[FanCtrl.scala 19:34]
      r_reduction_add_1 <= 1'h0; // @[FanCtrl.scala 19:34]
    end else begin
      r_reduction_add_1 <= _GEN_178;
    end
    if (reset) begin // @[FanCtrl.scala 19:34]
      r_reduction_add_2 <= 1'h0; // @[FanCtrl.scala 19:34]
    end else begin
      r_reduction_add_2 <= _GEN_371;
    end
    if (reset) begin // @[FanCtrl.scala 20:34]
      r_reduction_cmd_0 <= 3'h0; // @[FanCtrl.scala 20:34]
    end else if (r_valid_1) begin // @[FanCtrl.scala 41:34]
      if (_T_33) begin // @[FanCtrl.scala 51:42]
        r_reduction_cmd_0 <= 3'h5; // @[FanCtrl.scala 53:37]
      end else begin
        r_reduction_cmd_0 <= {{1'd0}, _GEN_49};
      end
    end else begin
      r_reduction_cmd_0 <= 3'h0; // @[FanCtrl.scala 68:33]
    end
    if (reset) begin // @[FanCtrl.scala 20:34]
      r_reduction_cmd_1 <= 3'h0; // @[FanCtrl.scala 20:34]
    end else if (r_valid_1) begin // @[FanCtrl.scala 81:34]
      if (_T_200) begin // @[FanCtrl.scala 89:66]
        r_reduction_cmd_1 <= 3'h5; // @[FanCtrl.scala 91:36]
      end else if (_T_219) begin // @[FanCtrl.scala 94:66]
        r_reduction_cmd_1 <= 3'h4; // @[FanCtrl.scala 96:35]
      end else begin
        r_reduction_cmd_1 <= 3'h0; // @[FanCtrl.scala 99:35]
      end
    end else begin
      r_reduction_cmd_1 <= 3'h0; // @[FanCtrl.scala 103:33]
    end
    if (reset) begin // @[FanCtrl.scala 20:34]
      r_reduction_cmd_2 <= 3'h0; // @[FanCtrl.scala 20:34]
    end else if (r_valid_1) begin // @[FanCtrl.scala 116:32]
      if (_T_279) begin // @[FanCtrl.scala 126:66]
        r_reduction_cmd_2 <= 3'h5;
      end else if (_T_310) begin // @[FanCtrl.scala 132:72]
        r_reduction_cmd_2 <= 3'h4;
      end else begin
        r_reduction_cmd_2 <= _GEN_356;
      end
    end else begin
      r_reduction_cmd_2 <= 3'h0;
    end
    if (reset) begin // @[FanCtrl.scala 23:33]
      r_add_lvl_0Reg_6 <= 1'h0; // @[FanCtrl.scala 23:33]
    end else begin
      r_add_lvl_0Reg_6 <= r_reduction_add_0; // @[FanCtrl.scala 157:20]
    end
    if (reset) begin // @[FanCtrl.scala 23:33]
      r_add_lvl_0Reg_7 <= 1'h0; // @[FanCtrl.scala 23:33]
    end else begin
      r_add_lvl_0Reg_7 <= r_reduction_add_1; // @[FanCtrl.scala 157:20]
    end
    if (reset) begin // @[FanCtrl.scala 24:33]
      r_add_lvl_1Reg_4 <= 1'h0; // @[FanCtrl.scala 24:33]
    end else begin
      r_add_lvl_1Reg_4 <= r_reduction_add_2; // @[FanCtrl.scala 168:20]
    end
    if (reset) begin // @[FanCtrl.scala 27:33]
      r_cmd_lvl_0Reg_6 <= 3'h0; // @[FanCtrl.scala 27:33]
    end else begin
      r_cmd_lvl_0Reg_6 <= r_reduction_cmd_0; // @[FanCtrl.scala 185:20]
    end
    if (reset) begin // @[FanCtrl.scala 27:33]
      r_cmd_lvl_0Reg_7 <= 3'h0; // @[FanCtrl.scala 27:33]
    end else begin
      r_cmd_lvl_0Reg_7 <= r_reduction_cmd_1; // @[FanCtrl.scala 185:20]
    end
    if (reset) begin // @[FanCtrl.scala 28:33]
      r_cmd_lvl_1Reg_4 <= 3'h0; // @[FanCtrl.scala 28:33]
    end else begin
      r_cmd_lvl_1Reg_4 <= r_reduction_cmd_2; // @[FanCtrl.scala 199:20]
    end
    if (reset) begin // @[FanCtrl.scala 34:23]
      w_vn_0 <= 5'h0; // @[FanCtrl.scala 34:23]
    end else begin
      w_vn_0 <= 5'h1; // @[FanCtrl.scala 37:10]
    end
    if (reset) begin // @[FanCtrl.scala 34:23]
      w_vn_1 <= 5'h0; // @[FanCtrl.scala 34:23]
    end else begin
      w_vn_1 <= 5'h1; // @[FanCtrl.scala 37:10]
    end
    if (reset) begin // @[FanCtrl.scala 34:23]
      w_vn_2 <= 5'h0; // @[FanCtrl.scala 34:23]
    end else begin
      w_vn_2 <= 5'h1; // @[FanCtrl.scala 37:10]
    end
    if (reset) begin // @[FanCtrl.scala 34:23]
      w_vn_3 <= 5'h0; // @[FanCtrl.scala 34:23]
    end else begin
      w_vn_3 <= 5'h1; // @[FanCtrl.scala 37:10]
    end
    if (reset) begin // @[FanCtrl.scala 35:26]
      r_valid_0 <= 1'h0; // @[FanCtrl.scala 35:26]
    end else begin
      r_valid_0 <= io_i_data_valid;
    end
    if (reset) begin // @[FanCtrl.scala 35:26]
      r_valid_1 <= 1'h0; // @[FanCtrl.scala 35:26]
    end else begin
      r_valid_1 <= r_valid_0; // @[FanCtrl.scala 222:24]
    end
    if (reset) begin // @[FanCtrl.scala 35:26]
      r_valid_2 <= 1'h0; // @[FanCtrl.scala 35:26]
    end else begin
      r_valid_2 <= r_valid_1; // @[FanCtrl.scala 222:24]
    end
    if (reset) begin // @[FanCtrl.scala 35:26]
      r_valid_3 <= 1'h0; // @[FanCtrl.scala 35:26]
    end else begin
      r_valid_3 <= r_valid_2; // @[FanCtrl.scala 222:24]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_reduction_add_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  r_reduction_add_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  r_reduction_add_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  r_reduction_cmd_0 = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  r_reduction_cmd_1 = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  r_reduction_cmd_2 = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  r_add_lvl_0Reg_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  r_add_lvl_0Reg_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  r_add_lvl_1Reg_4 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  r_cmd_lvl_0Reg_6 = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  r_cmd_lvl_0Reg_7 = _RAND_10[2:0];
  _RAND_11 = {1{`RANDOM}};
  r_cmd_lvl_1Reg_4 = _RAND_11[2:0];
  _RAND_12 = {1{`RANDOM}};
  w_vn_0 = _RAND_12[4:0];
  _RAND_13 = {1{`RANDOM}};
  w_vn_1 = _RAND_13[4:0];
  _RAND_14 = {1{`RANDOM}};
  w_vn_2 = _RAND_14[4:0];
  _RAND_15 = {1{`RANDOM}};
  w_vn_3 = _RAND_15[4:0];
  _RAND_16 = {1{`RANDOM}};
  r_valid_0 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  r_valid_1 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  r_valid_2 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  r_valid_3 = _RAND_19[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Benes(
  input  [15:0] io_i_data_bus2_0,
  input  [15:0] io_i_data_bus2_1,
  input  [15:0] io_i_data_bus2_2,
  input  [15:0] io_i_data_bus2_3,
  input  [15:0] io_i_data_bus1_0,
  input  [15:0] io_i_data_bus1_1,
  input  [15:0] io_i_data_bus1_2,
  input  [15:0] io_i_data_bus1_3,
  input  [3:0]  io_i_mux_bus_0,
  input  [3:0]  io_i_mux_bus_1,
  input  [3:0]  io_i_mux_bus_2,
  input  [3:0]  io_i_mux_bus_3,
  output [15:0] io_o_dist_bus1_0,
  output [15:0] io_o_dist_bus1_1,
  output [15:0] io_o_dist_bus1_2,
  output [15:0] io_o_dist_bus1_3,
  output [15:0] io_o_dist_bus2_0,
  output [15:0] io_o_dist_bus2_1,
  output [15:0] io_o_dist_bus2_2,
  output [15:0] io_o_dist_bus2_3
);
  wire  _T_2 = io_i_data_bus2_1 == io_i_data_bus2_0; // @[Benes.scala 60:36]
  wire [1:0] _GEN_4 = 2'h0 % 2'h2; // @[Benes.scala 24:52]
  wire  parsedindexvalue_first_stage = io_i_mux_bus_1[0] & (~_GEN_4[0] | 1'h0 - 1'h1); // @[Benes.scala 24:26]
  wire  parsedindexvalue_boolArray__0 = io_i_mux_bus_1[1]; // @[Benes.scala 28:92]
  wire  parsedindexvalue_boolArray__1 = io_i_mux_bus_1[2]; // @[Benes.scala 28:92]
  wire [2:0] _GEN_9 = {{2'd0}, parsedindexvalue_first_stage}; // @[Benes.scala 33:40]
  wire [2:0] _GEN_14 = _GEN_9 % 3'h4; // @[Benes.scala 33:40]
  wire  parsedindexvalue_calculation = _GEN_14[0]; // @[Benes.scala 33:40]
  wire  _parsedindexvalue_nextIndex_T = ~parsedindexvalue_calculation; // @[Benes.scala 35:27]
  wire  _parsedindexvalue_nextIndex_T_1 = ~parsedindexvalue_boolArray__0; // @[Benes.scala 35:53]
  wire  _parsedindexvalue_nextIndex_T_2 = ~parsedindexvalue_calculation & ~parsedindexvalue_boolArray__0; // @[Benes.scala 35:36]
  wire  _parsedindexvalue_nextIndex_T_5 = parsedindexvalue_calculation & _parsedindexvalue_nextIndex_T_1; // @[Benes.scala 36:36]
  wire [1:0] _GEN_88 = {{1'd0}, parsedindexvalue_calculation}; // @[Benes.scala 37:27]
  wire  _parsedindexvalue_nextIndex_T_6 = _GEN_88 == 2'h2; // @[Benes.scala 37:27]
  wire  _parsedindexvalue_nextIndex_T_8 = _GEN_88 == 2'h2 & _parsedindexvalue_nextIndex_T_1; // @[Benes.scala 37:36]
  wire  _parsedindexvalue_nextIndex_T_9 = _GEN_88 == 2'h3; // @[Benes.scala 38:27]
  wire  _parsedindexvalue_nextIndex_T_11 = _GEN_88 == 2'h3 & _parsedindexvalue_nextIndex_T_1; // @[Benes.scala 38:36]
  wire  _parsedindexvalue_nextIndex_T_14 = _parsedindexvalue_nextIndex_T & parsedindexvalue_boolArray__0; // @[Benes.scala 39:36]
  wire [1:0] _GEN_90 = {{1'd0}, parsedindexvalue_first_stage}; // @[Benes.scala 39:76]
  wire [1:0] _parsedindexvalue_nextIndex_T_16 = _GEN_90 + 2'h2; // @[Benes.scala 39:76]
  wire  _parsedindexvalue_nextIndex_T_19 = parsedindexvalue_calculation & parsedindexvalue_boolArray__0; // @[Benes.scala 40:36]
  wire  _parsedindexvalue_nextIndex_T_24 = _parsedindexvalue_nextIndex_T_6 & parsedindexvalue_boolArray__0; // @[Benes.scala 41:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_26 = _GEN_90 - 2'h2; // @[Benes.scala 41:76]
  wire  _parsedindexvalue_nextIndex_T_29 = _parsedindexvalue_nextIndex_T_9 & parsedindexvalue_boolArray__0; // @[Benes.scala 42:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_32 = _parsedindexvalue_nextIndex_T_29 ? _parsedindexvalue_nextIndex_T_26 : {{
    1'd0}, parsedindexvalue_first_stage}; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_33 = _parsedindexvalue_nextIndex_T_24 ? _parsedindexvalue_nextIndex_T_26 :
    _parsedindexvalue_nextIndex_T_32; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_34 = _parsedindexvalue_nextIndex_T_19 ? _parsedindexvalue_nextIndex_T_16 :
    _parsedindexvalue_nextIndex_T_33; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_35 = _parsedindexvalue_nextIndex_T_14 ? _parsedindexvalue_nextIndex_T_16 :
    _parsedindexvalue_nextIndex_T_34; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_36 = _parsedindexvalue_nextIndex_T_11 ? {{1'd0}, parsedindexvalue_first_stage
    } : _parsedindexvalue_nextIndex_T_35; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_37 = _parsedindexvalue_nextIndex_T_8 ? {{1'd0}, parsedindexvalue_first_stage}
     : _parsedindexvalue_nextIndex_T_36; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_38 = _parsedindexvalue_nextIndex_T_5 ? {{1'd0}, parsedindexvalue_first_stage}
     : _parsedindexvalue_nextIndex_T_37; // @[Mux.scala 101:16]
  wire [1:0] parsedindexvalue_nextIndex = _parsedindexvalue_nextIndex_T_2 ? {{1'd0}, parsedindexvalue_first_stage} :
    _parsedindexvalue_nextIndex_T_38; // @[Mux.scala 101:16]
  wire [2:0] _GEN_20 = {{1'd0}, parsedindexvalue_nextIndex}; // @[Benes.scala 33:40]
  wire [2:0] _GEN_25 = _GEN_20 % 3'h4; // @[Benes.scala 33:40]
  wire [1:0] parsedindexvalue_calculation_1 = _GEN_25[1:0]; // @[Benes.scala 33:40]
  wire  _parsedindexvalue_nextIndex_T_39 = parsedindexvalue_calculation_1 == 2'h0; // @[Benes.scala 35:27]
  wire  _parsedindexvalue_nextIndex_T_40 = ~parsedindexvalue_boolArray__1; // @[Benes.scala 35:53]
  wire  _parsedindexvalue_nextIndex_T_41 = parsedindexvalue_calculation_1 == 2'h0 & ~parsedindexvalue_boolArray__1; // @[Benes.scala 35:36]
  wire  _parsedindexvalue_nextIndex_T_42 = parsedindexvalue_calculation_1 == 2'h1; // @[Benes.scala 36:27]
  wire  _parsedindexvalue_nextIndex_T_44 = parsedindexvalue_calculation_1 == 2'h1 & _parsedindexvalue_nextIndex_T_40; // @[Benes.scala 36:36]
  wire  _parsedindexvalue_nextIndex_T_45 = parsedindexvalue_calculation_1 == 2'h2; // @[Benes.scala 37:27]
  wire  _parsedindexvalue_nextIndex_T_47 = parsedindexvalue_calculation_1 == 2'h2 & _parsedindexvalue_nextIndex_T_40; // @[Benes.scala 37:36]
  wire  _parsedindexvalue_nextIndex_T_48 = parsedindexvalue_calculation_1 == 2'h3; // @[Benes.scala 38:27]
  wire  _parsedindexvalue_nextIndex_T_50 = parsedindexvalue_calculation_1 == 2'h3 & _parsedindexvalue_nextIndex_T_40; // @[Benes.scala 38:36]
  wire  _parsedindexvalue_nextIndex_T_53 = _parsedindexvalue_nextIndex_T_39 & parsedindexvalue_boolArray__1; // @[Benes.scala 39:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_55 = parsedindexvalue_nextIndex + 2'h2; // @[Benes.scala 39:76]
  wire  _parsedindexvalue_nextIndex_T_58 = _parsedindexvalue_nextIndex_T_42 & parsedindexvalue_boolArray__1; // @[Benes.scala 40:36]
  wire  _parsedindexvalue_nextIndex_T_63 = _parsedindexvalue_nextIndex_T_45 & parsedindexvalue_boolArray__1; // @[Benes.scala 41:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_65 = parsedindexvalue_nextIndex - 2'h2; // @[Benes.scala 41:76]
  wire  _parsedindexvalue_nextIndex_T_68 = _parsedindexvalue_nextIndex_T_48 & parsedindexvalue_boolArray__1; // @[Benes.scala 42:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_71 = _parsedindexvalue_nextIndex_T_68 ? _parsedindexvalue_nextIndex_T_65 :
    parsedindexvalue_nextIndex; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_72 = _parsedindexvalue_nextIndex_T_63 ? _parsedindexvalue_nextIndex_T_65 :
    _parsedindexvalue_nextIndex_T_71; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_73 = _parsedindexvalue_nextIndex_T_58 ? _parsedindexvalue_nextIndex_T_55 :
    _parsedindexvalue_nextIndex_T_72; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_74 = _parsedindexvalue_nextIndex_T_53 ? _parsedindexvalue_nextIndex_T_55 :
    _parsedindexvalue_nextIndex_T_73; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_75 = _parsedindexvalue_nextIndex_T_50 ? parsedindexvalue_nextIndex :
    _parsedindexvalue_nextIndex_T_74; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_76 = _parsedindexvalue_nextIndex_T_47 ? parsedindexvalue_nextIndex :
    _parsedindexvalue_nextIndex_T_75; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_77 = _parsedindexvalue_nextIndex_T_44 ? parsedindexvalue_nextIndex :
    _parsedindexvalue_nextIndex_T_76; // @[Mux.scala 101:16]
  wire [1:0] parsedindexvalue_nextIndex_1 = _parsedindexvalue_nextIndex_T_41 ? parsedindexvalue_nextIndex :
    _parsedindexvalue_nextIndex_T_77; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_third_stage_T_1 = parsedindexvalue_nextIndex_1 % 2'h2; // @[Benes.scala 48:61]
  wire [1:0] _parsedindexvalue_third_stage_T_4 = parsedindexvalue_nextIndex_1 + 2'h1; // @[Benes.scala 48:89]
  wire [1:0] _parsedindexvalue_third_stage_T_6 = parsedindexvalue_nextIndex_1 - 2'h1; // @[Benes.scala 48:109]
  wire [1:0] _parsedindexvalue_third_stage_T_7 = _parsedindexvalue_third_stage_T_1 == 2'h0 ?
    _parsedindexvalue_third_stage_T_4 : _parsedindexvalue_third_stage_T_6; // @[Benes.scala 48:47]
  wire [1:0] parsedindexvalue = io_i_mux_bus_1[3] ? _parsedindexvalue_third_stage_T_7 : parsedindexvalue_nextIndex_1; // @[Benes.scala 48:24]
  wire [2:0] _T_3 = {{1'd0}, parsedindexvalue};
  wire [15:0] _GEN_0 = 3'h0 == _T_3 ? io_i_data_bus2_1 : 16'h0; // @[Benes.scala 63:{47,47}]
  wire [15:0] _GEN_1 = 3'h1 == _T_3 ? io_i_data_bus2_1 : 16'h0; // @[Benes.scala 63:{47,47}]
  wire [15:0] _GEN_2 = 3'h2 == _T_3 ? io_i_data_bus2_1 : 16'h0; // @[Benes.scala 63:{47,47}]
  wire [15:0] _GEN_3 = 3'h3 == _T_3 ? io_i_data_bus2_1 : 16'h0; // @[Benes.scala 63:{47,47}]
  wire  parsedindexvalue_first_stage_1 = io_i_mux_bus_1[0] ? 1'h0 : 1'h1; // @[Benes.scala 24:26]
  wire [2:0] _GEN_30 = {{2'd0}, parsedindexvalue_first_stage_1}; // @[Benes.scala 33:40]
  wire [2:0] _GEN_35 = _GEN_30 % 3'h4; // @[Benes.scala 33:40]
  wire  parsedindexvalue_calculation_2 = _GEN_35[0]; // @[Benes.scala 33:40]
  wire  _parsedindexvalue_nextIndex_T_78 = ~parsedindexvalue_calculation_2; // @[Benes.scala 35:27]
  wire  _parsedindexvalue_nextIndex_T_80 = ~parsedindexvalue_calculation_2 & ~parsedindexvalue_boolArray__0; // @[Benes.scala 35:36]
  wire  _parsedindexvalue_nextIndex_T_83 = parsedindexvalue_calculation_2 & _parsedindexvalue_nextIndex_T_1; // @[Benes.scala 36:36]
  wire [1:0] _GEN_96 = {{1'd0}, parsedindexvalue_calculation_2}; // @[Benes.scala 37:27]
  wire  _parsedindexvalue_nextIndex_T_84 = _GEN_96 == 2'h2; // @[Benes.scala 37:27]
  wire  _parsedindexvalue_nextIndex_T_86 = _GEN_96 == 2'h2 & _parsedindexvalue_nextIndex_T_1; // @[Benes.scala 37:36]
  wire  _parsedindexvalue_nextIndex_T_87 = _GEN_96 == 2'h3; // @[Benes.scala 38:27]
  wire  _parsedindexvalue_nextIndex_T_89 = _GEN_96 == 2'h3 & _parsedindexvalue_nextIndex_T_1; // @[Benes.scala 38:36]
  wire  _parsedindexvalue_nextIndex_T_92 = _parsedindexvalue_nextIndex_T_78 & parsedindexvalue_boolArray__0; // @[Benes.scala 39:36]
  wire [1:0] _GEN_98 = {{1'd0}, parsedindexvalue_first_stage_1}; // @[Benes.scala 39:76]
  wire [1:0] _parsedindexvalue_nextIndex_T_94 = _GEN_98 + 2'h2; // @[Benes.scala 39:76]
  wire  _parsedindexvalue_nextIndex_T_97 = parsedindexvalue_calculation_2 & parsedindexvalue_boolArray__0; // @[Benes.scala 40:36]
  wire  _parsedindexvalue_nextIndex_T_102 = _parsedindexvalue_nextIndex_T_84 & parsedindexvalue_boolArray__0; // @[Benes.scala 41:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_104 = _GEN_98 - 2'h2; // @[Benes.scala 41:76]
  wire  _parsedindexvalue_nextIndex_T_107 = _parsedindexvalue_nextIndex_T_87 & parsedindexvalue_boolArray__0; // @[Benes.scala 42:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_110 = _parsedindexvalue_nextIndex_T_107 ? _parsedindexvalue_nextIndex_T_104
     : {{1'd0}, parsedindexvalue_first_stage_1}; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_111 = _parsedindexvalue_nextIndex_T_102 ? _parsedindexvalue_nextIndex_T_104
     : _parsedindexvalue_nextIndex_T_110; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_112 = _parsedindexvalue_nextIndex_T_97 ? _parsedindexvalue_nextIndex_T_94 :
    _parsedindexvalue_nextIndex_T_111; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_113 = _parsedindexvalue_nextIndex_T_92 ? _parsedindexvalue_nextIndex_T_94 :
    _parsedindexvalue_nextIndex_T_112; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_114 = _parsedindexvalue_nextIndex_T_89 ? {{1'd0},
    parsedindexvalue_first_stage_1} : _parsedindexvalue_nextIndex_T_113; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_115 = _parsedindexvalue_nextIndex_T_86 ? {{1'd0},
    parsedindexvalue_first_stage_1} : _parsedindexvalue_nextIndex_T_114; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_116 = _parsedindexvalue_nextIndex_T_83 ? {{1'd0},
    parsedindexvalue_first_stage_1} : _parsedindexvalue_nextIndex_T_115; // @[Mux.scala 101:16]
  wire [1:0] parsedindexvalue_nextIndex_2 = _parsedindexvalue_nextIndex_T_80 ? {{1'd0}, parsedindexvalue_first_stage_1}
     : _parsedindexvalue_nextIndex_T_116; // @[Mux.scala 101:16]
  wire [2:0] _GEN_40 = {{1'd0}, parsedindexvalue_nextIndex_2}; // @[Benes.scala 33:40]
  wire [2:0] _GEN_46 = _GEN_40 % 3'h4; // @[Benes.scala 33:40]
  wire [1:0] parsedindexvalue_calculation_3 = _GEN_46[1:0]; // @[Benes.scala 33:40]
  wire  _parsedindexvalue_nextIndex_T_117 = parsedindexvalue_calculation_3 == 2'h0; // @[Benes.scala 35:27]
  wire  _parsedindexvalue_nextIndex_T_119 = parsedindexvalue_calculation_3 == 2'h0 & ~parsedindexvalue_boolArray__1; // @[Benes.scala 35:36]
  wire  _parsedindexvalue_nextIndex_T_120 = parsedindexvalue_calculation_3 == 2'h1; // @[Benes.scala 36:27]
  wire  _parsedindexvalue_nextIndex_T_122 = parsedindexvalue_calculation_3 == 2'h1 & _parsedindexvalue_nextIndex_T_40; // @[Benes.scala 36:36]
  wire  _parsedindexvalue_nextIndex_T_123 = parsedindexvalue_calculation_3 == 2'h2; // @[Benes.scala 37:27]
  wire  _parsedindexvalue_nextIndex_T_125 = parsedindexvalue_calculation_3 == 2'h2 & _parsedindexvalue_nextIndex_T_40; // @[Benes.scala 37:36]
  wire  _parsedindexvalue_nextIndex_T_126 = parsedindexvalue_calculation_3 == 2'h3; // @[Benes.scala 38:27]
  wire  _parsedindexvalue_nextIndex_T_128 = parsedindexvalue_calculation_3 == 2'h3 & _parsedindexvalue_nextIndex_T_40; // @[Benes.scala 38:36]
  wire  _parsedindexvalue_nextIndex_T_131 = _parsedindexvalue_nextIndex_T_117 & parsedindexvalue_boolArray__1; // @[Benes.scala 39:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_133 = parsedindexvalue_nextIndex_2 + 2'h2; // @[Benes.scala 39:76]
  wire  _parsedindexvalue_nextIndex_T_136 = _parsedindexvalue_nextIndex_T_120 & parsedindexvalue_boolArray__1; // @[Benes.scala 40:36]
  wire  _parsedindexvalue_nextIndex_T_141 = _parsedindexvalue_nextIndex_T_123 & parsedindexvalue_boolArray__1; // @[Benes.scala 41:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_143 = parsedindexvalue_nextIndex_2 - 2'h2; // @[Benes.scala 41:76]
  wire  _parsedindexvalue_nextIndex_T_146 = _parsedindexvalue_nextIndex_T_126 & parsedindexvalue_boolArray__1; // @[Benes.scala 42:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_149 = _parsedindexvalue_nextIndex_T_146 ? _parsedindexvalue_nextIndex_T_143
     : parsedindexvalue_nextIndex_2; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_150 = _parsedindexvalue_nextIndex_T_141 ? _parsedindexvalue_nextIndex_T_143
     : _parsedindexvalue_nextIndex_T_149; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_151 = _parsedindexvalue_nextIndex_T_136 ? _parsedindexvalue_nextIndex_T_133
     : _parsedindexvalue_nextIndex_T_150; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_152 = _parsedindexvalue_nextIndex_T_131 ? _parsedindexvalue_nextIndex_T_133
     : _parsedindexvalue_nextIndex_T_151; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_153 = _parsedindexvalue_nextIndex_T_128 ? parsedindexvalue_nextIndex_2 :
    _parsedindexvalue_nextIndex_T_152; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_154 = _parsedindexvalue_nextIndex_T_125 ? parsedindexvalue_nextIndex_2 :
    _parsedindexvalue_nextIndex_T_153; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_155 = _parsedindexvalue_nextIndex_T_122 ? parsedindexvalue_nextIndex_2 :
    _parsedindexvalue_nextIndex_T_154; // @[Mux.scala 101:16]
  wire [1:0] parsedindexvalue_nextIndex_3 = _parsedindexvalue_nextIndex_T_119 ? parsedindexvalue_nextIndex_2 :
    _parsedindexvalue_nextIndex_T_155; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_third_stage_T_9 = parsedindexvalue_nextIndex_3 % 2'h2; // @[Benes.scala 48:61]
  wire [1:0] _parsedindexvalue_third_stage_T_12 = parsedindexvalue_nextIndex_3 + 2'h1; // @[Benes.scala 48:89]
  wire [1:0] _parsedindexvalue_third_stage_T_14 = parsedindexvalue_nextIndex_3 - 2'h1; // @[Benes.scala 48:109]
  wire [1:0] _parsedindexvalue_third_stage_T_15 = _parsedindexvalue_third_stage_T_9 == 2'h0 ?
    _parsedindexvalue_third_stage_T_12 : _parsedindexvalue_third_stage_T_14; // @[Benes.scala 48:47]
  wire [1:0] parsedindexvalue_1 = io_i_mux_bus_1[3] ? _parsedindexvalue_third_stage_T_15 : parsedindexvalue_nextIndex_3; // @[Benes.scala 48:24]
  wire [2:0] _T_5 = {{1'd0}, parsedindexvalue_1};
  wire [15:0] _GEN_5 = 3'h0 == _T_5 ? io_i_data_bus2_1 : 16'h0; // @[Benes.scala 67:{47,47}]
  wire [15:0] _GEN_6 = 3'h1 == _T_5 ? io_i_data_bus2_1 : 16'h0; // @[Benes.scala 67:{47,47}]
  wire [15:0] _GEN_7 = 3'h2 == _T_5 ? io_i_data_bus2_1 : 16'h0; // @[Benes.scala 67:{47,47}]
  wire [15:0] _GEN_8 = 3'h3 == _T_5 ? io_i_data_bus2_1 : 16'h0; // @[Benes.scala 67:{47,47}]
  wire [15:0] _GEN_10 = io_i_data_bus2_1 == io_i_data_bus2_0 ? _GEN_0 : _GEN_5; // @[Benes.scala 60:61]
  wire [15:0] _GEN_11 = io_i_data_bus2_1 == io_i_data_bus2_0 ? _GEN_1 : _GEN_6; // @[Benes.scala 60:61]
  wire [15:0] _GEN_12 = io_i_data_bus2_1 == io_i_data_bus2_0 ? _GEN_2 : _GEN_7; // @[Benes.scala 60:61]
  wire [15:0] _GEN_13 = io_i_data_bus2_1 == io_i_data_bus2_0 ? _GEN_3 : _GEN_8; // @[Benes.scala 60:61]
  wire [15:0] _GEN_15 = _T_2 ? 16'h0 : io_i_data_bus2_1; // @[Benes.scala 72:60 74:28 78:28]
  wire [15:0] _GEN_16 = |io_i_mux_bus_1 ? _GEN_10 : 16'h0; // @[Benes.scala 58:35]
  wire [15:0] _GEN_17 = |io_i_mux_bus_1 ? _GEN_11 : _GEN_15; // @[Benes.scala 58:35]
  wire [15:0] _GEN_18 = |io_i_mux_bus_1 ? _GEN_12 : 16'h0; // @[Benes.scala 58:35]
  wire [15:0] _GEN_19 = |io_i_mux_bus_1 ? _GEN_13 : 16'h0; // @[Benes.scala 58:35]
  wire [15:0] _GEN_21 = io_i_data_bus2_1 != 16'h0 ? _GEN_16 : 16'h0; // @[Benes.scala 56:39]
  wire [15:0] _GEN_22 = io_i_data_bus2_1 != 16'h0 ? _GEN_17 : 16'h0; // @[Benes.scala 56:39]
  wire [15:0] _GEN_23 = io_i_data_bus2_1 != 16'h0 ? _GEN_18 : 16'h0; // @[Benes.scala 56:39]
  wire [15:0] _GEN_24 = io_i_data_bus2_1 != 16'h0 ? _GEN_19 : 16'h0; // @[Benes.scala 56:39]
  wire  _T_10 = io_i_data_bus2_2 == io_i_data_bus2_1; // @[Benes.scala 60:36]
  wire [1:0] _parsedindexvalue_T_5 = 2'h2 - 2'h1; // @[Benes.scala 62:97]
  wire [1:0] _parsedindexvalue_first_stage_T_17 = _parsedindexvalue_T_5 % 2'h2; // @[Benes.scala 24:52]
  wire [1:0] _parsedindexvalue_first_stage_T_20 = _parsedindexvalue_T_5 + 2'h1; // @[Benes.scala 24:78]
  wire [1:0] _parsedindexvalue_first_stage_T_22 = _parsedindexvalue_T_5 - 2'h1; // @[Benes.scala 24:96]
  wire [1:0] _parsedindexvalue_first_stage_T_23 = _parsedindexvalue_first_stage_T_17 == 2'h0 ?
    _parsedindexvalue_first_stage_T_20 : _parsedindexvalue_first_stage_T_22; // @[Benes.scala 24:40]
  wire [1:0] parsedindexvalue_first_stage_2 = io_i_mux_bus_2[0] ? _parsedindexvalue_first_stage_T_23 :
    _parsedindexvalue_T_5; // @[Benes.scala 24:26]
  wire  parsedindexvalue_boolArray_2_0 = io_i_mux_bus_2[1]; // @[Benes.scala 28:92]
  wire  parsedindexvalue_boolArray_2_1 = io_i_mux_bus_2[2]; // @[Benes.scala 28:92]
  wire [2:0] _GEN_51 = {{1'd0}, parsedindexvalue_first_stage_2}; // @[Benes.scala 33:40]
  wire [2:0] _GEN_56 = _GEN_51 % 3'h4; // @[Benes.scala 33:40]
  wire [1:0] parsedindexvalue_calculation_4 = _GEN_56[1:0]; // @[Benes.scala 33:40]
  wire  _parsedindexvalue_nextIndex_T_156 = parsedindexvalue_calculation_4 == 2'h0; // @[Benes.scala 35:27]
  wire  _parsedindexvalue_nextIndex_T_157 = ~parsedindexvalue_boolArray_2_0; // @[Benes.scala 35:53]
  wire  _parsedindexvalue_nextIndex_T_158 = parsedindexvalue_calculation_4 == 2'h0 & ~parsedindexvalue_boolArray_2_0; // @[Benes.scala 35:36]
  wire  _parsedindexvalue_nextIndex_T_159 = parsedindexvalue_calculation_4 == 2'h1; // @[Benes.scala 36:27]
  wire  _parsedindexvalue_nextIndex_T_161 = parsedindexvalue_calculation_4 == 2'h1 & _parsedindexvalue_nextIndex_T_157; // @[Benes.scala 36:36]
  wire  _parsedindexvalue_nextIndex_T_162 = parsedindexvalue_calculation_4 == 2'h2; // @[Benes.scala 37:27]
  wire  _parsedindexvalue_nextIndex_T_164 = parsedindexvalue_calculation_4 == 2'h2 & _parsedindexvalue_nextIndex_T_157; // @[Benes.scala 37:36]
  wire  _parsedindexvalue_nextIndex_T_165 = parsedindexvalue_calculation_4 == 2'h3; // @[Benes.scala 38:27]
  wire  _parsedindexvalue_nextIndex_T_167 = parsedindexvalue_calculation_4 == 2'h3 & _parsedindexvalue_nextIndex_T_157; // @[Benes.scala 38:36]
  wire  _parsedindexvalue_nextIndex_T_170 = _parsedindexvalue_nextIndex_T_156 & parsedindexvalue_boolArray_2_0; // @[Benes.scala 39:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_172 = parsedindexvalue_first_stage_2 + 2'h2; // @[Benes.scala 39:76]
  wire  _parsedindexvalue_nextIndex_T_175 = _parsedindexvalue_nextIndex_T_159 & parsedindexvalue_boolArray_2_0; // @[Benes.scala 40:36]
  wire  _parsedindexvalue_nextIndex_T_180 = _parsedindexvalue_nextIndex_T_162 & parsedindexvalue_boolArray_2_0; // @[Benes.scala 41:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_182 = parsedindexvalue_first_stage_2 - 2'h2; // @[Benes.scala 41:76]
  wire  _parsedindexvalue_nextIndex_T_185 = _parsedindexvalue_nextIndex_T_165 & parsedindexvalue_boolArray_2_0; // @[Benes.scala 42:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_188 = _parsedindexvalue_nextIndex_T_185 ? _parsedindexvalue_nextIndex_T_182
     : parsedindexvalue_first_stage_2; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_189 = _parsedindexvalue_nextIndex_T_180 ? _parsedindexvalue_nextIndex_T_182
     : _parsedindexvalue_nextIndex_T_188; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_190 = _parsedindexvalue_nextIndex_T_175 ? _parsedindexvalue_nextIndex_T_172
     : _parsedindexvalue_nextIndex_T_189; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_191 = _parsedindexvalue_nextIndex_T_170 ? _parsedindexvalue_nextIndex_T_172
     : _parsedindexvalue_nextIndex_T_190; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_192 = _parsedindexvalue_nextIndex_T_167 ? parsedindexvalue_first_stage_2 :
    _parsedindexvalue_nextIndex_T_191; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_193 = _parsedindexvalue_nextIndex_T_164 ? parsedindexvalue_first_stage_2 :
    _parsedindexvalue_nextIndex_T_192; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_194 = _parsedindexvalue_nextIndex_T_161 ? parsedindexvalue_first_stage_2 :
    _parsedindexvalue_nextIndex_T_193; // @[Mux.scala 101:16]
  wire [1:0] parsedindexvalue_nextIndex_4 = _parsedindexvalue_nextIndex_T_158 ? parsedindexvalue_first_stage_2 :
    _parsedindexvalue_nextIndex_T_194; // @[Mux.scala 101:16]
  wire [2:0] _GEN_61 = {{1'd0}, parsedindexvalue_nextIndex_4}; // @[Benes.scala 33:40]
  wire [2:0] _GEN_66 = _GEN_61 % 3'h4; // @[Benes.scala 33:40]
  wire [1:0] parsedindexvalue_calculation_5 = _GEN_66[1:0]; // @[Benes.scala 33:40]
  wire  _parsedindexvalue_nextIndex_T_195 = parsedindexvalue_calculation_5 == 2'h0; // @[Benes.scala 35:27]
  wire  _parsedindexvalue_nextIndex_T_196 = ~parsedindexvalue_boolArray_2_1; // @[Benes.scala 35:53]
  wire  _parsedindexvalue_nextIndex_T_197 = parsedindexvalue_calculation_5 == 2'h0 & ~parsedindexvalue_boolArray_2_1; // @[Benes.scala 35:36]
  wire  _parsedindexvalue_nextIndex_T_198 = parsedindexvalue_calculation_5 == 2'h1; // @[Benes.scala 36:27]
  wire  _parsedindexvalue_nextIndex_T_200 = parsedindexvalue_calculation_5 == 2'h1 & _parsedindexvalue_nextIndex_T_196; // @[Benes.scala 36:36]
  wire  _parsedindexvalue_nextIndex_T_201 = parsedindexvalue_calculation_5 == 2'h2; // @[Benes.scala 37:27]
  wire  _parsedindexvalue_nextIndex_T_203 = parsedindexvalue_calculation_5 == 2'h2 & _parsedindexvalue_nextIndex_T_196; // @[Benes.scala 37:36]
  wire  _parsedindexvalue_nextIndex_T_204 = parsedindexvalue_calculation_5 == 2'h3; // @[Benes.scala 38:27]
  wire  _parsedindexvalue_nextIndex_T_206 = parsedindexvalue_calculation_5 == 2'h3 & _parsedindexvalue_nextIndex_T_196; // @[Benes.scala 38:36]
  wire  _parsedindexvalue_nextIndex_T_209 = _parsedindexvalue_nextIndex_T_195 & parsedindexvalue_boolArray_2_1; // @[Benes.scala 39:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_211 = parsedindexvalue_nextIndex_4 + 2'h2; // @[Benes.scala 39:76]
  wire  _parsedindexvalue_nextIndex_T_214 = _parsedindexvalue_nextIndex_T_198 & parsedindexvalue_boolArray_2_1; // @[Benes.scala 40:36]
  wire  _parsedindexvalue_nextIndex_T_219 = _parsedindexvalue_nextIndex_T_201 & parsedindexvalue_boolArray_2_1; // @[Benes.scala 41:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_221 = parsedindexvalue_nextIndex_4 - 2'h2; // @[Benes.scala 41:76]
  wire  _parsedindexvalue_nextIndex_T_224 = _parsedindexvalue_nextIndex_T_204 & parsedindexvalue_boolArray_2_1; // @[Benes.scala 42:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_227 = _parsedindexvalue_nextIndex_T_224 ? _parsedindexvalue_nextIndex_T_221
     : parsedindexvalue_nextIndex_4; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_228 = _parsedindexvalue_nextIndex_T_219 ? _parsedindexvalue_nextIndex_T_221
     : _parsedindexvalue_nextIndex_T_227; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_229 = _parsedindexvalue_nextIndex_T_214 ? _parsedindexvalue_nextIndex_T_211
     : _parsedindexvalue_nextIndex_T_228; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_230 = _parsedindexvalue_nextIndex_T_209 ? _parsedindexvalue_nextIndex_T_211
     : _parsedindexvalue_nextIndex_T_229; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_231 = _parsedindexvalue_nextIndex_T_206 ? parsedindexvalue_nextIndex_4 :
    _parsedindexvalue_nextIndex_T_230; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_232 = _parsedindexvalue_nextIndex_T_203 ? parsedindexvalue_nextIndex_4 :
    _parsedindexvalue_nextIndex_T_231; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_233 = _parsedindexvalue_nextIndex_T_200 ? parsedindexvalue_nextIndex_4 :
    _parsedindexvalue_nextIndex_T_232; // @[Mux.scala 101:16]
  wire [1:0] parsedindexvalue_nextIndex_5 = _parsedindexvalue_nextIndex_T_197 ? parsedindexvalue_nextIndex_4 :
    _parsedindexvalue_nextIndex_T_233; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_third_stage_T_17 = parsedindexvalue_nextIndex_5 % 2'h2; // @[Benes.scala 48:61]
  wire [1:0] _parsedindexvalue_third_stage_T_20 = parsedindexvalue_nextIndex_5 + 2'h1; // @[Benes.scala 48:89]
  wire [1:0] _parsedindexvalue_third_stage_T_22 = parsedindexvalue_nextIndex_5 - 2'h1; // @[Benes.scala 48:109]
  wire [1:0] _parsedindexvalue_third_stage_T_23 = _parsedindexvalue_third_stage_T_17 == 2'h0 ?
    _parsedindexvalue_third_stage_T_20 : _parsedindexvalue_third_stage_T_22; // @[Benes.scala 48:47]
  wire [1:0] parsedindexvalue_2 = io_i_mux_bus_2[3] ? _parsedindexvalue_third_stage_T_23 : parsedindexvalue_nextIndex_5; // @[Benes.scala 48:24]
  wire [2:0] _T_11 = {{1'd0}, parsedindexvalue_2};
  wire [15:0] _GEN_26 = 3'h0 == _T_11 ? io_i_data_bus2_2 : _GEN_21; // @[Benes.scala 63:{47,47}]
  wire [15:0] _GEN_27 = 3'h1 == _T_11 ? io_i_data_bus2_2 : _GEN_22; // @[Benes.scala 63:{47,47}]
  wire [15:0] _GEN_28 = 3'h2 == _T_11 ? io_i_data_bus2_2 : _GEN_23; // @[Benes.scala 63:{47,47}]
  wire [15:0] _GEN_29 = 3'h3 == _T_11 ? io_i_data_bus2_2 : _GEN_24; // @[Benes.scala 63:{47,47}]
  wire [1:0] parsedindexvalue_first_stage_3 = io_i_mux_bus_2[0] ? 2'h3 : 2'h2; // @[Benes.scala 24:26]
  wire [2:0] _GEN_72 = {{1'd0}, parsedindexvalue_first_stage_3}; // @[Benes.scala 33:40]
  wire [2:0] _GEN_77 = _GEN_72 % 3'h4; // @[Benes.scala 33:40]
  wire [1:0] parsedindexvalue_calculation_6 = _GEN_77[1:0]; // @[Benes.scala 33:40]
  wire  _parsedindexvalue_nextIndex_T_234 = parsedindexvalue_calculation_6 == 2'h0; // @[Benes.scala 35:27]
  wire  _parsedindexvalue_nextIndex_T_236 = parsedindexvalue_calculation_6 == 2'h0 & ~parsedindexvalue_boolArray_2_0; // @[Benes.scala 35:36]
  wire  _parsedindexvalue_nextIndex_T_237 = parsedindexvalue_calculation_6 == 2'h1; // @[Benes.scala 36:27]
  wire  _parsedindexvalue_nextIndex_T_239 = parsedindexvalue_calculation_6 == 2'h1 & _parsedindexvalue_nextIndex_T_157; // @[Benes.scala 36:36]
  wire  _parsedindexvalue_nextIndex_T_240 = parsedindexvalue_calculation_6 == 2'h2; // @[Benes.scala 37:27]
  wire  _parsedindexvalue_nextIndex_T_242 = parsedindexvalue_calculation_6 == 2'h2 & _parsedindexvalue_nextIndex_T_157; // @[Benes.scala 37:36]
  wire  _parsedindexvalue_nextIndex_T_243 = parsedindexvalue_calculation_6 == 2'h3; // @[Benes.scala 38:27]
  wire  _parsedindexvalue_nextIndex_T_245 = parsedindexvalue_calculation_6 == 2'h3 & _parsedindexvalue_nextIndex_T_157; // @[Benes.scala 38:36]
  wire  _parsedindexvalue_nextIndex_T_248 = _parsedindexvalue_nextIndex_T_234 & parsedindexvalue_boolArray_2_0; // @[Benes.scala 39:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_250 = parsedindexvalue_first_stage_3 + 2'h2; // @[Benes.scala 39:76]
  wire  _parsedindexvalue_nextIndex_T_253 = _parsedindexvalue_nextIndex_T_237 & parsedindexvalue_boolArray_2_0; // @[Benes.scala 40:36]
  wire  _parsedindexvalue_nextIndex_T_258 = _parsedindexvalue_nextIndex_T_240 & parsedindexvalue_boolArray_2_0; // @[Benes.scala 41:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_260 = parsedindexvalue_first_stage_3 - 2'h2; // @[Benes.scala 41:76]
  wire  _parsedindexvalue_nextIndex_T_263 = _parsedindexvalue_nextIndex_T_243 & parsedindexvalue_boolArray_2_0; // @[Benes.scala 42:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_266 = _parsedindexvalue_nextIndex_T_263 ? _parsedindexvalue_nextIndex_T_260
     : parsedindexvalue_first_stage_3; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_267 = _parsedindexvalue_nextIndex_T_258 ? _parsedindexvalue_nextIndex_T_260
     : _parsedindexvalue_nextIndex_T_266; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_268 = _parsedindexvalue_nextIndex_T_253 ? _parsedindexvalue_nextIndex_T_250
     : _parsedindexvalue_nextIndex_T_267; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_269 = _parsedindexvalue_nextIndex_T_248 ? _parsedindexvalue_nextIndex_T_250
     : _parsedindexvalue_nextIndex_T_268; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_270 = _parsedindexvalue_nextIndex_T_245 ? parsedindexvalue_first_stage_3 :
    _parsedindexvalue_nextIndex_T_269; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_271 = _parsedindexvalue_nextIndex_T_242 ? parsedindexvalue_first_stage_3 :
    _parsedindexvalue_nextIndex_T_270; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_272 = _parsedindexvalue_nextIndex_T_239 ? parsedindexvalue_first_stage_3 :
    _parsedindexvalue_nextIndex_T_271; // @[Mux.scala 101:16]
  wire [1:0] parsedindexvalue_nextIndex_6 = _parsedindexvalue_nextIndex_T_236 ? parsedindexvalue_first_stage_3 :
    _parsedindexvalue_nextIndex_T_272; // @[Mux.scala 101:16]
  wire [2:0] _GEN_82 = {{1'd0}, parsedindexvalue_nextIndex_6}; // @[Benes.scala 33:40]
  wire [2:0] _GEN_83 = _GEN_82 % 3'h4; // @[Benes.scala 33:40]
  wire [1:0] parsedindexvalue_calculation_7 = _GEN_83[1:0]; // @[Benes.scala 33:40]
  wire  _parsedindexvalue_nextIndex_T_273 = parsedindexvalue_calculation_7 == 2'h0; // @[Benes.scala 35:27]
  wire  _parsedindexvalue_nextIndex_T_275 = parsedindexvalue_calculation_7 == 2'h0 & ~parsedindexvalue_boolArray_2_1; // @[Benes.scala 35:36]
  wire  _parsedindexvalue_nextIndex_T_276 = parsedindexvalue_calculation_7 == 2'h1; // @[Benes.scala 36:27]
  wire  _parsedindexvalue_nextIndex_T_278 = parsedindexvalue_calculation_7 == 2'h1 & _parsedindexvalue_nextIndex_T_196; // @[Benes.scala 36:36]
  wire  _parsedindexvalue_nextIndex_T_279 = parsedindexvalue_calculation_7 == 2'h2; // @[Benes.scala 37:27]
  wire  _parsedindexvalue_nextIndex_T_281 = parsedindexvalue_calculation_7 == 2'h2 & _parsedindexvalue_nextIndex_T_196; // @[Benes.scala 37:36]
  wire  _parsedindexvalue_nextIndex_T_282 = parsedindexvalue_calculation_7 == 2'h3; // @[Benes.scala 38:27]
  wire  _parsedindexvalue_nextIndex_T_284 = parsedindexvalue_calculation_7 == 2'h3 & _parsedindexvalue_nextIndex_T_196; // @[Benes.scala 38:36]
  wire  _parsedindexvalue_nextIndex_T_287 = _parsedindexvalue_nextIndex_T_273 & parsedindexvalue_boolArray_2_1; // @[Benes.scala 39:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_289 = parsedindexvalue_nextIndex_6 + 2'h2; // @[Benes.scala 39:76]
  wire  _parsedindexvalue_nextIndex_T_292 = _parsedindexvalue_nextIndex_T_276 & parsedindexvalue_boolArray_2_1; // @[Benes.scala 40:36]
  wire  _parsedindexvalue_nextIndex_T_297 = _parsedindexvalue_nextIndex_T_279 & parsedindexvalue_boolArray_2_1; // @[Benes.scala 41:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_299 = parsedindexvalue_nextIndex_6 - 2'h2; // @[Benes.scala 41:76]
  wire  _parsedindexvalue_nextIndex_T_302 = _parsedindexvalue_nextIndex_T_282 & parsedindexvalue_boolArray_2_1; // @[Benes.scala 42:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_305 = _parsedindexvalue_nextIndex_T_302 ? _parsedindexvalue_nextIndex_T_299
     : parsedindexvalue_nextIndex_6; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_306 = _parsedindexvalue_nextIndex_T_297 ? _parsedindexvalue_nextIndex_T_299
     : _parsedindexvalue_nextIndex_T_305; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_307 = _parsedindexvalue_nextIndex_T_292 ? _parsedindexvalue_nextIndex_T_289
     : _parsedindexvalue_nextIndex_T_306; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_308 = _parsedindexvalue_nextIndex_T_287 ? _parsedindexvalue_nextIndex_T_289
     : _parsedindexvalue_nextIndex_T_307; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_309 = _parsedindexvalue_nextIndex_T_284 ? parsedindexvalue_nextIndex_6 :
    _parsedindexvalue_nextIndex_T_308; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_310 = _parsedindexvalue_nextIndex_T_281 ? parsedindexvalue_nextIndex_6 :
    _parsedindexvalue_nextIndex_T_309; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_311 = _parsedindexvalue_nextIndex_T_278 ? parsedindexvalue_nextIndex_6 :
    _parsedindexvalue_nextIndex_T_310; // @[Mux.scala 101:16]
  wire [1:0] parsedindexvalue_nextIndex_7 = _parsedindexvalue_nextIndex_T_275 ? parsedindexvalue_nextIndex_6 :
    _parsedindexvalue_nextIndex_T_311; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_third_stage_T_25 = parsedindexvalue_nextIndex_7 % 2'h2; // @[Benes.scala 48:61]
  wire [1:0] _parsedindexvalue_third_stage_T_28 = parsedindexvalue_nextIndex_7 + 2'h1; // @[Benes.scala 48:89]
  wire [1:0] _parsedindexvalue_third_stage_T_30 = parsedindexvalue_nextIndex_7 - 2'h1; // @[Benes.scala 48:109]
  wire [1:0] _parsedindexvalue_third_stage_T_31 = _parsedindexvalue_third_stage_T_25 == 2'h0 ?
    _parsedindexvalue_third_stage_T_28 : _parsedindexvalue_third_stage_T_30; // @[Benes.scala 48:47]
  wire [1:0] parsedindexvalue_3 = io_i_mux_bus_2[3] ? _parsedindexvalue_third_stage_T_31 : parsedindexvalue_nextIndex_7; // @[Benes.scala 48:24]
  wire [2:0] _T_13 = {{1'd0}, parsedindexvalue_3};
  wire [15:0] _GEN_31 = 3'h0 == _T_13 ? io_i_data_bus2_2 : _GEN_21; // @[Benes.scala 67:{47,47}]
  wire [15:0] _GEN_32 = 3'h1 == _T_13 ? io_i_data_bus2_2 : _GEN_22; // @[Benes.scala 67:{47,47}]
  wire [15:0] _GEN_33 = 3'h2 == _T_13 ? io_i_data_bus2_2 : _GEN_23; // @[Benes.scala 67:{47,47}]
  wire [15:0] _GEN_34 = 3'h3 == _T_13 ? io_i_data_bus2_2 : _GEN_24; // @[Benes.scala 67:{47,47}]
  wire [15:0] _GEN_36 = io_i_data_bus2_2 == io_i_data_bus2_1 ? _GEN_26 : _GEN_31; // @[Benes.scala 60:61]
  wire [15:0] _GEN_37 = io_i_data_bus2_2 == io_i_data_bus2_1 ? _GEN_27 : _GEN_32; // @[Benes.scala 60:61]
  wire [15:0] _GEN_38 = io_i_data_bus2_2 == io_i_data_bus2_1 ? _GEN_28 : _GEN_33; // @[Benes.scala 60:61]
  wire [15:0] _GEN_39 = io_i_data_bus2_2 == io_i_data_bus2_1 ? _GEN_29 : _GEN_34; // @[Benes.scala 60:61]
  wire [15:0] _GEN_41 = _T_10 ? 16'h0 : io_i_data_bus2_2; // @[Benes.scala 72:60 74:28 78:28]
  wire [15:0] _GEN_42 = |io_i_mux_bus_2 ? _GEN_36 : _GEN_21; // @[Benes.scala 58:35]
  wire [15:0] _GEN_43 = |io_i_mux_bus_2 ? _GEN_37 : _GEN_22; // @[Benes.scala 58:35]
  wire [15:0] _GEN_44 = |io_i_mux_bus_2 ? _GEN_38 : _GEN_41; // @[Benes.scala 58:35]
  wire [15:0] _GEN_45 = |io_i_mux_bus_2 ? _GEN_39 : _GEN_24; // @[Benes.scala 58:35]
  wire [15:0] _GEN_47 = io_i_data_bus2_2 != 16'h0 ? _GEN_42 : _GEN_21; // @[Benes.scala 56:39]
  wire [15:0] _GEN_48 = io_i_data_bus2_2 != 16'h0 ? _GEN_43 : _GEN_22; // @[Benes.scala 56:39]
  wire [15:0] _GEN_49 = io_i_data_bus2_2 != 16'h0 ? _GEN_44 : _GEN_23; // @[Benes.scala 56:39]
  wire [15:0] _GEN_50 = io_i_data_bus2_2 != 16'h0 ? _GEN_45 : _GEN_24; // @[Benes.scala 56:39]
  wire  _T_18 = io_i_data_bus2_3 == io_i_data_bus2_2; // @[Benes.scala 60:36]
  wire [1:0] _parsedindexvalue_T_9 = 2'h3 - 2'h1; // @[Benes.scala 62:97]
  wire [1:0] _parsedindexvalue_first_stage_T_33 = _parsedindexvalue_T_9 % 2'h2; // @[Benes.scala 24:52]
  wire [1:0] _parsedindexvalue_first_stage_T_36 = _parsedindexvalue_T_9 + 2'h1; // @[Benes.scala 24:78]
  wire [1:0] _parsedindexvalue_first_stage_T_38 = _parsedindexvalue_T_9 - 2'h1; // @[Benes.scala 24:96]
  wire [1:0] _parsedindexvalue_first_stage_T_39 = _parsedindexvalue_first_stage_T_33 == 2'h0 ?
    _parsedindexvalue_first_stage_T_36 : _parsedindexvalue_first_stage_T_38; // @[Benes.scala 24:40]
  wire [1:0] parsedindexvalue_first_stage_4 = io_i_mux_bus_3[0] ? _parsedindexvalue_first_stage_T_39 :
    _parsedindexvalue_T_9; // @[Benes.scala 24:26]
  wire  parsedindexvalue_boolArray_4_0 = io_i_mux_bus_3[1]; // @[Benes.scala 28:92]
  wire  parsedindexvalue_boolArray_4_1 = io_i_mux_bus_3[2]; // @[Benes.scala 28:92]
  wire [2:0] _GEN_84 = {{1'd0}, parsedindexvalue_first_stage_4}; // @[Benes.scala 33:40]
  wire [2:0] _GEN_85 = _GEN_84 % 3'h4; // @[Benes.scala 33:40]
  wire [1:0] parsedindexvalue_calculation_8 = _GEN_85[1:0]; // @[Benes.scala 33:40]
  wire  _parsedindexvalue_nextIndex_T_312 = parsedindexvalue_calculation_8 == 2'h0; // @[Benes.scala 35:27]
  wire  _parsedindexvalue_nextIndex_T_313 = ~parsedindexvalue_boolArray_4_0; // @[Benes.scala 35:53]
  wire  _parsedindexvalue_nextIndex_T_314 = parsedindexvalue_calculation_8 == 2'h0 & ~parsedindexvalue_boolArray_4_0; // @[Benes.scala 35:36]
  wire  _parsedindexvalue_nextIndex_T_315 = parsedindexvalue_calculation_8 == 2'h1; // @[Benes.scala 36:27]
  wire  _parsedindexvalue_nextIndex_T_317 = parsedindexvalue_calculation_8 == 2'h1 & _parsedindexvalue_nextIndex_T_313; // @[Benes.scala 36:36]
  wire  _parsedindexvalue_nextIndex_T_318 = parsedindexvalue_calculation_8 == 2'h2; // @[Benes.scala 37:27]
  wire  _parsedindexvalue_nextIndex_T_320 = parsedindexvalue_calculation_8 == 2'h2 & _parsedindexvalue_nextIndex_T_313; // @[Benes.scala 37:36]
  wire  _parsedindexvalue_nextIndex_T_321 = parsedindexvalue_calculation_8 == 2'h3; // @[Benes.scala 38:27]
  wire  _parsedindexvalue_nextIndex_T_323 = parsedindexvalue_calculation_8 == 2'h3 & _parsedindexvalue_nextIndex_T_313; // @[Benes.scala 38:36]
  wire  _parsedindexvalue_nextIndex_T_326 = _parsedindexvalue_nextIndex_T_312 & parsedindexvalue_boolArray_4_0; // @[Benes.scala 39:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_328 = parsedindexvalue_first_stage_4 + 2'h2; // @[Benes.scala 39:76]
  wire  _parsedindexvalue_nextIndex_T_331 = _parsedindexvalue_nextIndex_T_315 & parsedindexvalue_boolArray_4_0; // @[Benes.scala 40:36]
  wire  _parsedindexvalue_nextIndex_T_336 = _parsedindexvalue_nextIndex_T_318 & parsedindexvalue_boolArray_4_0; // @[Benes.scala 41:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_338 = parsedindexvalue_first_stage_4 - 2'h2; // @[Benes.scala 41:76]
  wire  _parsedindexvalue_nextIndex_T_341 = _parsedindexvalue_nextIndex_T_321 & parsedindexvalue_boolArray_4_0; // @[Benes.scala 42:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_344 = _parsedindexvalue_nextIndex_T_341 ? _parsedindexvalue_nextIndex_T_338
     : parsedindexvalue_first_stage_4; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_345 = _parsedindexvalue_nextIndex_T_336 ? _parsedindexvalue_nextIndex_T_338
     : _parsedindexvalue_nextIndex_T_344; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_346 = _parsedindexvalue_nextIndex_T_331 ? _parsedindexvalue_nextIndex_T_328
     : _parsedindexvalue_nextIndex_T_345; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_347 = _parsedindexvalue_nextIndex_T_326 ? _parsedindexvalue_nextIndex_T_328
     : _parsedindexvalue_nextIndex_T_346; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_348 = _parsedindexvalue_nextIndex_T_323 ? parsedindexvalue_first_stage_4 :
    _parsedindexvalue_nextIndex_T_347; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_349 = _parsedindexvalue_nextIndex_T_320 ? parsedindexvalue_first_stage_4 :
    _parsedindexvalue_nextIndex_T_348; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_350 = _parsedindexvalue_nextIndex_T_317 ? parsedindexvalue_first_stage_4 :
    _parsedindexvalue_nextIndex_T_349; // @[Mux.scala 101:16]
  wire [1:0] parsedindexvalue_nextIndex_8 = _parsedindexvalue_nextIndex_T_314 ? parsedindexvalue_first_stage_4 :
    _parsedindexvalue_nextIndex_T_350; // @[Mux.scala 101:16]
  wire [2:0] _GEN_86 = {{1'd0}, parsedindexvalue_nextIndex_8}; // @[Benes.scala 33:40]
  wire [2:0] _GEN_87 = _GEN_86 % 3'h4; // @[Benes.scala 33:40]
  wire [1:0] parsedindexvalue_calculation_9 = _GEN_87[1:0]; // @[Benes.scala 33:40]
  wire  _parsedindexvalue_nextIndex_T_351 = parsedindexvalue_calculation_9 == 2'h0; // @[Benes.scala 35:27]
  wire  _parsedindexvalue_nextIndex_T_352 = ~parsedindexvalue_boolArray_4_1; // @[Benes.scala 35:53]
  wire  _parsedindexvalue_nextIndex_T_353 = parsedindexvalue_calculation_9 == 2'h0 & ~parsedindexvalue_boolArray_4_1; // @[Benes.scala 35:36]
  wire  _parsedindexvalue_nextIndex_T_354 = parsedindexvalue_calculation_9 == 2'h1; // @[Benes.scala 36:27]
  wire  _parsedindexvalue_nextIndex_T_356 = parsedindexvalue_calculation_9 == 2'h1 & _parsedindexvalue_nextIndex_T_352; // @[Benes.scala 36:36]
  wire  _parsedindexvalue_nextIndex_T_357 = parsedindexvalue_calculation_9 == 2'h2; // @[Benes.scala 37:27]
  wire  _parsedindexvalue_nextIndex_T_359 = parsedindexvalue_calculation_9 == 2'h2 & _parsedindexvalue_nextIndex_T_352; // @[Benes.scala 37:36]
  wire  _parsedindexvalue_nextIndex_T_360 = parsedindexvalue_calculation_9 == 2'h3; // @[Benes.scala 38:27]
  wire  _parsedindexvalue_nextIndex_T_362 = parsedindexvalue_calculation_9 == 2'h3 & _parsedindexvalue_nextIndex_T_352; // @[Benes.scala 38:36]
  wire  _parsedindexvalue_nextIndex_T_365 = _parsedindexvalue_nextIndex_T_351 & parsedindexvalue_boolArray_4_1; // @[Benes.scala 39:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_367 = parsedindexvalue_nextIndex_8 + 2'h2; // @[Benes.scala 39:76]
  wire  _parsedindexvalue_nextIndex_T_370 = _parsedindexvalue_nextIndex_T_354 & parsedindexvalue_boolArray_4_1; // @[Benes.scala 40:36]
  wire  _parsedindexvalue_nextIndex_T_375 = _parsedindexvalue_nextIndex_T_357 & parsedindexvalue_boolArray_4_1; // @[Benes.scala 41:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_377 = parsedindexvalue_nextIndex_8 - 2'h2; // @[Benes.scala 41:76]
  wire  _parsedindexvalue_nextIndex_T_380 = _parsedindexvalue_nextIndex_T_360 & parsedindexvalue_boolArray_4_1; // @[Benes.scala 42:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_383 = _parsedindexvalue_nextIndex_T_380 ? _parsedindexvalue_nextIndex_T_377
     : parsedindexvalue_nextIndex_8; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_384 = _parsedindexvalue_nextIndex_T_375 ? _parsedindexvalue_nextIndex_T_377
     : _parsedindexvalue_nextIndex_T_383; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_385 = _parsedindexvalue_nextIndex_T_370 ? _parsedindexvalue_nextIndex_T_367
     : _parsedindexvalue_nextIndex_T_384; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_386 = _parsedindexvalue_nextIndex_T_365 ? _parsedindexvalue_nextIndex_T_367
     : _parsedindexvalue_nextIndex_T_385; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_387 = _parsedindexvalue_nextIndex_T_362 ? parsedindexvalue_nextIndex_8 :
    _parsedindexvalue_nextIndex_T_386; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_388 = _parsedindexvalue_nextIndex_T_359 ? parsedindexvalue_nextIndex_8 :
    _parsedindexvalue_nextIndex_T_387; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_389 = _parsedindexvalue_nextIndex_T_356 ? parsedindexvalue_nextIndex_8 :
    _parsedindexvalue_nextIndex_T_388; // @[Mux.scala 101:16]
  wire [1:0] parsedindexvalue_nextIndex_9 = _parsedindexvalue_nextIndex_T_353 ? parsedindexvalue_nextIndex_8 :
    _parsedindexvalue_nextIndex_T_389; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_third_stage_T_33 = parsedindexvalue_nextIndex_9 % 2'h2; // @[Benes.scala 48:61]
  wire [1:0] _parsedindexvalue_third_stage_T_36 = parsedindexvalue_nextIndex_9 + 2'h1; // @[Benes.scala 48:89]
  wire [1:0] _parsedindexvalue_third_stage_T_38 = parsedindexvalue_nextIndex_9 - 2'h1; // @[Benes.scala 48:109]
  wire [1:0] _parsedindexvalue_third_stage_T_39 = _parsedindexvalue_third_stage_T_33 == 2'h0 ?
    _parsedindexvalue_third_stage_T_36 : _parsedindexvalue_third_stage_T_38; // @[Benes.scala 48:47]
  wire [1:0] parsedindexvalue_4 = io_i_mux_bus_3[3] ? _parsedindexvalue_third_stage_T_39 : parsedindexvalue_nextIndex_9; // @[Benes.scala 48:24]
  wire [2:0] _T_19 = {{1'd0}, parsedindexvalue_4};
  wire [15:0] _GEN_52 = 3'h0 == _T_19 ? io_i_data_bus2_3 : _GEN_47; // @[Benes.scala 63:{47,47}]
  wire [15:0] _GEN_53 = 3'h1 == _T_19 ? io_i_data_bus2_3 : _GEN_48; // @[Benes.scala 63:{47,47}]
  wire [15:0] _GEN_54 = 3'h2 == _T_19 ? io_i_data_bus2_3 : _GEN_49; // @[Benes.scala 63:{47,47}]
  wire [15:0] _GEN_55 = 3'h3 == _T_19 ? io_i_data_bus2_3 : _GEN_50; // @[Benes.scala 63:{47,47}]
  wire [1:0] _parsedindexvalue_first_stage_T_41 = 2'h3 % 2'h2; // @[Benes.scala 24:52]
  wire [1:0] _parsedindexvalue_first_stage_T_47 = _parsedindexvalue_first_stage_T_41 == 2'h0 ? 2'h0 :
    _parsedindexvalue_T_9; // @[Benes.scala 24:40]
  wire [1:0] parsedindexvalue_first_stage_5 = io_i_mux_bus_3[0] ? _parsedindexvalue_first_stage_T_47 : 2'h3; // @[Benes.scala 24:26]
  wire [2:0] _GEN_89 = {{1'd0}, parsedindexvalue_first_stage_5}; // @[Benes.scala 33:40]
  wire [2:0] _GEN_91 = _GEN_89 % 3'h4; // @[Benes.scala 33:40]
  wire [1:0] parsedindexvalue_calculation_10 = _GEN_91[1:0]; // @[Benes.scala 33:40]
  wire  _parsedindexvalue_nextIndex_T_390 = parsedindexvalue_calculation_10 == 2'h0; // @[Benes.scala 35:27]
  wire  _parsedindexvalue_nextIndex_T_392 = parsedindexvalue_calculation_10 == 2'h0 & ~parsedindexvalue_boolArray_4_0; // @[Benes.scala 35:36]
  wire  _parsedindexvalue_nextIndex_T_393 = parsedindexvalue_calculation_10 == 2'h1; // @[Benes.scala 36:27]
  wire  _parsedindexvalue_nextIndex_T_395 = parsedindexvalue_calculation_10 == 2'h1 & _parsedindexvalue_nextIndex_T_313; // @[Benes.scala 36:36]
  wire  _parsedindexvalue_nextIndex_T_396 = parsedindexvalue_calculation_10 == 2'h2; // @[Benes.scala 37:27]
  wire  _parsedindexvalue_nextIndex_T_398 = parsedindexvalue_calculation_10 == 2'h2 & _parsedindexvalue_nextIndex_T_313; // @[Benes.scala 37:36]
  wire  _parsedindexvalue_nextIndex_T_399 = parsedindexvalue_calculation_10 == 2'h3; // @[Benes.scala 38:27]
  wire  _parsedindexvalue_nextIndex_T_401 = parsedindexvalue_calculation_10 == 2'h3 & _parsedindexvalue_nextIndex_T_313; // @[Benes.scala 38:36]
  wire  _parsedindexvalue_nextIndex_T_404 = _parsedindexvalue_nextIndex_T_390 & parsedindexvalue_boolArray_4_0; // @[Benes.scala 39:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_406 = parsedindexvalue_first_stage_5 + 2'h2; // @[Benes.scala 39:76]
  wire  _parsedindexvalue_nextIndex_T_409 = _parsedindexvalue_nextIndex_T_393 & parsedindexvalue_boolArray_4_0; // @[Benes.scala 40:36]
  wire  _parsedindexvalue_nextIndex_T_414 = _parsedindexvalue_nextIndex_T_396 & parsedindexvalue_boolArray_4_0; // @[Benes.scala 41:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_416 = parsedindexvalue_first_stage_5 - 2'h2; // @[Benes.scala 41:76]
  wire  _parsedindexvalue_nextIndex_T_419 = _parsedindexvalue_nextIndex_T_399 & parsedindexvalue_boolArray_4_0; // @[Benes.scala 42:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_422 = _parsedindexvalue_nextIndex_T_419 ? _parsedindexvalue_nextIndex_T_416
     : parsedindexvalue_first_stage_5; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_423 = _parsedindexvalue_nextIndex_T_414 ? _parsedindexvalue_nextIndex_T_416
     : _parsedindexvalue_nextIndex_T_422; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_424 = _parsedindexvalue_nextIndex_T_409 ? _parsedindexvalue_nextIndex_T_406
     : _parsedindexvalue_nextIndex_T_423; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_425 = _parsedindexvalue_nextIndex_T_404 ? _parsedindexvalue_nextIndex_T_406
     : _parsedindexvalue_nextIndex_T_424; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_426 = _parsedindexvalue_nextIndex_T_401 ? parsedindexvalue_first_stage_5 :
    _parsedindexvalue_nextIndex_T_425; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_427 = _parsedindexvalue_nextIndex_T_398 ? parsedindexvalue_first_stage_5 :
    _parsedindexvalue_nextIndex_T_426; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_428 = _parsedindexvalue_nextIndex_T_395 ? parsedindexvalue_first_stage_5 :
    _parsedindexvalue_nextIndex_T_427; // @[Mux.scala 101:16]
  wire [1:0] parsedindexvalue_nextIndex_10 = _parsedindexvalue_nextIndex_T_392 ? parsedindexvalue_first_stage_5 :
    _parsedindexvalue_nextIndex_T_428; // @[Mux.scala 101:16]
  wire [2:0] _GEN_92 = {{1'd0}, parsedindexvalue_nextIndex_10}; // @[Benes.scala 33:40]
  wire [2:0] _GEN_93 = _GEN_92 % 3'h4; // @[Benes.scala 33:40]
  wire [1:0] parsedindexvalue_calculation_11 = _GEN_93[1:0]; // @[Benes.scala 33:40]
  wire  _parsedindexvalue_nextIndex_T_429 = parsedindexvalue_calculation_11 == 2'h0; // @[Benes.scala 35:27]
  wire  _parsedindexvalue_nextIndex_T_431 = parsedindexvalue_calculation_11 == 2'h0 & ~parsedindexvalue_boolArray_4_1; // @[Benes.scala 35:36]
  wire  _parsedindexvalue_nextIndex_T_432 = parsedindexvalue_calculation_11 == 2'h1; // @[Benes.scala 36:27]
  wire  _parsedindexvalue_nextIndex_T_434 = parsedindexvalue_calculation_11 == 2'h1 & _parsedindexvalue_nextIndex_T_352; // @[Benes.scala 36:36]
  wire  _parsedindexvalue_nextIndex_T_435 = parsedindexvalue_calculation_11 == 2'h2; // @[Benes.scala 37:27]
  wire  _parsedindexvalue_nextIndex_T_437 = parsedindexvalue_calculation_11 == 2'h2 & _parsedindexvalue_nextIndex_T_352; // @[Benes.scala 37:36]
  wire  _parsedindexvalue_nextIndex_T_438 = parsedindexvalue_calculation_11 == 2'h3; // @[Benes.scala 38:27]
  wire  _parsedindexvalue_nextIndex_T_440 = parsedindexvalue_calculation_11 == 2'h3 & _parsedindexvalue_nextIndex_T_352; // @[Benes.scala 38:36]
  wire  _parsedindexvalue_nextIndex_T_443 = _parsedindexvalue_nextIndex_T_429 & parsedindexvalue_boolArray_4_1; // @[Benes.scala 39:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_445 = parsedindexvalue_nextIndex_10 + 2'h2; // @[Benes.scala 39:76]
  wire  _parsedindexvalue_nextIndex_T_448 = _parsedindexvalue_nextIndex_T_432 & parsedindexvalue_boolArray_4_1; // @[Benes.scala 40:36]
  wire  _parsedindexvalue_nextIndex_T_453 = _parsedindexvalue_nextIndex_T_435 & parsedindexvalue_boolArray_4_1; // @[Benes.scala 41:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_455 = parsedindexvalue_nextIndex_10 - 2'h2; // @[Benes.scala 41:76]
  wire  _parsedindexvalue_nextIndex_T_458 = _parsedindexvalue_nextIndex_T_438 & parsedindexvalue_boolArray_4_1; // @[Benes.scala 42:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_461 = _parsedindexvalue_nextIndex_T_458 ? _parsedindexvalue_nextIndex_T_455
     : parsedindexvalue_nextIndex_10; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_462 = _parsedindexvalue_nextIndex_T_453 ? _parsedindexvalue_nextIndex_T_455
     : _parsedindexvalue_nextIndex_T_461; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_463 = _parsedindexvalue_nextIndex_T_448 ? _parsedindexvalue_nextIndex_T_445
     : _parsedindexvalue_nextIndex_T_462; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_464 = _parsedindexvalue_nextIndex_T_443 ? _parsedindexvalue_nextIndex_T_445
     : _parsedindexvalue_nextIndex_T_463; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_465 = _parsedindexvalue_nextIndex_T_440 ? parsedindexvalue_nextIndex_10 :
    _parsedindexvalue_nextIndex_T_464; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_466 = _parsedindexvalue_nextIndex_T_437 ? parsedindexvalue_nextIndex_10 :
    _parsedindexvalue_nextIndex_T_465; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_467 = _parsedindexvalue_nextIndex_T_434 ? parsedindexvalue_nextIndex_10 :
    _parsedindexvalue_nextIndex_T_466; // @[Mux.scala 101:16]
  wire [1:0] parsedindexvalue_nextIndex_11 = _parsedindexvalue_nextIndex_T_431 ? parsedindexvalue_nextIndex_10 :
    _parsedindexvalue_nextIndex_T_467; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_third_stage_T_41 = parsedindexvalue_nextIndex_11 % 2'h2; // @[Benes.scala 48:61]
  wire [1:0] _parsedindexvalue_third_stage_T_44 = parsedindexvalue_nextIndex_11 + 2'h1; // @[Benes.scala 48:89]
  wire [1:0] _parsedindexvalue_third_stage_T_46 = parsedindexvalue_nextIndex_11 - 2'h1; // @[Benes.scala 48:109]
  wire [1:0] _parsedindexvalue_third_stage_T_47 = _parsedindexvalue_third_stage_T_41 == 2'h0 ?
    _parsedindexvalue_third_stage_T_44 : _parsedindexvalue_third_stage_T_46; // @[Benes.scala 48:47]
  wire [1:0] parsedindexvalue_5 = io_i_mux_bus_3[3] ? _parsedindexvalue_third_stage_T_47 : parsedindexvalue_nextIndex_11
    ; // @[Benes.scala 48:24]
  wire [2:0] _T_21 = {{1'd0}, parsedindexvalue_5};
  wire [15:0] _GEN_57 = 3'h0 == _T_21 ? io_i_data_bus2_3 : _GEN_47; // @[Benes.scala 67:{47,47}]
  wire [15:0] _GEN_58 = 3'h1 == _T_21 ? io_i_data_bus2_3 : _GEN_48; // @[Benes.scala 67:{47,47}]
  wire [15:0] _GEN_59 = 3'h2 == _T_21 ? io_i_data_bus2_3 : _GEN_49; // @[Benes.scala 67:{47,47}]
  wire [15:0] _GEN_60 = 3'h3 == _T_21 ? io_i_data_bus2_3 : _GEN_50; // @[Benes.scala 67:{47,47}]
  wire [15:0] _GEN_62 = io_i_data_bus2_3 == io_i_data_bus2_2 ? _GEN_52 : _GEN_57; // @[Benes.scala 60:61]
  wire [15:0] _GEN_63 = io_i_data_bus2_3 == io_i_data_bus2_2 ? _GEN_53 : _GEN_58; // @[Benes.scala 60:61]
  wire [15:0] _GEN_64 = io_i_data_bus2_3 == io_i_data_bus2_2 ? _GEN_54 : _GEN_59; // @[Benes.scala 60:61]
  wire [15:0] _GEN_65 = io_i_data_bus2_3 == io_i_data_bus2_2 ? _GEN_55 : _GEN_60; // @[Benes.scala 60:61]
  wire [15:0] _GEN_67 = _T_18 ? 16'h0 : io_i_data_bus2_3; // @[Benes.scala 72:60 74:28 78:28]
  wire [15:0] _GEN_68 = |io_i_mux_bus_3 ? _GEN_62 : _GEN_47; // @[Benes.scala 58:35]
  wire [15:0] _GEN_69 = |io_i_mux_bus_3 ? _GEN_63 : _GEN_48; // @[Benes.scala 58:35]
  wire [15:0] _GEN_70 = |io_i_mux_bus_3 ? _GEN_64 : _GEN_49; // @[Benes.scala 58:35]
  wire [15:0] _GEN_71 = |io_i_mux_bus_3 ? _GEN_65 : _GEN_67; // @[Benes.scala 58:35]
  wire [15:0] _GEN_73 = io_i_data_bus2_3 != 16'h0 ? _GEN_68 : _GEN_47; // @[Benes.scala 56:39]
  wire [15:0] _GEN_74 = io_i_data_bus2_3 != 16'h0 ? _GEN_69 : _GEN_48; // @[Benes.scala 56:39]
  wire [15:0] _GEN_75 = io_i_data_bus2_3 != 16'h0 ? _GEN_70 : _GEN_49; // @[Benes.scala 56:39]
  wire [15:0] _GEN_76 = io_i_data_bus2_3 != 16'h0 ? _GEN_71 : _GEN_50; // @[Benes.scala 56:39]
  wire  parsedindexvalue_first_stage_6 = io_i_mux_bus_0[0] & (~_GEN_4[0] | 1'h0 - 1'h1); // @[Benes.scala 24:26]
  wire  parsedindexvalue_boolArray_6_0 = io_i_mux_bus_0[1]; // @[Benes.scala 28:92]
  wire  parsedindexvalue_boolArray_6_1 = io_i_mux_bus_0[2]; // @[Benes.scala 28:92]
  wire [2:0] _GEN_94 = {{2'd0}, parsedindexvalue_first_stage_6}; // @[Benes.scala 33:40]
  wire [2:0] _GEN_95 = _GEN_94 % 3'h4; // @[Benes.scala 33:40]
  wire  parsedindexvalue_calculation_12 = _GEN_95[0]; // @[Benes.scala 33:40]
  wire  _parsedindexvalue_nextIndex_T_468 = ~parsedindexvalue_calculation_12; // @[Benes.scala 35:27]
  wire  _parsedindexvalue_nextIndex_T_469 = ~parsedindexvalue_boolArray_6_0; // @[Benes.scala 35:53]
  wire  _parsedindexvalue_nextIndex_T_470 = ~parsedindexvalue_calculation_12 & ~parsedindexvalue_boolArray_6_0; // @[Benes.scala 35:36]
  wire  _parsedindexvalue_nextIndex_T_473 = parsedindexvalue_calculation_12 & _parsedindexvalue_nextIndex_T_469; // @[Benes.scala 36:36]
  wire [1:0] _GEN_104 = {{1'd0}, parsedindexvalue_calculation_12}; // @[Benes.scala 37:27]
  wire  _parsedindexvalue_nextIndex_T_474 = _GEN_104 == 2'h2; // @[Benes.scala 37:27]
  wire  _parsedindexvalue_nextIndex_T_476 = _GEN_104 == 2'h2 & _parsedindexvalue_nextIndex_T_469; // @[Benes.scala 37:36]
  wire  _parsedindexvalue_nextIndex_T_477 = _GEN_104 == 2'h3; // @[Benes.scala 38:27]
  wire  _parsedindexvalue_nextIndex_T_479 = _GEN_104 == 2'h3 & _parsedindexvalue_nextIndex_T_469; // @[Benes.scala 38:36]
  wire  _parsedindexvalue_nextIndex_T_482 = _parsedindexvalue_nextIndex_T_468 & parsedindexvalue_boolArray_6_0; // @[Benes.scala 39:36]
  wire [1:0] _GEN_106 = {{1'd0}, parsedindexvalue_first_stage_6}; // @[Benes.scala 39:76]
  wire [1:0] _parsedindexvalue_nextIndex_T_484 = _GEN_106 + 2'h2; // @[Benes.scala 39:76]
  wire  _parsedindexvalue_nextIndex_T_487 = parsedindexvalue_calculation_12 & parsedindexvalue_boolArray_6_0; // @[Benes.scala 40:36]
  wire  _parsedindexvalue_nextIndex_T_492 = _parsedindexvalue_nextIndex_T_474 & parsedindexvalue_boolArray_6_0; // @[Benes.scala 41:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_494 = _GEN_106 - 2'h2; // @[Benes.scala 41:76]
  wire  _parsedindexvalue_nextIndex_T_497 = _parsedindexvalue_nextIndex_T_477 & parsedindexvalue_boolArray_6_0; // @[Benes.scala 42:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_500 = _parsedindexvalue_nextIndex_T_497 ? _parsedindexvalue_nextIndex_T_494
     : {{1'd0}, parsedindexvalue_first_stage_6}; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_501 = _parsedindexvalue_nextIndex_T_492 ? _parsedindexvalue_nextIndex_T_494
     : _parsedindexvalue_nextIndex_T_500; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_502 = _parsedindexvalue_nextIndex_T_487 ? _parsedindexvalue_nextIndex_T_484
     : _parsedindexvalue_nextIndex_T_501; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_503 = _parsedindexvalue_nextIndex_T_482 ? _parsedindexvalue_nextIndex_T_484
     : _parsedindexvalue_nextIndex_T_502; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_504 = _parsedindexvalue_nextIndex_T_479 ? {{1'd0},
    parsedindexvalue_first_stage_6} : _parsedindexvalue_nextIndex_T_503; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_505 = _parsedindexvalue_nextIndex_T_476 ? {{1'd0},
    parsedindexvalue_first_stage_6} : _parsedindexvalue_nextIndex_T_504; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_506 = _parsedindexvalue_nextIndex_T_473 ? {{1'd0},
    parsedindexvalue_first_stage_6} : _parsedindexvalue_nextIndex_T_505; // @[Mux.scala 101:16]
  wire [1:0] parsedindexvalue_nextIndex_12 = _parsedindexvalue_nextIndex_T_470 ? {{1'd0}, parsedindexvalue_first_stage_6
    } : _parsedindexvalue_nextIndex_T_506; // @[Mux.scala 101:16]
  wire [2:0] _GEN_97 = {{1'd0}, parsedindexvalue_nextIndex_12}; // @[Benes.scala 33:40]
  wire [2:0] _GEN_99 = _GEN_97 % 3'h4; // @[Benes.scala 33:40]
  wire [1:0] parsedindexvalue_calculation_13 = _GEN_99[1:0]; // @[Benes.scala 33:40]
  wire  _parsedindexvalue_nextIndex_T_507 = parsedindexvalue_calculation_13 == 2'h0; // @[Benes.scala 35:27]
  wire  _parsedindexvalue_nextIndex_T_508 = ~parsedindexvalue_boolArray_6_1; // @[Benes.scala 35:53]
  wire  _parsedindexvalue_nextIndex_T_509 = parsedindexvalue_calculation_13 == 2'h0 & ~parsedindexvalue_boolArray_6_1; // @[Benes.scala 35:36]
  wire  _parsedindexvalue_nextIndex_T_510 = parsedindexvalue_calculation_13 == 2'h1; // @[Benes.scala 36:27]
  wire  _parsedindexvalue_nextIndex_T_512 = parsedindexvalue_calculation_13 == 2'h1 & _parsedindexvalue_nextIndex_T_508; // @[Benes.scala 36:36]
  wire  _parsedindexvalue_nextIndex_T_513 = parsedindexvalue_calculation_13 == 2'h2; // @[Benes.scala 37:27]
  wire  _parsedindexvalue_nextIndex_T_515 = parsedindexvalue_calculation_13 == 2'h2 & _parsedindexvalue_nextIndex_T_508; // @[Benes.scala 37:36]
  wire  _parsedindexvalue_nextIndex_T_516 = parsedindexvalue_calculation_13 == 2'h3; // @[Benes.scala 38:27]
  wire  _parsedindexvalue_nextIndex_T_518 = parsedindexvalue_calculation_13 == 2'h3 & _parsedindexvalue_nextIndex_T_508; // @[Benes.scala 38:36]
  wire  _parsedindexvalue_nextIndex_T_521 = _parsedindexvalue_nextIndex_T_507 & parsedindexvalue_boolArray_6_1; // @[Benes.scala 39:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_523 = parsedindexvalue_nextIndex_12 + 2'h2; // @[Benes.scala 39:76]
  wire  _parsedindexvalue_nextIndex_T_526 = _parsedindexvalue_nextIndex_T_510 & parsedindexvalue_boolArray_6_1; // @[Benes.scala 40:36]
  wire  _parsedindexvalue_nextIndex_T_531 = _parsedindexvalue_nextIndex_T_513 & parsedindexvalue_boolArray_6_1; // @[Benes.scala 41:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_533 = parsedindexvalue_nextIndex_12 - 2'h2; // @[Benes.scala 41:76]
  wire  _parsedindexvalue_nextIndex_T_536 = _parsedindexvalue_nextIndex_T_516 & parsedindexvalue_boolArray_6_1; // @[Benes.scala 42:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_539 = _parsedindexvalue_nextIndex_T_536 ? _parsedindexvalue_nextIndex_T_533
     : parsedindexvalue_nextIndex_12; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_540 = _parsedindexvalue_nextIndex_T_531 ? _parsedindexvalue_nextIndex_T_533
     : _parsedindexvalue_nextIndex_T_539; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_541 = _parsedindexvalue_nextIndex_T_526 ? _parsedindexvalue_nextIndex_T_523
     : _parsedindexvalue_nextIndex_T_540; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_542 = _parsedindexvalue_nextIndex_T_521 ? _parsedindexvalue_nextIndex_T_523
     : _parsedindexvalue_nextIndex_T_541; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_543 = _parsedindexvalue_nextIndex_T_518 ? parsedindexvalue_nextIndex_12 :
    _parsedindexvalue_nextIndex_T_542; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_544 = _parsedindexvalue_nextIndex_T_515 ? parsedindexvalue_nextIndex_12 :
    _parsedindexvalue_nextIndex_T_543; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_545 = _parsedindexvalue_nextIndex_T_512 ? parsedindexvalue_nextIndex_12 :
    _parsedindexvalue_nextIndex_T_544; // @[Mux.scala 101:16]
  wire [1:0] parsedindexvalue_nextIndex_13 = _parsedindexvalue_nextIndex_T_509 ? parsedindexvalue_nextIndex_12 :
    _parsedindexvalue_nextIndex_T_545; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_third_stage_T_49 = parsedindexvalue_nextIndex_13 % 2'h2; // @[Benes.scala 48:61]
  wire [1:0] _parsedindexvalue_third_stage_T_52 = parsedindexvalue_nextIndex_13 + 2'h1; // @[Benes.scala 48:89]
  wire [1:0] _parsedindexvalue_third_stage_T_54 = parsedindexvalue_nextIndex_13 - 2'h1; // @[Benes.scala 48:109]
  wire [1:0] _parsedindexvalue_third_stage_T_55 = _parsedindexvalue_third_stage_T_49 == 2'h0 ?
    _parsedindexvalue_third_stage_T_52 : _parsedindexvalue_third_stage_T_54; // @[Benes.scala 48:47]
  wire [1:0] parsedindexvalue_6 = io_i_mux_bus_0[3] ? _parsedindexvalue_third_stage_T_55 : parsedindexvalue_nextIndex_13
    ; // @[Benes.scala 48:24]
  wire [2:0] _T_25 = {{1'd0}, parsedindexvalue_6};
  wire [15:0] _GEN_78 = 3'h0 == _T_25 ? io_i_data_bus2_0 : _GEN_73; // @[Benes.scala 94:{35,35}]
  wire [15:0] _GEN_79 = 3'h1 == _T_25 ? io_i_data_bus2_0 : _GEN_74; // @[Benes.scala 94:{35,35}]
  wire [15:0] _GEN_80 = 3'h2 == _T_25 ? io_i_data_bus2_0 : _GEN_75; // @[Benes.scala 94:{35,35}]
  wire [15:0] _GEN_81 = 3'h3 == _T_25 ? io_i_data_bus2_0 : _GEN_76; // @[Benes.scala 94:{35,35}]
  assign io_o_dist_bus1_0 = io_i_data_bus1_0; // @[Benes.scala 16:18]
  assign io_o_dist_bus1_1 = io_i_data_bus1_1; // @[Benes.scala 16:18]
  assign io_o_dist_bus1_2 = io_i_data_bus1_2; // @[Benes.scala 16:18]
  assign io_o_dist_bus1_3 = io_i_data_bus1_3; // @[Benes.scala 16:18]
  assign io_o_dist_bus2_0 = io_i_data_bus2_0 != 16'h0 ? _GEN_78 : _GEN_73; // @[Benes.scala 91:35]
  assign io_o_dist_bus2_1 = io_i_data_bus2_0 != 16'h0 ? _GEN_79 : _GEN_74; // @[Benes.scala 91:35]
  assign io_o_dist_bus2_2 = io_i_data_bus2_0 != 16'h0 ? _GEN_80 : _GEN_75; // @[Benes.scala 91:35]
  assign io_o_dist_bus2_3 = io_i_data_bus2_0 != 16'h0 ? _GEN_81 : _GEN_76; // @[Benes.scala 91:35]
endmodule
module buffer_multiplication(
  input  [15:0] io_buffer1_0,
  input  [15:0] io_buffer1_1,
  input  [15:0] io_buffer1_2,
  input  [15:0] io_buffer1_3,
  input  [15:0] io_buffer2_0,
  input  [15:0] io_buffer2_1,
  input  [15:0] io_buffer2_2,
  input  [15:0] io_buffer2_3,
  output [15:0] io_out_0,
  output [15:0] io_out_1,
  output [15:0] io_out_2,
  output [15:0] io_out_3
);
  wire [31:0] elementMul = io_buffer1_0 * io_buffer2_0; // @[buffer_multiplication.scala 17:42]
  wire [31:0] result_elementMul = io_buffer1_1 * io_buffer2_1; // @[buffer_multiplication.scala 17:42]
  wire [31:0] result_result_elementMul = io_buffer1_2 * io_buffer2_2; // @[buffer_multiplication.scala 17:42]
  wire [31:0] result_result_result_elementMul = io_buffer1_3 * io_buffer2_3; // @[buffer_multiplication.scala 17:42]
  assign io_out_0 = elementMul[15:0]; // @[buffer_multiplication.scala 15:20 19:27]
  assign io_out_1 = result_elementMul[15:0]; // @[buffer_multiplication.scala 15:20 19:27]
  assign io_out_2 = result_result_elementMul[15:0]; // @[buffer_multiplication.scala 15:20 19:27]
  assign io_out_3 = result_result_result_elementMul[15:0]; // @[buffer_multiplication.scala 15:20 19:27]
endmodule
module ReductionMux(
  input  [31:0] io_i_data_0,
  input  [31:0] io_i_data_1,
  output [31:0] io_o_data_0,
  output [31:0] io_o_data_1
);
  assign io_o_data_0 = io_i_data_0; // @[ReductionMux.scala 31:39 33:18 35:18]
  assign io_o_data_1 = io_i_data_1; // @[ReductionMux.scala 37:22]
endmodule
module SimpleAdder(
  input  [31:0] io_A,
  input  [31:0] io_B,
  output [31:0] io_O
);
  assign io_O = io_A + io_B; // @[SimpleAdder.scala 14:18]
endmodule
module EdgeAdderSwitch(
  input         clock,
  input         reset,
  input         io_i_valid,
  input  [63:0] io_i_data_bus_0,
  input  [63:0] io_i_data_bus_1,
  input  [2:0]  io_i_add_en,
  input  [4:0]  io_i_cmd,
  output [31:0] io_o_adder
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] reductionMux_io_i_data_0; // @[EdgeAdderSwitch.scala 19:28]
  wire [31:0] reductionMux_io_i_data_1; // @[EdgeAdderSwitch.scala 19:28]
  wire [31:0] reductionMux_io_o_data_0; // @[EdgeAdderSwitch.scala 19:28]
  wire [31:0] reductionMux_io_o_data_1; // @[EdgeAdderSwitch.scala 19:28]
  wire [31:0] adder32_io_A; // @[EdgeAdderSwitch.scala 23:23]
  wire [31:0] adder32_io_B; // @[EdgeAdderSwitch.scala 23:23]
  wire [31:0] adder32_io_O; // @[EdgeAdderSwitch.scala 23:23]
  reg  r_valid; // @[EdgeAdderSwitch.scala 27:24]
  reg [31:0] r_adder; // @[EdgeAdderSwitch.scala 28:24]
  reg [2:0] r_add_en; // @[EdgeAdderSwitch.scala 31:25]
  wire [31:0] _GEN_3 = 5'h4 == io_i_cmd ? reductionMux_io_o_data_0 : r_adder; // @[EdgeAdderSwitch.scala 38:23 45:17 28:24]
  wire [31:0] _GEN_15 = r_add_en == 3'h0 ? r_adder : adder32_io_O; // @[EdgeAdderSwitch.scala 64:22 65:18 67:18]
  ReductionMux reductionMux ( // @[EdgeAdderSwitch.scala 19:28]
    .io_i_data_0(reductionMux_io_i_data_0),
    .io_i_data_1(reductionMux_io_i_data_1),
    .io_o_data_0(reductionMux_io_o_data_0),
    .io_o_data_1(reductionMux_io_o_data_1)
  );
  SimpleAdder adder32 ( // @[EdgeAdderSwitch.scala 23:23]
    .io_A(adder32_io_A),
    .io_B(adder32_io_B),
    .io_O(adder32_io_O)
  );
  assign io_o_adder = reset ? 32'h0 : _GEN_15; // @[EdgeAdderSwitch.scala 59:14 60:16]
  assign reductionMux_io_i_data_0 = io_i_data_bus_0[31:0]; // @[EdgeAdderSwitch.scala 20:26]
  assign reductionMux_io_i_data_1 = io_i_data_bus_1[31:0]; // @[EdgeAdderSwitch.scala 20:26]
  assign adder32_io_A = reductionMux_io_o_data_1; // @[EdgeAdderSwitch.scala 24:16]
  assign adder32_io_B = reductionMux_io_o_data_0; // @[EdgeAdderSwitch.scala 25:16]
  always @(posedge clock) begin
    if (reset) begin // @[EdgeAdderSwitch.scala 27:24]
      r_valid <= 1'h0; // @[EdgeAdderSwitch.scala 27:24]
    end else begin
      r_valid <= io_i_valid; // @[EdgeAdderSwitch.scala 27:24]
    end
    if (reset) begin // @[EdgeAdderSwitch.scala 28:24]
      r_adder <= 32'h0; // @[EdgeAdderSwitch.scala 28:24]
    end else if (reset) begin // @[EdgeAdderSwitch.scala 33:14]
      r_adder <= 32'h0; // @[EdgeAdderSwitch.scala 34:13]
    end else if (r_valid) begin // @[EdgeAdderSwitch.scala 37:25]
      if (5'h3 == io_i_cmd) begin // @[EdgeAdderSwitch.scala 38:23]
        r_adder <= reductionMux_io_o_data_1; // @[EdgeAdderSwitch.scala 40:17]
      end else begin
        r_adder <= _GEN_3;
      end
    end
    if (reset) begin // @[EdgeAdderSwitch.scala 31:25]
      r_add_en <= 3'h0; // @[EdgeAdderSwitch.scala 31:25]
    end else begin
      r_add_en <= io_i_add_en; // @[EdgeAdderSwitch.scala 31:25]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  r_adder = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  r_add_en = _RAND_2[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Fan4(
  input         clock,
  input         reset,
  input         io_i_valid,
  input  [31:0] io_i_data_bus_0,
  input  [31:0] io_i_data_bus_1,
  input  [31:0] io_i_data_bus_2,
  input  [31:0] io_i_data_bus_3,
  input         io_i_add_en_bus_0,
  input         io_i_add_en_bus_1,
  input         io_i_add_en_bus_2,
  input  [2:0]  io_i_cmd_bus_0,
  input  [2:0]  io_i_cmd_bus_1,
  input  [2:0]  io_i_cmd_bus_2,
  output [31:0] io_o_adder_0,
  output [31:0] io_o_adder_1,
  output [31:0] io_o_adder_2
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  my_adder_0_clock; // @[FanNetwork.scala 119:28]
  wire  my_adder_0_reset; // @[FanNetwork.scala 119:28]
  wire  my_adder_0_io_i_valid; // @[FanNetwork.scala 119:28]
  wire [63:0] my_adder_0_io_i_data_bus_0; // @[FanNetwork.scala 119:28]
  wire [63:0] my_adder_0_io_i_data_bus_1; // @[FanNetwork.scala 119:28]
  wire [2:0] my_adder_0_io_i_add_en; // @[FanNetwork.scala 119:28]
  wire [4:0] my_adder_0_io_i_cmd; // @[FanNetwork.scala 119:28]
  wire [31:0] my_adder_0_io_o_adder; // @[FanNetwork.scala 119:28]
  wire  my_adder_1_clock; // @[FanNetwork.scala 132:28]
  wire  my_adder_1_reset; // @[FanNetwork.scala 132:28]
  wire  my_adder_1_io_i_valid; // @[FanNetwork.scala 132:28]
  wire [63:0] my_adder_1_io_i_data_bus_0; // @[FanNetwork.scala 132:28]
  wire [63:0] my_adder_1_io_i_data_bus_1; // @[FanNetwork.scala 132:28]
  wire [2:0] my_adder_1_io_i_add_en; // @[FanNetwork.scala 132:28]
  wire [4:0] my_adder_1_io_i_cmd; // @[FanNetwork.scala 132:28]
  wire [31:0] my_adder_1_io_o_adder; // @[FanNetwork.scala 132:28]
  wire  my_adder_2_clock; // @[FanNetwork.scala 145:28]
  wire  my_adder_2_reset; // @[FanNetwork.scala 145:28]
  wire  my_adder_2_io_i_valid; // @[FanNetwork.scala 145:28]
  wire [63:0] my_adder_2_io_i_data_bus_0; // @[FanNetwork.scala 145:28]
  wire [63:0] my_adder_2_io_i_data_bus_1; // @[FanNetwork.scala 145:28]
  wire [2:0] my_adder_2_io_i_add_en; // @[FanNetwork.scala 145:28]
  wire [4:0] my_adder_2_io_i_cmd; // @[FanNetwork.scala 145:28]
  wire [31:0] my_adder_2_io_o_adder; // @[FanNetwork.scala 145:28]
  reg  r_valid_0; // @[FanNetwork.scala 30:26]
  reg  r_valid_1; // @[FanNetwork.scala 30:26]
  wire [63:0] w_fan_lvl_0_0 = {{32'd0}, my_adder_0_io_o_adder};
  wire [63:0] w_fan_lvl_0_1 = {{32'd0}, my_adder_2_io_o_adder};
  EdgeAdderSwitch my_adder_0 ( // @[FanNetwork.scala 119:28]
    .clock(my_adder_0_clock),
    .reset(my_adder_0_reset),
    .io_i_valid(my_adder_0_io_i_valid),
    .io_i_data_bus_0(my_adder_0_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_0_io_i_data_bus_1),
    .io_i_add_en(my_adder_0_io_i_add_en),
    .io_i_cmd(my_adder_0_io_i_cmd),
    .io_o_adder(my_adder_0_io_o_adder)
  );
  EdgeAdderSwitch my_adder_1 ( // @[FanNetwork.scala 132:28]
    .clock(my_adder_1_clock),
    .reset(my_adder_1_reset),
    .io_i_valid(my_adder_1_io_i_valid),
    .io_i_data_bus_0(my_adder_1_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_1_io_i_data_bus_1),
    .io_i_add_en(my_adder_1_io_i_add_en),
    .io_i_cmd(my_adder_1_io_i_cmd),
    .io_o_adder(my_adder_1_io_o_adder)
  );
  EdgeAdderSwitch my_adder_2 ( // @[FanNetwork.scala 145:28]
    .clock(my_adder_2_clock),
    .reset(my_adder_2_reset),
    .io_i_valid(my_adder_2_io_i_valid),
    .io_i_data_bus_0(my_adder_2_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_2_io_i_data_bus_1),
    .io_i_add_en(my_adder_2_io_i_add_en),
    .io_i_cmd(my_adder_2_io_i_cmd),
    .io_o_adder(my_adder_2_io_o_adder)
  );
  assign io_o_adder_0 = w_fan_lvl_0_0[31:0]; // @[FanNetwork.scala 207:19]
  assign io_o_adder_1 = my_adder_1_io_o_adder; // @[FanNetwork.scala 208:19]
  assign io_o_adder_2 = w_fan_lvl_0_1[31:0]; // @[FanNetwork.scala 209:19]
  assign my_adder_0_clock = clock;
  assign my_adder_0_reset = reset;
  assign my_adder_0_io_i_valid = r_valid_0; // @[FanNetwork.scala 121:27]
  assign my_adder_0_io_i_data_bus_0 = {{32'd0}, io_i_data_bus_1}; // @[FanNetwork.scala 122:30]
  assign my_adder_0_io_i_data_bus_1 = {{32'd0}, io_i_data_bus_0}; // @[FanNetwork.scala 122:30]
  assign my_adder_0_io_i_add_en = {{2'd0}, io_i_add_en_bus_0}; // @[FanNetwork.scala 123:28]
  assign my_adder_0_io_i_cmd = {{2'd0}, io_i_cmd_bus_0}; // @[FanNetwork.scala 124:25]
  assign my_adder_1_clock = clock;
  assign my_adder_1_reset = reset;
  assign my_adder_1_io_i_valid = r_valid_1; // @[FanNetwork.scala 134:27]
  assign my_adder_1_io_i_data_bus_0 = {{32'd0}, my_adder_2_io_o_adder}; // @[FanNetwork.scala 135:{40,40}]
  assign my_adder_1_io_i_data_bus_1 = {{32'd0}, my_adder_0_io_o_adder}; // @[FanNetwork.scala 135:{40,40}]
  assign my_adder_1_io_i_add_en = {{2'd0}, io_i_add_en_bus_2}; // @[FanNetwork.scala 136:28]
  assign my_adder_1_io_i_cmd = {{2'd0}, io_i_cmd_bus_2}; // @[FanNetwork.scala 137:26]
  assign my_adder_2_clock = clock;
  assign my_adder_2_reset = reset;
  assign my_adder_2_io_i_valid = r_valid_0; // @[FanNetwork.scala 147:27]
  assign my_adder_2_io_i_data_bus_0 = {{32'd0}, io_i_data_bus_3}; // @[FanNetwork.scala 148:30]
  assign my_adder_2_io_i_data_bus_1 = {{32'd0}, io_i_data_bus_2}; // @[FanNetwork.scala 148:30]
  assign my_adder_2_io_i_add_en = {{2'd0}, io_i_add_en_bus_1}; // @[FanNetwork.scala 149:28]
  assign my_adder_2_io_i_cmd = {{2'd0}, io_i_cmd_bus_1}; // @[FanNetwork.scala 150:25]
  always @(posedge clock) begin
    if (reset) begin // @[FanNetwork.scala 30:26]
      r_valid_0 <= 1'h0; // @[FanNetwork.scala 30:26]
    end else begin
      r_valid_0 <= io_i_valid;
    end
    if (reset) begin // @[FanNetwork.scala 30:26]
      r_valid_1 <= 1'h0; // @[FanNetwork.scala 30:26]
    end else begin
      r_valid_1 <= r_valid_0; // @[FanNetwork.scala 114:24]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_valid_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  r_valid_1 = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module flexdpecom4(
  input         clock,
  input         reset,
  input         io_i_data_valid,
  input  [15:0] io_i_data_bus_0,
  input  [15:0] io_i_data_bus_1,
  input  [15:0] io_i_data_bus_2,
  input  [15:0] io_i_data_bus_3,
  input  [15:0] io_i_data_bus2_0,
  input  [15:0] io_i_data_bus2_1,
  input  [15:0] io_i_data_bus2_2,
  input  [15:0] io_i_data_bus2_3,
  output [15:0] io_o_adder_0,
  output [15:0] io_o_adder_1,
  output [15:0] io_o_adder_2,
  input  [3:0]  io_i_mux_bus_0,
  input  [3:0]  io_i_mux_bus_1,
  input  [3:0]  io_i_mux_bus_2,
  input  [3:0]  io_i_mux_bus_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
`endif // RANDOMIZE_REG_INIT
  wire  my_controller_clock; // @[FlexDPE.scala 55:31]
  wire  my_controller_reset; // @[FlexDPE.scala 55:31]
  wire  my_controller_io_i_data_valid; // @[FlexDPE.scala 55:31]
  wire  my_controller_io_o_reduction_add_0; // @[FlexDPE.scala 55:31]
  wire  my_controller_io_o_reduction_add_1; // @[FlexDPE.scala 55:31]
  wire  my_controller_io_o_reduction_add_2; // @[FlexDPE.scala 55:31]
  wire [2:0] my_controller_io_o_reduction_cmd_0; // @[FlexDPE.scala 55:31]
  wire [2:0] my_controller_io_o_reduction_cmd_1; // @[FlexDPE.scala 55:31]
  wire [2:0] my_controller_io_o_reduction_cmd_2; // @[FlexDPE.scala 55:31]
  wire  my_controller_io_o_reduction_valid; // @[FlexDPE.scala 55:31]
  wire [15:0] my_Benes_io_i_data_bus2_0; // @[FlexDPE.scala 64:26]
  wire [15:0] my_Benes_io_i_data_bus2_1; // @[FlexDPE.scala 64:26]
  wire [15:0] my_Benes_io_i_data_bus2_2; // @[FlexDPE.scala 64:26]
  wire [15:0] my_Benes_io_i_data_bus2_3; // @[FlexDPE.scala 64:26]
  wire [15:0] my_Benes_io_i_data_bus1_0; // @[FlexDPE.scala 64:26]
  wire [15:0] my_Benes_io_i_data_bus1_1; // @[FlexDPE.scala 64:26]
  wire [15:0] my_Benes_io_i_data_bus1_2; // @[FlexDPE.scala 64:26]
  wire [15:0] my_Benes_io_i_data_bus1_3; // @[FlexDPE.scala 64:26]
  wire [3:0] my_Benes_io_i_mux_bus_0; // @[FlexDPE.scala 64:26]
  wire [3:0] my_Benes_io_i_mux_bus_1; // @[FlexDPE.scala 64:26]
  wire [3:0] my_Benes_io_i_mux_bus_2; // @[FlexDPE.scala 64:26]
  wire [3:0] my_Benes_io_i_mux_bus_3; // @[FlexDPE.scala 64:26]
  wire [15:0] my_Benes_io_o_dist_bus1_0; // @[FlexDPE.scala 64:26]
  wire [15:0] my_Benes_io_o_dist_bus1_1; // @[FlexDPE.scala 64:26]
  wire [15:0] my_Benes_io_o_dist_bus1_2; // @[FlexDPE.scala 64:26]
  wire [15:0] my_Benes_io_o_dist_bus1_3; // @[FlexDPE.scala 64:26]
  wire [15:0] my_Benes_io_o_dist_bus2_0; // @[FlexDPE.scala 64:26]
  wire [15:0] my_Benes_io_o_dist_bus2_1; // @[FlexDPE.scala 64:26]
  wire [15:0] my_Benes_io_o_dist_bus2_2; // @[FlexDPE.scala 64:26]
  wire [15:0] my_Benes_io_o_dist_bus2_3; // @[FlexDPE.scala 64:26]
  wire [15:0] buffer_mult_io_buffer1_0; // @[FlexDPE.scala 75:30]
  wire [15:0] buffer_mult_io_buffer1_1; // @[FlexDPE.scala 75:30]
  wire [15:0] buffer_mult_io_buffer1_2; // @[FlexDPE.scala 75:30]
  wire [15:0] buffer_mult_io_buffer1_3; // @[FlexDPE.scala 75:30]
  wire [15:0] buffer_mult_io_buffer2_0; // @[FlexDPE.scala 75:30]
  wire [15:0] buffer_mult_io_buffer2_1; // @[FlexDPE.scala 75:30]
  wire [15:0] buffer_mult_io_buffer2_2; // @[FlexDPE.scala 75:30]
  wire [15:0] buffer_mult_io_buffer2_3; // @[FlexDPE.scala 75:30]
  wire [15:0] buffer_mult_io_out_0; // @[FlexDPE.scala 75:30]
  wire [15:0] buffer_mult_io_out_1; // @[FlexDPE.scala 75:30]
  wire [15:0] buffer_mult_io_out_2; // @[FlexDPE.scala 75:30]
  wire [15:0] buffer_mult_io_out_3; // @[FlexDPE.scala 75:30]
  wire  my_fan_network_clock; // @[FlexDPE.scala 87:32]
  wire  my_fan_network_reset; // @[FlexDPE.scala 87:32]
  wire  my_fan_network_io_i_valid; // @[FlexDPE.scala 87:32]
  wire [31:0] my_fan_network_io_i_data_bus_0; // @[FlexDPE.scala 87:32]
  wire [31:0] my_fan_network_io_i_data_bus_1; // @[FlexDPE.scala 87:32]
  wire [31:0] my_fan_network_io_i_data_bus_2; // @[FlexDPE.scala 87:32]
  wire [31:0] my_fan_network_io_i_data_bus_3; // @[FlexDPE.scala 87:32]
  wire  my_fan_network_io_i_add_en_bus_0; // @[FlexDPE.scala 87:32]
  wire  my_fan_network_io_i_add_en_bus_1; // @[FlexDPE.scala 87:32]
  wire  my_fan_network_io_i_add_en_bus_2; // @[FlexDPE.scala 87:32]
  wire [2:0] my_fan_network_io_i_cmd_bus_0; // @[FlexDPE.scala 87:32]
  wire [2:0] my_fan_network_io_i_cmd_bus_1; // @[FlexDPE.scala 87:32]
  wire [2:0] my_fan_network_io_i_cmd_bus_2; // @[FlexDPE.scala 87:32]
  wire [31:0] my_fan_network_io_o_adder_0; // @[FlexDPE.scala 87:32]
  wire [31:0] my_fan_network_io_o_adder_1; // @[FlexDPE.scala 87:32]
  wire [31:0] my_fan_network_io_o_adder_2; // @[FlexDPE.scala 87:32]
  reg [14:0] r_mult_0; // @[FlexDPE.scala 32:26]
  reg [14:0] r_mult_1; // @[FlexDPE.scala 32:26]
  reg [14:0] r_mult_2; // @[FlexDPE.scala 32:26]
  reg [14:0] r_mult_3; // @[FlexDPE.scala 32:26]
  reg [15:0] matrix_0_0; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_0_1; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_0_2; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_0_3; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_0_4; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_0_5; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_0_6; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_0_7; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_1_0; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_1_1; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_1_2; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_1_3; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_1_4; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_1_5; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_1_6; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_1_7; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_2_0; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_2_1; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_2_2; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_2_3; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_2_4; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_2_5; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_2_6; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_2_7; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_3_0; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_3_1; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_3_2; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_3_3; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_3_4; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_3_5; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_3_6; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_3_7; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_4_0; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_4_1; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_4_2; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_4_3; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_4_4; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_4_5; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_4_6; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_4_7; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_5_0; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_5_1; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_5_2; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_5_3; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_5_4; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_5_5; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_5_6; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_5_7; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_6_0; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_6_1; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_6_2; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_6_3; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_6_4; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_6_5; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_6_6; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_6_7; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_7_0; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_7_1; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_7_2; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_7_3; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_7_4; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_7_5; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_7_6; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_7_7; // @[FlexDPE.scala 33:21]
  wire [15:0] _GEN_0 = reset ? 16'h0 : buffer_mult_io_out_0; // @[FlexDPE.scala 32:{26,26} 81:14]
  wire [15:0] _GEN_1 = reset ? 16'h0 : buffer_mult_io_out_1; // @[FlexDPE.scala 32:{26,26} 81:14]
  wire [15:0] _GEN_2 = reset ? 16'h0 : buffer_mult_io_out_2; // @[FlexDPE.scala 32:{26,26} 81:14]
  wire [15:0] _GEN_3 = reset ? 16'h0 : buffer_mult_io_out_3; // @[FlexDPE.scala 32:{26,26} 81:14]
  fancontrol4 my_controller ( // @[FlexDPE.scala 55:31]
    .clock(my_controller_clock),
    .reset(my_controller_reset),
    .io_i_data_valid(my_controller_io_i_data_valid),
    .io_o_reduction_add_0(my_controller_io_o_reduction_add_0),
    .io_o_reduction_add_1(my_controller_io_o_reduction_add_1),
    .io_o_reduction_add_2(my_controller_io_o_reduction_add_2),
    .io_o_reduction_cmd_0(my_controller_io_o_reduction_cmd_0),
    .io_o_reduction_cmd_1(my_controller_io_o_reduction_cmd_1),
    .io_o_reduction_cmd_2(my_controller_io_o_reduction_cmd_2),
    .io_o_reduction_valid(my_controller_io_o_reduction_valid)
  );
  Benes my_Benes ( // @[FlexDPE.scala 64:26]
    .io_i_data_bus2_0(my_Benes_io_i_data_bus2_0),
    .io_i_data_bus2_1(my_Benes_io_i_data_bus2_1),
    .io_i_data_bus2_2(my_Benes_io_i_data_bus2_2),
    .io_i_data_bus2_3(my_Benes_io_i_data_bus2_3),
    .io_i_data_bus1_0(my_Benes_io_i_data_bus1_0),
    .io_i_data_bus1_1(my_Benes_io_i_data_bus1_1),
    .io_i_data_bus1_2(my_Benes_io_i_data_bus1_2),
    .io_i_data_bus1_3(my_Benes_io_i_data_bus1_3),
    .io_i_mux_bus_0(my_Benes_io_i_mux_bus_0),
    .io_i_mux_bus_1(my_Benes_io_i_mux_bus_1),
    .io_i_mux_bus_2(my_Benes_io_i_mux_bus_2),
    .io_i_mux_bus_3(my_Benes_io_i_mux_bus_3),
    .io_o_dist_bus1_0(my_Benes_io_o_dist_bus1_0),
    .io_o_dist_bus1_1(my_Benes_io_o_dist_bus1_1),
    .io_o_dist_bus1_2(my_Benes_io_o_dist_bus1_2),
    .io_o_dist_bus1_3(my_Benes_io_o_dist_bus1_3),
    .io_o_dist_bus2_0(my_Benes_io_o_dist_bus2_0),
    .io_o_dist_bus2_1(my_Benes_io_o_dist_bus2_1),
    .io_o_dist_bus2_2(my_Benes_io_o_dist_bus2_2),
    .io_o_dist_bus2_3(my_Benes_io_o_dist_bus2_3)
  );
  buffer_multiplication buffer_mult ( // @[FlexDPE.scala 75:30]
    .io_buffer1_0(buffer_mult_io_buffer1_0),
    .io_buffer1_1(buffer_mult_io_buffer1_1),
    .io_buffer1_2(buffer_mult_io_buffer1_2),
    .io_buffer1_3(buffer_mult_io_buffer1_3),
    .io_buffer2_0(buffer_mult_io_buffer2_0),
    .io_buffer2_1(buffer_mult_io_buffer2_1),
    .io_buffer2_2(buffer_mult_io_buffer2_2),
    .io_buffer2_3(buffer_mult_io_buffer2_3),
    .io_out_0(buffer_mult_io_out_0),
    .io_out_1(buffer_mult_io_out_1),
    .io_out_2(buffer_mult_io_out_2),
    .io_out_3(buffer_mult_io_out_3)
  );
  Fan4 my_fan_network ( // @[FlexDPE.scala 87:32]
    .clock(my_fan_network_clock),
    .reset(my_fan_network_reset),
    .io_i_valid(my_fan_network_io_i_valid),
    .io_i_data_bus_0(my_fan_network_io_i_data_bus_0),
    .io_i_data_bus_1(my_fan_network_io_i_data_bus_1),
    .io_i_data_bus_2(my_fan_network_io_i_data_bus_2),
    .io_i_data_bus_3(my_fan_network_io_i_data_bus_3),
    .io_i_add_en_bus_0(my_fan_network_io_i_add_en_bus_0),
    .io_i_add_en_bus_1(my_fan_network_io_i_add_en_bus_1),
    .io_i_add_en_bus_2(my_fan_network_io_i_add_en_bus_2),
    .io_i_cmd_bus_0(my_fan_network_io_i_cmd_bus_0),
    .io_i_cmd_bus_1(my_fan_network_io_i_cmd_bus_1),
    .io_i_cmd_bus_2(my_fan_network_io_i_cmd_bus_2),
    .io_o_adder_0(my_fan_network_io_o_adder_0),
    .io_o_adder_1(my_fan_network_io_o_adder_1),
    .io_o_adder_2(my_fan_network_io_o_adder_2)
  );
  assign io_o_adder_0 = my_fan_network_io_o_adder_0[15:0]; // @[FlexDPE.scala 96:16]
  assign io_o_adder_1 = my_fan_network_io_o_adder_1[15:0]; // @[FlexDPE.scala 96:16]
  assign io_o_adder_2 = my_fan_network_io_o_adder_2[15:0]; // @[FlexDPE.scala 96:16]
  assign my_controller_clock = clock;
  assign my_controller_reset = reset;
  assign my_controller_io_i_data_valid = io_i_data_valid; // @[FlexDPE.scala 59:35]
  assign my_Benes_io_i_data_bus2_0 = io_i_data_bus2_0; // @[FlexDPE.scala 67:29]
  assign my_Benes_io_i_data_bus2_1 = io_i_data_bus2_1; // @[FlexDPE.scala 67:29]
  assign my_Benes_io_i_data_bus2_2 = io_i_data_bus2_2; // @[FlexDPE.scala 67:29]
  assign my_Benes_io_i_data_bus2_3 = io_i_data_bus2_3; // @[FlexDPE.scala 67:29]
  assign my_Benes_io_i_data_bus1_0 = io_i_data_bus_0; // @[FlexDPE.scala 66:29]
  assign my_Benes_io_i_data_bus1_1 = io_i_data_bus_1; // @[FlexDPE.scala 66:29]
  assign my_Benes_io_i_data_bus1_2 = io_i_data_bus_2; // @[FlexDPE.scala 66:29]
  assign my_Benes_io_i_data_bus1_3 = io_i_data_bus_3; // @[FlexDPE.scala 66:29]
  assign my_Benes_io_i_mux_bus_0 = io_i_mux_bus_0; // @[FlexDPE.scala 68:27]
  assign my_Benes_io_i_mux_bus_1 = io_i_mux_bus_1; // @[FlexDPE.scala 68:27]
  assign my_Benes_io_i_mux_bus_2 = io_i_mux_bus_2; // @[FlexDPE.scala 68:27]
  assign my_Benes_io_i_mux_bus_3 = io_i_mux_bus_3; // @[FlexDPE.scala 68:27]
  assign buffer_mult_io_buffer1_0 = my_Benes_io_o_dist_bus1_0; // @[FlexDPE.scala 78:30]
  assign buffer_mult_io_buffer1_1 = my_Benes_io_o_dist_bus1_1; // @[FlexDPE.scala 78:30]
  assign buffer_mult_io_buffer1_2 = my_Benes_io_o_dist_bus1_2; // @[FlexDPE.scala 78:30]
  assign buffer_mult_io_buffer1_3 = my_Benes_io_o_dist_bus1_3; // @[FlexDPE.scala 78:30]
  assign buffer_mult_io_buffer2_0 = my_Benes_io_o_dist_bus2_0; // @[FlexDPE.scala 79:30]
  assign buffer_mult_io_buffer2_1 = my_Benes_io_o_dist_bus2_1; // @[FlexDPE.scala 79:30]
  assign buffer_mult_io_buffer2_2 = my_Benes_io_o_dist_bus2_2; // @[FlexDPE.scala 79:30]
  assign buffer_mult_io_buffer2_3 = my_Benes_io_o_dist_bus2_3; // @[FlexDPE.scala 79:30]
  assign my_fan_network_clock = clock;
  assign my_fan_network_reset = reset;
  assign my_fan_network_io_i_valid = my_controller_io_o_reduction_valid; // @[FlexDPE.scala 89:31]
  assign my_fan_network_io_i_data_bus_0 = {{17'd0}, r_mult_0}; // @[FlexDPE.scala 90:34]
  assign my_fan_network_io_i_data_bus_1 = {{17'd0}, r_mult_1}; // @[FlexDPE.scala 90:34]
  assign my_fan_network_io_i_data_bus_2 = {{17'd0}, r_mult_2}; // @[FlexDPE.scala 90:34]
  assign my_fan_network_io_i_data_bus_3 = {{17'd0}, r_mult_3}; // @[FlexDPE.scala 90:34]
  assign my_fan_network_io_i_add_en_bus_0 = my_controller_io_o_reduction_add_0; // @[FlexDPE.scala 91:36]
  assign my_fan_network_io_i_add_en_bus_1 = my_controller_io_o_reduction_add_1; // @[FlexDPE.scala 91:36]
  assign my_fan_network_io_i_add_en_bus_2 = my_controller_io_o_reduction_add_2; // @[FlexDPE.scala 91:36]
  assign my_fan_network_io_i_cmd_bus_0 = my_controller_io_o_reduction_cmd_0; // @[FlexDPE.scala 92:33]
  assign my_fan_network_io_i_cmd_bus_1 = my_controller_io_o_reduction_cmd_1; // @[FlexDPE.scala 92:33]
  assign my_fan_network_io_i_cmd_bus_2 = my_controller_io_o_reduction_cmd_2; // @[FlexDPE.scala 92:33]
  always @(posedge clock) begin
    r_mult_0 <= _GEN_0[14:0]; // @[FlexDPE.scala 32:{26,26} 81:14]
    r_mult_1 <= _GEN_1[14:0]; // @[FlexDPE.scala 32:{26,26} 81:14]
    r_mult_2 <= _GEN_2[14:0]; // @[FlexDPE.scala 32:{26,26} 81:14]
    r_mult_3 <= _GEN_3[14:0]; // @[FlexDPE.scala 32:{26,26} 81:14]
    matrix_0_0 <= matrix_0_0; // @[FlexDPE.scala 33:21]
    matrix_0_1 <= matrix_0_1; // @[FlexDPE.scala 33:21]
    matrix_0_2 <= matrix_0_2; // @[FlexDPE.scala 33:21]
    matrix_0_3 <= matrix_0_3; // @[FlexDPE.scala 33:21]
    matrix_0_4 <= matrix_0_4; // @[FlexDPE.scala 33:21]
    matrix_0_5 <= matrix_0_5; // @[FlexDPE.scala 33:21]
    matrix_0_6 <= matrix_0_6; // @[FlexDPE.scala 33:21]
    matrix_0_7 <= matrix_0_7; // @[FlexDPE.scala 33:21]
    matrix_1_0 <= matrix_1_0; // @[FlexDPE.scala 33:21]
    matrix_1_1 <= matrix_1_1; // @[FlexDPE.scala 33:21]
    matrix_1_2 <= matrix_1_2; // @[FlexDPE.scala 33:21]
    matrix_1_3 <= matrix_1_3; // @[FlexDPE.scala 33:21]
    matrix_1_4 <= matrix_1_4; // @[FlexDPE.scala 33:21]
    matrix_1_5 <= matrix_1_5; // @[FlexDPE.scala 33:21]
    matrix_1_6 <= matrix_1_6; // @[FlexDPE.scala 33:21]
    matrix_1_7 <= matrix_1_7; // @[FlexDPE.scala 33:21]
    matrix_2_0 <= matrix_2_0; // @[FlexDPE.scala 33:21]
    matrix_2_1 <= matrix_2_1; // @[FlexDPE.scala 33:21]
    matrix_2_2 <= matrix_2_2; // @[FlexDPE.scala 33:21]
    matrix_2_3 <= matrix_2_3; // @[FlexDPE.scala 33:21]
    matrix_2_4 <= matrix_2_4; // @[FlexDPE.scala 33:21]
    matrix_2_5 <= matrix_2_5; // @[FlexDPE.scala 33:21]
    matrix_2_6 <= matrix_2_6; // @[FlexDPE.scala 33:21]
    matrix_2_7 <= matrix_2_7; // @[FlexDPE.scala 33:21]
    matrix_3_0 <= matrix_3_0; // @[FlexDPE.scala 33:21]
    matrix_3_1 <= matrix_3_1; // @[FlexDPE.scala 33:21]
    matrix_3_2 <= matrix_3_2; // @[FlexDPE.scala 33:21]
    matrix_3_3 <= matrix_3_3; // @[FlexDPE.scala 33:21]
    matrix_3_4 <= matrix_3_4; // @[FlexDPE.scala 33:21]
    matrix_3_5 <= matrix_3_5; // @[FlexDPE.scala 33:21]
    matrix_3_6 <= matrix_3_6; // @[FlexDPE.scala 33:21]
    matrix_3_7 <= matrix_3_7; // @[FlexDPE.scala 33:21]
    matrix_4_0 <= matrix_4_0; // @[FlexDPE.scala 33:21]
    matrix_4_1 <= matrix_4_1; // @[FlexDPE.scala 33:21]
    matrix_4_2 <= matrix_4_2; // @[FlexDPE.scala 33:21]
    matrix_4_3 <= matrix_4_3; // @[FlexDPE.scala 33:21]
    matrix_4_4 <= matrix_4_4; // @[FlexDPE.scala 33:21]
    matrix_4_5 <= matrix_4_5; // @[FlexDPE.scala 33:21]
    matrix_4_6 <= matrix_4_6; // @[FlexDPE.scala 33:21]
    matrix_4_7 <= matrix_4_7; // @[FlexDPE.scala 33:21]
    matrix_5_0 <= matrix_5_0; // @[FlexDPE.scala 33:21]
    matrix_5_1 <= matrix_5_1; // @[FlexDPE.scala 33:21]
    matrix_5_2 <= matrix_5_2; // @[FlexDPE.scala 33:21]
    matrix_5_3 <= matrix_5_3; // @[FlexDPE.scala 33:21]
    matrix_5_4 <= matrix_5_4; // @[FlexDPE.scala 33:21]
    matrix_5_5 <= matrix_5_5; // @[FlexDPE.scala 33:21]
    matrix_5_6 <= matrix_5_6; // @[FlexDPE.scala 33:21]
    matrix_5_7 <= matrix_5_7; // @[FlexDPE.scala 33:21]
    matrix_6_0 <= matrix_6_0; // @[FlexDPE.scala 33:21]
    matrix_6_1 <= matrix_6_1; // @[FlexDPE.scala 33:21]
    matrix_6_2 <= matrix_6_2; // @[FlexDPE.scala 33:21]
    matrix_6_3 <= matrix_6_3; // @[FlexDPE.scala 33:21]
    matrix_6_4 <= matrix_6_4; // @[FlexDPE.scala 33:21]
    matrix_6_5 <= matrix_6_5; // @[FlexDPE.scala 33:21]
    matrix_6_6 <= matrix_6_6; // @[FlexDPE.scala 33:21]
    matrix_6_7 <= matrix_6_7; // @[FlexDPE.scala 33:21]
    matrix_7_0 <= matrix_7_0; // @[FlexDPE.scala 33:21]
    matrix_7_1 <= matrix_7_1; // @[FlexDPE.scala 33:21]
    matrix_7_2 <= matrix_7_2; // @[FlexDPE.scala 33:21]
    matrix_7_3 <= matrix_7_3; // @[FlexDPE.scala 33:21]
    matrix_7_4 <= matrix_7_4; // @[FlexDPE.scala 33:21]
    matrix_7_5 <= matrix_7_5; // @[FlexDPE.scala 33:21]
    matrix_7_6 <= matrix_7_6; // @[FlexDPE.scala 33:21]
    matrix_7_7 <= matrix_7_7; // @[FlexDPE.scala 33:21]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_mult_0 = _RAND_0[14:0];
  _RAND_1 = {1{`RANDOM}};
  r_mult_1 = _RAND_1[14:0];
  _RAND_2 = {1{`RANDOM}};
  r_mult_2 = _RAND_2[14:0];
  _RAND_3 = {1{`RANDOM}};
  r_mult_3 = _RAND_3[14:0];
  _RAND_4 = {1{`RANDOM}};
  matrix_0_0 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  matrix_0_1 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  matrix_0_2 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  matrix_0_3 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  matrix_0_4 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  matrix_0_5 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  matrix_0_6 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  matrix_0_7 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  matrix_1_0 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  matrix_1_1 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  matrix_1_2 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  matrix_1_3 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  matrix_1_4 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  matrix_1_5 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  matrix_1_6 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  matrix_1_7 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  matrix_2_0 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  matrix_2_1 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  matrix_2_2 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  matrix_2_3 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  matrix_2_4 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  matrix_2_5 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  matrix_2_6 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  matrix_2_7 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  matrix_3_0 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  matrix_3_1 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  matrix_3_2 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  matrix_3_3 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  matrix_3_4 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  matrix_3_5 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  matrix_3_6 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  matrix_3_7 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  matrix_4_0 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  matrix_4_1 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  matrix_4_2 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  matrix_4_3 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  matrix_4_4 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  matrix_4_5 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  matrix_4_6 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  matrix_4_7 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  matrix_5_0 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  matrix_5_1 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  matrix_5_2 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  matrix_5_3 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  matrix_5_4 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  matrix_5_5 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  matrix_5_6 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  matrix_5_7 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  matrix_6_0 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  matrix_6_1 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  matrix_6_2 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  matrix_6_3 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  matrix_6_4 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  matrix_6_5 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  matrix_6_6 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  matrix_6_7 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  matrix_7_0 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  matrix_7_1 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  matrix_7_2 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  matrix_7_3 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  matrix_7_4 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  matrix_7_5 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  matrix_7_6 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  matrix_7_7 = _RAND_67[15:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FlexDPU(
  input         clock,
  input         reset,
  input  [31:0] io_CalFDE,
  input         io_i_stationary,
  input         io_i_data_valid,
  input  [15:0] io_Stationary_matrix_0_0,
  input  [15:0] io_Stationary_matrix_0_1,
  input  [15:0] io_Stationary_matrix_0_2,
  input  [15:0] io_Stationary_matrix_0_3,
  input  [15:0] io_Stationary_matrix_0_4,
  input  [15:0] io_Stationary_matrix_0_5,
  input  [15:0] io_Stationary_matrix_0_6,
  input  [15:0] io_Stationary_matrix_0_7,
  input  [15:0] io_Stationary_matrix_1_0,
  input  [15:0] io_Stationary_matrix_1_1,
  input  [15:0] io_Stationary_matrix_1_2,
  input  [15:0] io_Stationary_matrix_1_3,
  input  [15:0] io_Stationary_matrix_1_4,
  input  [15:0] io_Stationary_matrix_1_5,
  input  [15:0] io_Stationary_matrix_1_6,
  input  [15:0] io_Stationary_matrix_1_7,
  input  [15:0] io_Stationary_matrix_2_0,
  input  [15:0] io_Stationary_matrix_2_1,
  input  [15:0] io_Stationary_matrix_2_2,
  input  [15:0] io_Stationary_matrix_2_3,
  input  [15:0] io_Stationary_matrix_2_4,
  input  [15:0] io_Stationary_matrix_2_5,
  input  [15:0] io_Stationary_matrix_2_6,
  input  [15:0] io_Stationary_matrix_2_7,
  input  [15:0] io_Stationary_matrix_3_0,
  input  [15:0] io_Stationary_matrix_3_1,
  input  [15:0] io_Stationary_matrix_3_2,
  input  [15:0] io_Stationary_matrix_3_3,
  input  [15:0] io_Stationary_matrix_3_4,
  input  [15:0] io_Stationary_matrix_3_5,
  input  [15:0] io_Stationary_matrix_3_6,
  input  [15:0] io_Stationary_matrix_3_7,
  input  [15:0] io_Stationary_matrix_4_0,
  input  [15:0] io_Stationary_matrix_4_1,
  input  [15:0] io_Stationary_matrix_4_2,
  input  [15:0] io_Stationary_matrix_4_3,
  input  [15:0] io_Stationary_matrix_4_4,
  input  [15:0] io_Stationary_matrix_4_5,
  input  [15:0] io_Stationary_matrix_4_6,
  input  [15:0] io_Stationary_matrix_4_7,
  input  [15:0] io_Stationary_matrix_5_0,
  input  [15:0] io_Stationary_matrix_5_1,
  input  [15:0] io_Stationary_matrix_5_2,
  input  [15:0] io_Stationary_matrix_5_3,
  input  [15:0] io_Stationary_matrix_5_4,
  input  [15:0] io_Stationary_matrix_5_5,
  input  [15:0] io_Stationary_matrix_5_6,
  input  [15:0] io_Stationary_matrix_5_7,
  input  [15:0] io_Stationary_matrix_6_0,
  input  [15:0] io_Stationary_matrix_6_1,
  input  [15:0] io_Stationary_matrix_6_2,
  input  [15:0] io_Stationary_matrix_6_3,
  input  [15:0] io_Stationary_matrix_6_4,
  input  [15:0] io_Stationary_matrix_6_5,
  input  [15:0] io_Stationary_matrix_6_6,
  input  [15:0] io_Stationary_matrix_6_7,
  input  [15:0] io_Stationary_matrix_7_0,
  input  [15:0] io_Stationary_matrix_7_1,
  input  [15:0] io_Stationary_matrix_7_2,
  input  [15:0] io_Stationary_matrix_7_3,
  input  [15:0] io_Stationary_matrix_7_4,
  input  [15:0] io_Stationary_matrix_7_5,
  input  [15:0] io_Stationary_matrix_7_6,
  input  [15:0] io_Stationary_matrix_7_7,
  input  [15:0] io_Streaming_matrix_0_0,
  input  [15:0] io_Streaming_matrix_0_1,
  input  [15:0] io_Streaming_matrix_0_2,
  input  [15:0] io_Streaming_matrix_0_3,
  input  [15:0] io_Streaming_matrix_0_4,
  input  [15:0] io_Streaming_matrix_0_5,
  input  [15:0] io_Streaming_matrix_0_6,
  input  [15:0] io_Streaming_matrix_0_7,
  input  [15:0] io_Streaming_matrix_1_0,
  input  [15:0] io_Streaming_matrix_1_1,
  input  [15:0] io_Streaming_matrix_1_2,
  input  [15:0] io_Streaming_matrix_1_3,
  input  [15:0] io_Streaming_matrix_1_4,
  input  [15:0] io_Streaming_matrix_1_5,
  input  [15:0] io_Streaming_matrix_1_6,
  input  [15:0] io_Streaming_matrix_1_7,
  input  [15:0] io_Streaming_matrix_2_0,
  input  [15:0] io_Streaming_matrix_2_1,
  input  [15:0] io_Streaming_matrix_2_2,
  input  [15:0] io_Streaming_matrix_2_3,
  input  [15:0] io_Streaming_matrix_2_4,
  input  [15:0] io_Streaming_matrix_2_5,
  input  [15:0] io_Streaming_matrix_2_6,
  input  [15:0] io_Streaming_matrix_2_7,
  input  [15:0] io_Streaming_matrix_3_0,
  input  [15:0] io_Streaming_matrix_3_1,
  input  [15:0] io_Streaming_matrix_3_2,
  input  [15:0] io_Streaming_matrix_3_3,
  input  [15:0] io_Streaming_matrix_3_4,
  input  [15:0] io_Streaming_matrix_3_5,
  input  [15:0] io_Streaming_matrix_3_6,
  input  [15:0] io_Streaming_matrix_3_7,
  input  [15:0] io_Streaming_matrix_4_0,
  input  [15:0] io_Streaming_matrix_4_1,
  input  [15:0] io_Streaming_matrix_4_2,
  input  [15:0] io_Streaming_matrix_4_3,
  input  [15:0] io_Streaming_matrix_4_4,
  input  [15:0] io_Streaming_matrix_4_5,
  input  [15:0] io_Streaming_matrix_4_6,
  input  [15:0] io_Streaming_matrix_4_7,
  input  [15:0] io_Streaming_matrix_5_0,
  input  [15:0] io_Streaming_matrix_5_1,
  input  [15:0] io_Streaming_matrix_5_2,
  input  [15:0] io_Streaming_matrix_5_3,
  input  [15:0] io_Streaming_matrix_5_4,
  input  [15:0] io_Streaming_matrix_5_5,
  input  [15:0] io_Streaming_matrix_5_6,
  input  [15:0] io_Streaming_matrix_5_7,
  input  [15:0] io_Streaming_matrix_6_0,
  input  [15:0] io_Streaming_matrix_6_1,
  input  [15:0] io_Streaming_matrix_6_2,
  input  [15:0] io_Streaming_matrix_6_3,
  input  [15:0] io_Streaming_matrix_6_4,
  input  [15:0] io_Streaming_matrix_6_5,
  input  [15:0] io_Streaming_matrix_6_6,
  input  [15:0] io_Streaming_matrix_6_7,
  input  [15:0] io_Streaming_matrix_7_0,
  input  [15:0] io_Streaming_matrix_7_1,
  input  [15:0] io_Streaming_matrix_7_2,
  input  [15:0] io_Streaming_matrix_7_3,
  input  [15:0] io_Streaming_matrix_7_4,
  input  [15:0] io_Streaming_matrix_7_5,
  input  [15:0] io_Streaming_matrix_7_6,
  input  [15:0] io_Streaming_matrix_7_7,
  output [15:0] io_output_0_0,
  output [15:0] io_output_0_1,
  output [15:0] io_output_0_2,
  output [15:0] io_output_0_3,
  output [15:0] io_output_0_4,
  output [15:0] io_output_0_5,
  output [15:0] io_output_0_6,
  output [15:0] io_output_0_7,
  output [15:0] io_output_1_0,
  output [15:0] io_output_1_1,
  output [15:0] io_output_1_2,
  output [15:0] io_output_1_3,
  output [15:0] io_output_1_4,
  output [15:0] io_output_1_5,
  output [15:0] io_output_1_6,
  output [15:0] io_output_1_7,
  output [15:0] io_output_2_0,
  output [15:0] io_output_2_1,
  output [15:0] io_output_2_2,
  output [15:0] io_output_2_3,
  output [15:0] io_output_2_4,
  output [15:0] io_output_2_5,
  output [15:0] io_output_2_6,
  output [15:0] io_output_2_7,
  output [15:0] io_output_3_0,
  output [15:0] io_output_3_1,
  output [15:0] io_output_3_2,
  output [15:0] io_output_3_3,
  output [15:0] io_output_3_4,
  output [15:0] io_output_3_5,
  output [15:0] io_output_3_6,
  output [15:0] io_output_3_7,
  output [15:0] io_output_4_0,
  output [15:0] io_output_4_1,
  output [15:0] io_output_4_2,
  output [15:0] io_output_4_3,
  output [15:0] io_output_4_4,
  output [15:0] io_output_4_5,
  output [15:0] io_output_4_6,
  output [15:0] io_output_4_7,
  output [15:0] io_output_5_0,
  output [15:0] io_output_5_1,
  output [15:0] io_output_5_2,
  output [15:0] io_output_5_3,
  output [15:0] io_output_5_4,
  output [15:0] io_output_5_5,
  output [15:0] io_output_5_6,
  output [15:0] io_output_5_7,
  output [15:0] io_output_6_0,
  output [15:0] io_output_6_1,
  output [15:0] io_output_6_2,
  output [15:0] io_output_6_3,
  output [15:0] io_output_6_4,
  output [15:0] io_output_6_5,
  output [15:0] io_output_6_6,
  output [15:0] io_output_6_7,
  output [15:0] io_output_7_0,
  output [15:0] io_output_7_1,
  output [15:0] io_output_7_2,
  output [15:0] io_output_7_3,
  output [15:0] io_output_7_4,
  output [15:0] io_output_7_5,
  output [15:0] io_output_7_6,
  output [15:0] io_output_7_7
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
`endif // RANDOMIZE_REG_INIT
  wire  PathFinder_clock; // @[FlexDPU.scala 77:41]
  wire  PathFinder_reset; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_0_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_0_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_0_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_0_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_0_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_0_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_0_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_0_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_1_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_1_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_1_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_1_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_1_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_1_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_1_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_1_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_2_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_2_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_2_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_2_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_2_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_2_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_2_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_2_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_3_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_3_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_3_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_3_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_3_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_3_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_3_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_3_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_4_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_4_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_4_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_4_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_4_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_4_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_4_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_4_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_5_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_5_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_5_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_5_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_5_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_5_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_5_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_5_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_6_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_6_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_6_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_6_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_6_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_6_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_6_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_6_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_7_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_7_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_7_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_7_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_7_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_7_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_7_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_7_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Streaming_matrix_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Streaming_matrix_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Streaming_matrix_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Streaming_matrix_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Streaming_matrix_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Streaming_matrix_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Streaming_matrix_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Streaming_matrix_7; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_io_i_mux_bus_0; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_io_i_mux_bus_1; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_io_i_mux_bus_2; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_io_i_mux_bus_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Source_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Source_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Source_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Source_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_destination_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_destination_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_destination_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_destination_3; // @[FlexDPU.scala 77:41]
  wire  PathFinder_io_PF_Valid; // @[FlexDPU.scala 77:41]
  wire [31:0] PathFinder_io_NoDPE; // @[FlexDPU.scala 77:41]
  wire  PathFinder_io_DataValid; // @[FlexDPU.scala 77:41]
  wire  PathFinder_1_clock; // @[FlexDPU.scala 77:41]
  wire  PathFinder_1_reset; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_0_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_0_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_0_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_0_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_0_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_0_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_0_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_0_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_1_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_1_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_1_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_1_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_1_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_1_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_1_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_1_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_2_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_2_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_2_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_2_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_2_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_2_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_2_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_2_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_3_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_3_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_3_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_3_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_3_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_3_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_3_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_3_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_4_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_4_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_4_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_4_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_4_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_4_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_4_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_4_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_5_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_5_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_5_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_5_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_5_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_5_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_5_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_5_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_6_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_6_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_6_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_6_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_6_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_6_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_6_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_6_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_7_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_7_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_7_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_7_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_7_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_7_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_7_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_7_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Streaming_matrix_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Streaming_matrix_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Streaming_matrix_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Streaming_matrix_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Streaming_matrix_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Streaming_matrix_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Streaming_matrix_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Streaming_matrix_7; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_1_io_i_mux_bus_0; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_1_io_i_mux_bus_1; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_1_io_i_mux_bus_2; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_1_io_i_mux_bus_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Source_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Source_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Source_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Source_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_destination_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_destination_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_destination_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_destination_3; // @[FlexDPU.scala 77:41]
  wire  PathFinder_1_io_PF_Valid; // @[FlexDPU.scala 77:41]
  wire [31:0] PathFinder_1_io_NoDPE; // @[FlexDPU.scala 77:41]
  wire  PathFinder_1_io_DataValid; // @[FlexDPU.scala 77:41]
  wire  PathFinder_2_clock; // @[FlexDPU.scala 77:41]
  wire  PathFinder_2_reset; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_0_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_0_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_0_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_0_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_0_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_0_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_0_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_0_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_1_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_1_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_1_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_1_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_1_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_1_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_1_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_1_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_2_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_2_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_2_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_2_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_2_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_2_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_2_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_2_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_3_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_3_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_3_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_3_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_3_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_3_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_3_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_3_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_4_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_4_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_4_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_4_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_4_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_4_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_4_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_4_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_5_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_5_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_5_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_5_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_5_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_5_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_5_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_5_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_6_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_6_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_6_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_6_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_6_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_6_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_6_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_6_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_7_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_7_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_7_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_7_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_7_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_7_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_7_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_7_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Streaming_matrix_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Streaming_matrix_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Streaming_matrix_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Streaming_matrix_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Streaming_matrix_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Streaming_matrix_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Streaming_matrix_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Streaming_matrix_7; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_2_io_i_mux_bus_0; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_2_io_i_mux_bus_1; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_2_io_i_mux_bus_2; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_2_io_i_mux_bus_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Source_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Source_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Source_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Source_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_destination_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_destination_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_destination_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_destination_3; // @[FlexDPU.scala 77:41]
  wire  PathFinder_2_io_PF_Valid; // @[FlexDPU.scala 77:41]
  wire [31:0] PathFinder_2_io_NoDPE; // @[FlexDPU.scala 77:41]
  wire  PathFinder_2_io_DataValid; // @[FlexDPU.scala 77:41]
  wire  PathFinder_3_clock; // @[FlexDPU.scala 77:41]
  wire  PathFinder_3_reset; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_0_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_0_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_0_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_0_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_0_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_0_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_0_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_0_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_1_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_1_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_1_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_1_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_1_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_1_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_1_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_1_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_2_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_2_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_2_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_2_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_2_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_2_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_2_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_2_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_3_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_3_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_3_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_3_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_3_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_3_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_3_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_3_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_4_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_4_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_4_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_4_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_4_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_4_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_4_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_4_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_5_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_5_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_5_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_5_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_5_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_5_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_5_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_5_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_6_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_6_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_6_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_6_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_6_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_6_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_6_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_6_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_7_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_7_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_7_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_7_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_7_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_7_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_7_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_7_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Streaming_matrix_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Streaming_matrix_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Streaming_matrix_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Streaming_matrix_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Streaming_matrix_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Streaming_matrix_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Streaming_matrix_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Streaming_matrix_7; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_3_io_i_mux_bus_0; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_3_io_i_mux_bus_1; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_3_io_i_mux_bus_2; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_3_io_i_mux_bus_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Source_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Source_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Source_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Source_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_destination_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_destination_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_destination_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_destination_3; // @[FlexDPU.scala 77:41]
  wire  PathFinder_3_io_PF_Valid; // @[FlexDPU.scala 77:41]
  wire [31:0] PathFinder_3_io_NoDPE; // @[FlexDPU.scala 77:41]
  wire  PathFinder_3_io_DataValid; // @[FlexDPU.scala 77:41]
  wire  PathFinder_4_clock; // @[FlexDPU.scala 77:41]
  wire  PathFinder_4_reset; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_0_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_0_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_0_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_0_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_0_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_0_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_0_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_0_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_1_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_1_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_1_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_1_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_1_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_1_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_1_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_1_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_2_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_2_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_2_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_2_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_2_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_2_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_2_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_2_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_3_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_3_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_3_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_3_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_3_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_3_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_3_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_3_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_4_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_4_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_4_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_4_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_4_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_4_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_4_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_4_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_5_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_5_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_5_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_5_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_5_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_5_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_5_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_5_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_6_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_6_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_6_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_6_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_6_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_6_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_6_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_6_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_7_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_7_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_7_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_7_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_7_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_7_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_7_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_7_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Streaming_matrix_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Streaming_matrix_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Streaming_matrix_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Streaming_matrix_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Streaming_matrix_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Streaming_matrix_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Streaming_matrix_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Streaming_matrix_7; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_4_io_i_mux_bus_0; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_4_io_i_mux_bus_1; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_4_io_i_mux_bus_2; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_4_io_i_mux_bus_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Source_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Source_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Source_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Source_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_destination_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_destination_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_destination_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_destination_3; // @[FlexDPU.scala 77:41]
  wire  PathFinder_4_io_PF_Valid; // @[FlexDPU.scala 77:41]
  wire [31:0] PathFinder_4_io_NoDPE; // @[FlexDPU.scala 77:41]
  wire  PathFinder_4_io_DataValid; // @[FlexDPU.scala 77:41]
  wire  PathFinder_5_clock; // @[FlexDPU.scala 77:41]
  wire  PathFinder_5_reset; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_0_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_0_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_0_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_0_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_0_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_0_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_0_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_0_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_1_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_1_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_1_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_1_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_1_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_1_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_1_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_1_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_2_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_2_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_2_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_2_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_2_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_2_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_2_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_2_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_3_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_3_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_3_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_3_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_3_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_3_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_3_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_3_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_4_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_4_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_4_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_4_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_4_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_4_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_4_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_4_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_5_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_5_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_5_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_5_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_5_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_5_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_5_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_5_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_6_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_6_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_6_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_6_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_6_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_6_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_6_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_6_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_7_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_7_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_7_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_7_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_7_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_7_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_7_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_7_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Streaming_matrix_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Streaming_matrix_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Streaming_matrix_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Streaming_matrix_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Streaming_matrix_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Streaming_matrix_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Streaming_matrix_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Streaming_matrix_7; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_5_io_i_mux_bus_0; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_5_io_i_mux_bus_1; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_5_io_i_mux_bus_2; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_5_io_i_mux_bus_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Source_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Source_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Source_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Source_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_destination_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_destination_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_destination_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_destination_3; // @[FlexDPU.scala 77:41]
  wire  PathFinder_5_io_PF_Valid; // @[FlexDPU.scala 77:41]
  wire [31:0] PathFinder_5_io_NoDPE; // @[FlexDPU.scala 77:41]
  wire  PathFinder_5_io_DataValid; // @[FlexDPU.scala 77:41]
  wire  PathFinder_6_clock; // @[FlexDPU.scala 77:41]
  wire  PathFinder_6_reset; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_0_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_0_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_0_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_0_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_0_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_0_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_0_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_0_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_1_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_1_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_1_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_1_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_1_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_1_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_1_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_1_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_2_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_2_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_2_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_2_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_2_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_2_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_2_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_2_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_3_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_3_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_3_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_3_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_3_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_3_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_3_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_3_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_4_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_4_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_4_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_4_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_4_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_4_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_4_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_4_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_5_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_5_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_5_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_5_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_5_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_5_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_5_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_5_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_6_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_6_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_6_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_6_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_6_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_6_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_6_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_6_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_7_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_7_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_7_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_7_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_7_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_7_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_7_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_7_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Streaming_matrix_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Streaming_matrix_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Streaming_matrix_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Streaming_matrix_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Streaming_matrix_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Streaming_matrix_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Streaming_matrix_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Streaming_matrix_7; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_6_io_i_mux_bus_0; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_6_io_i_mux_bus_1; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_6_io_i_mux_bus_2; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_6_io_i_mux_bus_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Source_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Source_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Source_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Source_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_destination_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_destination_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_destination_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_destination_3; // @[FlexDPU.scala 77:41]
  wire  PathFinder_6_io_PF_Valid; // @[FlexDPU.scala 77:41]
  wire [31:0] PathFinder_6_io_NoDPE; // @[FlexDPU.scala 77:41]
  wire  PathFinder_6_io_DataValid; // @[FlexDPU.scala 77:41]
  wire  PathFinder_7_clock; // @[FlexDPU.scala 77:41]
  wire  PathFinder_7_reset; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_0_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_0_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_0_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_0_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_0_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_0_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_0_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_0_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_1_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_1_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_1_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_1_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_1_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_1_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_1_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_1_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_2_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_2_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_2_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_2_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_2_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_2_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_2_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_2_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_3_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_3_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_3_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_3_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_3_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_3_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_3_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_3_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_4_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_4_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_4_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_4_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_4_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_4_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_4_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_4_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_5_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_5_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_5_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_5_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_5_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_5_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_5_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_5_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_6_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_6_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_6_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_6_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_6_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_6_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_6_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_6_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_7_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_7_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_7_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_7_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_7_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_7_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_7_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_7_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Streaming_matrix_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Streaming_matrix_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Streaming_matrix_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Streaming_matrix_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Streaming_matrix_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Streaming_matrix_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Streaming_matrix_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Streaming_matrix_7; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_7_io_i_mux_bus_0; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_7_io_i_mux_bus_1; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_7_io_i_mux_bus_2; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_7_io_i_mux_bus_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Source_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Source_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Source_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Source_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_destination_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_destination_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_destination_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_destination_3; // @[FlexDPU.scala 77:41]
  wire  PathFinder_7_io_PF_Valid; // @[FlexDPU.scala 77:41]
  wire [31:0] PathFinder_7_io_NoDPE; // @[FlexDPU.scala 77:41]
  wire  PathFinder_7_io_DataValid; // @[FlexDPU.scala 77:41]
  wire  PathFinder_8_clock; // @[FlexDPU.scala 77:41]
  wire  PathFinder_8_reset; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_0_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_0_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_0_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_0_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_0_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_0_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_0_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_0_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_1_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_1_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_1_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_1_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_1_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_1_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_1_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_1_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_2_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_2_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_2_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_2_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_2_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_2_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_2_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_2_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_3_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_3_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_3_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_3_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_3_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_3_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_3_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_3_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_4_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_4_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_4_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_4_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_4_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_4_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_4_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_4_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_5_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_5_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_5_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_5_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_5_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_5_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_5_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_5_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_6_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_6_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_6_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_6_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_6_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_6_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_6_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_6_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_7_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_7_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_7_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_7_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_7_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_7_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_7_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_7_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Streaming_matrix_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Streaming_matrix_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Streaming_matrix_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Streaming_matrix_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Streaming_matrix_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Streaming_matrix_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Streaming_matrix_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Streaming_matrix_7; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_8_io_i_mux_bus_0; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_8_io_i_mux_bus_1; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_8_io_i_mux_bus_2; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_8_io_i_mux_bus_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Source_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Source_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Source_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Source_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_destination_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_destination_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_destination_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_destination_3; // @[FlexDPU.scala 77:41]
  wire  PathFinder_8_io_PF_Valid; // @[FlexDPU.scala 77:41]
  wire [31:0] PathFinder_8_io_NoDPE; // @[FlexDPU.scala 77:41]
  wire  PathFinder_8_io_DataValid; // @[FlexDPU.scala 77:41]
  wire  PathFinder_9_clock; // @[FlexDPU.scala 77:41]
  wire  PathFinder_9_reset; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_0_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_0_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_0_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_0_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_0_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_0_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_0_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_0_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_1_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_1_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_1_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_1_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_1_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_1_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_1_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_1_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_2_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_2_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_2_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_2_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_2_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_2_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_2_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_2_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_3_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_3_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_3_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_3_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_3_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_3_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_3_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_3_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_4_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_4_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_4_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_4_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_4_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_4_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_4_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_4_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_5_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_5_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_5_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_5_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_5_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_5_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_5_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_5_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_6_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_6_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_6_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_6_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_6_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_6_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_6_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_6_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_7_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_7_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_7_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_7_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_7_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_7_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_7_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_7_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Streaming_matrix_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Streaming_matrix_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Streaming_matrix_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Streaming_matrix_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Streaming_matrix_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Streaming_matrix_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Streaming_matrix_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Streaming_matrix_7; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_9_io_i_mux_bus_0; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_9_io_i_mux_bus_1; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_9_io_i_mux_bus_2; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_9_io_i_mux_bus_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Source_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Source_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Source_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Source_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_destination_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_destination_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_destination_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_destination_3; // @[FlexDPU.scala 77:41]
  wire  PathFinder_9_io_PF_Valid; // @[FlexDPU.scala 77:41]
  wire [31:0] PathFinder_9_io_NoDPE; // @[FlexDPU.scala 77:41]
  wire  PathFinder_9_io_DataValid; // @[FlexDPU.scala 77:41]
  wire  PathFinder_10_clock; // @[FlexDPU.scala 77:41]
  wire  PathFinder_10_reset; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_0_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_0_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_0_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_0_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_0_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_0_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_0_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_0_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_1_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_1_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_1_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_1_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_1_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_1_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_1_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_1_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_2_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_2_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_2_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_2_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_2_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_2_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_2_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_2_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_3_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_3_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_3_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_3_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_3_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_3_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_3_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_3_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_4_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_4_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_4_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_4_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_4_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_4_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_4_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_4_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_5_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_5_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_5_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_5_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_5_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_5_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_5_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_5_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_6_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_6_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_6_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_6_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_6_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_6_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_6_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_6_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_7_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_7_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_7_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_7_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_7_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_7_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_7_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_7_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Streaming_matrix_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Streaming_matrix_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Streaming_matrix_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Streaming_matrix_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Streaming_matrix_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Streaming_matrix_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Streaming_matrix_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Streaming_matrix_7; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_10_io_i_mux_bus_0; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_10_io_i_mux_bus_1; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_10_io_i_mux_bus_2; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_10_io_i_mux_bus_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Source_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Source_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Source_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Source_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_destination_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_destination_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_destination_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_destination_3; // @[FlexDPU.scala 77:41]
  wire  PathFinder_10_io_PF_Valid; // @[FlexDPU.scala 77:41]
  wire [31:0] PathFinder_10_io_NoDPE; // @[FlexDPU.scala 77:41]
  wire  PathFinder_10_io_DataValid; // @[FlexDPU.scala 77:41]
  wire  PathFinder_11_clock; // @[FlexDPU.scala 77:41]
  wire  PathFinder_11_reset; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_0_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_0_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_0_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_0_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_0_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_0_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_0_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_0_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_1_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_1_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_1_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_1_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_1_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_1_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_1_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_1_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_2_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_2_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_2_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_2_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_2_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_2_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_2_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_2_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_3_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_3_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_3_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_3_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_3_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_3_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_3_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_3_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_4_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_4_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_4_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_4_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_4_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_4_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_4_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_4_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_5_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_5_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_5_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_5_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_5_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_5_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_5_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_5_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_6_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_6_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_6_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_6_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_6_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_6_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_6_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_6_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_7_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_7_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_7_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_7_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_7_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_7_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_7_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_7_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Streaming_matrix_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Streaming_matrix_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Streaming_matrix_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Streaming_matrix_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Streaming_matrix_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Streaming_matrix_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Streaming_matrix_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Streaming_matrix_7; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_11_io_i_mux_bus_0; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_11_io_i_mux_bus_1; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_11_io_i_mux_bus_2; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_11_io_i_mux_bus_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Source_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Source_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Source_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Source_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_destination_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_destination_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_destination_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_destination_3; // @[FlexDPU.scala 77:41]
  wire  PathFinder_11_io_PF_Valid; // @[FlexDPU.scala 77:41]
  wire [31:0] PathFinder_11_io_NoDPE; // @[FlexDPU.scala 77:41]
  wire  PathFinder_11_io_DataValid; // @[FlexDPU.scala 77:41]
  wire  PathFinder_12_clock; // @[FlexDPU.scala 77:41]
  wire  PathFinder_12_reset; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_0_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_0_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_0_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_0_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_0_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_0_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_0_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_0_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_1_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_1_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_1_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_1_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_1_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_1_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_1_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_1_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_2_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_2_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_2_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_2_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_2_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_2_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_2_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_2_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_3_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_3_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_3_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_3_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_3_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_3_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_3_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_3_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_4_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_4_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_4_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_4_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_4_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_4_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_4_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_4_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_5_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_5_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_5_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_5_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_5_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_5_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_5_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_5_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_6_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_6_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_6_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_6_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_6_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_6_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_6_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_6_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_7_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_7_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_7_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_7_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_7_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_7_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_7_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_7_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Streaming_matrix_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Streaming_matrix_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Streaming_matrix_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Streaming_matrix_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Streaming_matrix_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Streaming_matrix_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Streaming_matrix_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Streaming_matrix_7; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_12_io_i_mux_bus_0; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_12_io_i_mux_bus_1; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_12_io_i_mux_bus_2; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_12_io_i_mux_bus_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Source_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Source_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Source_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Source_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_destination_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_destination_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_destination_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_destination_3; // @[FlexDPU.scala 77:41]
  wire  PathFinder_12_io_PF_Valid; // @[FlexDPU.scala 77:41]
  wire [31:0] PathFinder_12_io_NoDPE; // @[FlexDPU.scala 77:41]
  wire  PathFinder_12_io_DataValid; // @[FlexDPU.scala 77:41]
  wire  PathFinder_13_clock; // @[FlexDPU.scala 77:41]
  wire  PathFinder_13_reset; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_0_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_0_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_0_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_0_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_0_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_0_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_0_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_0_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_1_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_1_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_1_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_1_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_1_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_1_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_1_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_1_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_2_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_2_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_2_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_2_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_2_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_2_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_2_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_2_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_3_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_3_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_3_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_3_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_3_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_3_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_3_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_3_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_4_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_4_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_4_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_4_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_4_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_4_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_4_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_4_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_5_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_5_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_5_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_5_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_5_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_5_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_5_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_5_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_6_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_6_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_6_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_6_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_6_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_6_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_6_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_6_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_7_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_7_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_7_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_7_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_7_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_7_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_7_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_7_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Streaming_matrix_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Streaming_matrix_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Streaming_matrix_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Streaming_matrix_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Streaming_matrix_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Streaming_matrix_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Streaming_matrix_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Streaming_matrix_7; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_13_io_i_mux_bus_0; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_13_io_i_mux_bus_1; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_13_io_i_mux_bus_2; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_13_io_i_mux_bus_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Source_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Source_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Source_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Source_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_destination_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_destination_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_destination_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_destination_3; // @[FlexDPU.scala 77:41]
  wire  PathFinder_13_io_PF_Valid; // @[FlexDPU.scala 77:41]
  wire [31:0] PathFinder_13_io_NoDPE; // @[FlexDPU.scala 77:41]
  wire  PathFinder_13_io_DataValid; // @[FlexDPU.scala 77:41]
  wire  PathFinder_14_clock; // @[FlexDPU.scala 77:41]
  wire  PathFinder_14_reset; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_0_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_0_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_0_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_0_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_0_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_0_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_0_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_0_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_1_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_1_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_1_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_1_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_1_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_1_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_1_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_1_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_2_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_2_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_2_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_2_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_2_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_2_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_2_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_2_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_3_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_3_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_3_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_3_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_3_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_3_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_3_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_3_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_4_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_4_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_4_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_4_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_4_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_4_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_4_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_4_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_5_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_5_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_5_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_5_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_5_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_5_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_5_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_5_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_6_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_6_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_6_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_6_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_6_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_6_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_6_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_6_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_7_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_7_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_7_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_7_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_7_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_7_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_7_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_7_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Streaming_matrix_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Streaming_matrix_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Streaming_matrix_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Streaming_matrix_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Streaming_matrix_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Streaming_matrix_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Streaming_matrix_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Streaming_matrix_7; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_14_io_i_mux_bus_0; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_14_io_i_mux_bus_1; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_14_io_i_mux_bus_2; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_14_io_i_mux_bus_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Source_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Source_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Source_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Source_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_destination_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_destination_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_destination_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_destination_3; // @[FlexDPU.scala 77:41]
  wire  PathFinder_14_io_PF_Valid; // @[FlexDPU.scala 77:41]
  wire [31:0] PathFinder_14_io_NoDPE; // @[FlexDPU.scala 77:41]
  wire  PathFinder_14_io_DataValid; // @[FlexDPU.scala 77:41]
  wire  PathFinder_15_clock; // @[FlexDPU.scala 77:41]
  wire  PathFinder_15_reset; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_0_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_0_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_0_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_0_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_0_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_0_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_0_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_0_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_1_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_1_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_1_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_1_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_1_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_1_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_1_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_1_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_2_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_2_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_2_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_2_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_2_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_2_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_2_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_2_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_3_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_3_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_3_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_3_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_3_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_3_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_3_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_3_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_4_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_4_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_4_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_4_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_4_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_4_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_4_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_4_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_5_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_5_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_5_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_5_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_5_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_5_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_5_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_5_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_6_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_6_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_6_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_6_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_6_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_6_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_6_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_6_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_7_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_7_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_7_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_7_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_7_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_7_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_7_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_7_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Streaming_matrix_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Streaming_matrix_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Streaming_matrix_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Streaming_matrix_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Streaming_matrix_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Streaming_matrix_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Streaming_matrix_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Streaming_matrix_7; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_15_io_i_mux_bus_0; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_15_io_i_mux_bus_1; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_15_io_i_mux_bus_2; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_15_io_i_mux_bus_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Source_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Source_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Source_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Source_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_destination_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_destination_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_destination_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_destination_3; // @[FlexDPU.scala 77:41]
  wire  PathFinder_15_io_PF_Valid; // @[FlexDPU.scala 77:41]
  wire [31:0] PathFinder_15_io_NoDPE; // @[FlexDPU.scala 77:41]
  wire  PathFinder_15_io_DataValid; // @[FlexDPU.scala 77:41]
  wire  flexdpecom4_clock; // @[FlexDPU.scala 110:47]
  wire  flexdpecom4_reset; // @[FlexDPU.scala 110:47]
  wire  flexdpecom4_io_i_data_valid; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_io_i_data_bus_0; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_io_i_data_bus_1; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_io_i_data_bus_2; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_io_i_data_bus_3; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_io_i_data_bus2_0; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_io_i_data_bus2_1; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_io_i_data_bus2_2; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_io_i_data_bus2_3; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_io_o_adder_0; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_io_o_adder_1; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_io_o_adder_2; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_io_i_mux_bus_0; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_io_i_mux_bus_1; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_io_i_mux_bus_2; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_io_i_mux_bus_3; // @[FlexDPU.scala 110:47]
  wire  flexdpecom4_1_clock; // @[FlexDPU.scala 110:47]
  wire  flexdpecom4_1_reset; // @[FlexDPU.scala 110:47]
  wire  flexdpecom4_1_io_i_data_valid; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_1_io_i_data_bus_0; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_1_io_i_data_bus_1; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_1_io_i_data_bus_2; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_1_io_i_data_bus_3; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_1_io_i_data_bus2_0; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_1_io_i_data_bus2_1; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_1_io_i_data_bus2_2; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_1_io_i_data_bus2_3; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_1_io_o_adder_0; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_1_io_o_adder_1; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_1_io_o_adder_2; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_1_io_i_mux_bus_0; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_1_io_i_mux_bus_1; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_1_io_i_mux_bus_2; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_1_io_i_mux_bus_3; // @[FlexDPU.scala 110:47]
  wire  flexdpecom4_2_clock; // @[FlexDPU.scala 110:47]
  wire  flexdpecom4_2_reset; // @[FlexDPU.scala 110:47]
  wire  flexdpecom4_2_io_i_data_valid; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_2_io_i_data_bus_0; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_2_io_i_data_bus_1; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_2_io_i_data_bus_2; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_2_io_i_data_bus_3; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_2_io_i_data_bus2_0; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_2_io_i_data_bus2_1; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_2_io_i_data_bus2_2; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_2_io_i_data_bus2_3; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_2_io_o_adder_0; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_2_io_o_adder_1; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_2_io_o_adder_2; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_2_io_i_mux_bus_0; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_2_io_i_mux_bus_1; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_2_io_i_mux_bus_2; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_2_io_i_mux_bus_3; // @[FlexDPU.scala 110:47]
  wire  flexdpecom4_3_clock; // @[FlexDPU.scala 110:47]
  wire  flexdpecom4_3_reset; // @[FlexDPU.scala 110:47]
  wire  flexdpecom4_3_io_i_data_valid; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_3_io_i_data_bus_0; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_3_io_i_data_bus_1; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_3_io_i_data_bus_2; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_3_io_i_data_bus_3; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_3_io_i_data_bus2_0; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_3_io_i_data_bus2_1; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_3_io_i_data_bus2_2; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_3_io_i_data_bus2_3; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_3_io_o_adder_0; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_3_io_o_adder_1; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_3_io_o_adder_2; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_3_io_i_mux_bus_0; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_3_io_i_mux_bus_1; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_3_io_i_mux_bus_2; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_3_io_i_mux_bus_3; // @[FlexDPU.scala 110:47]
  wire  flexdpecom4_4_clock; // @[FlexDPU.scala 110:47]
  wire  flexdpecom4_4_reset; // @[FlexDPU.scala 110:47]
  wire  flexdpecom4_4_io_i_data_valid; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_4_io_i_data_bus_0; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_4_io_i_data_bus_1; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_4_io_i_data_bus_2; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_4_io_i_data_bus_3; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_4_io_i_data_bus2_0; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_4_io_i_data_bus2_1; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_4_io_i_data_bus2_2; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_4_io_i_data_bus2_3; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_4_io_o_adder_0; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_4_io_o_adder_1; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_4_io_o_adder_2; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_4_io_i_mux_bus_0; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_4_io_i_mux_bus_1; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_4_io_i_mux_bus_2; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_4_io_i_mux_bus_3; // @[FlexDPU.scala 110:47]
  wire  flexdpecom4_5_clock; // @[FlexDPU.scala 110:47]
  wire  flexdpecom4_5_reset; // @[FlexDPU.scala 110:47]
  wire  flexdpecom4_5_io_i_data_valid; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_5_io_i_data_bus_0; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_5_io_i_data_bus_1; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_5_io_i_data_bus_2; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_5_io_i_data_bus_3; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_5_io_i_data_bus2_0; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_5_io_i_data_bus2_1; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_5_io_i_data_bus2_2; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_5_io_i_data_bus2_3; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_5_io_o_adder_0; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_5_io_o_adder_1; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_5_io_o_adder_2; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_5_io_i_mux_bus_0; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_5_io_i_mux_bus_1; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_5_io_i_mux_bus_2; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_5_io_i_mux_bus_3; // @[FlexDPU.scala 110:47]
  wire  flexdpecom4_6_clock; // @[FlexDPU.scala 110:47]
  wire  flexdpecom4_6_reset; // @[FlexDPU.scala 110:47]
  wire  flexdpecom4_6_io_i_data_valid; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_6_io_i_data_bus_0; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_6_io_i_data_bus_1; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_6_io_i_data_bus_2; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_6_io_i_data_bus_3; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_6_io_i_data_bus2_0; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_6_io_i_data_bus2_1; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_6_io_i_data_bus2_2; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_6_io_i_data_bus2_3; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_6_io_o_adder_0; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_6_io_o_adder_1; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_6_io_o_adder_2; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_6_io_i_mux_bus_0; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_6_io_i_mux_bus_1; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_6_io_i_mux_bus_2; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_6_io_i_mux_bus_3; // @[FlexDPU.scala 110:47]
  wire  flexdpecom4_7_clock; // @[FlexDPU.scala 110:47]
  wire  flexdpecom4_7_reset; // @[FlexDPU.scala 110:47]
  wire  flexdpecom4_7_io_i_data_valid; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_7_io_i_data_bus_0; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_7_io_i_data_bus_1; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_7_io_i_data_bus_2; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_7_io_i_data_bus_3; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_7_io_i_data_bus2_0; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_7_io_i_data_bus2_1; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_7_io_i_data_bus2_2; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_7_io_i_data_bus2_3; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_7_io_o_adder_0; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_7_io_o_adder_1; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_7_io_o_adder_2; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_7_io_i_mux_bus_0; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_7_io_i_mux_bus_1; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_7_io_i_mux_bus_2; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_7_io_i_mux_bus_3; // @[FlexDPU.scala 110:47]
  wire  flexdpecom4_8_clock; // @[FlexDPU.scala 110:47]
  wire  flexdpecom4_8_reset; // @[FlexDPU.scala 110:47]
  wire  flexdpecom4_8_io_i_data_valid; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_8_io_i_data_bus_0; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_8_io_i_data_bus_1; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_8_io_i_data_bus_2; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_8_io_i_data_bus_3; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_8_io_i_data_bus2_0; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_8_io_i_data_bus2_1; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_8_io_i_data_bus2_2; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_8_io_i_data_bus2_3; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_8_io_o_adder_0; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_8_io_o_adder_1; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_8_io_o_adder_2; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_8_io_i_mux_bus_0; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_8_io_i_mux_bus_1; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_8_io_i_mux_bus_2; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_8_io_i_mux_bus_3; // @[FlexDPU.scala 110:47]
  wire  flexdpecom4_9_clock; // @[FlexDPU.scala 110:47]
  wire  flexdpecom4_9_reset; // @[FlexDPU.scala 110:47]
  wire  flexdpecom4_9_io_i_data_valid; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_9_io_i_data_bus_0; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_9_io_i_data_bus_1; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_9_io_i_data_bus_2; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_9_io_i_data_bus_3; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_9_io_i_data_bus2_0; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_9_io_i_data_bus2_1; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_9_io_i_data_bus2_2; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_9_io_i_data_bus2_3; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_9_io_o_adder_0; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_9_io_o_adder_1; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_9_io_o_adder_2; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_9_io_i_mux_bus_0; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_9_io_i_mux_bus_1; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_9_io_i_mux_bus_2; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_9_io_i_mux_bus_3; // @[FlexDPU.scala 110:47]
  wire  flexdpecom4_10_clock; // @[FlexDPU.scala 110:47]
  wire  flexdpecom4_10_reset; // @[FlexDPU.scala 110:47]
  wire  flexdpecom4_10_io_i_data_valid; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_10_io_i_data_bus_0; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_10_io_i_data_bus_1; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_10_io_i_data_bus_2; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_10_io_i_data_bus_3; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_10_io_i_data_bus2_0; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_10_io_i_data_bus2_1; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_10_io_i_data_bus2_2; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_10_io_i_data_bus2_3; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_10_io_o_adder_0; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_10_io_o_adder_1; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_10_io_o_adder_2; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_10_io_i_mux_bus_0; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_10_io_i_mux_bus_1; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_10_io_i_mux_bus_2; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_10_io_i_mux_bus_3; // @[FlexDPU.scala 110:47]
  wire  flexdpecom4_11_clock; // @[FlexDPU.scala 110:47]
  wire  flexdpecom4_11_reset; // @[FlexDPU.scala 110:47]
  wire  flexdpecom4_11_io_i_data_valid; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_11_io_i_data_bus_0; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_11_io_i_data_bus_1; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_11_io_i_data_bus_2; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_11_io_i_data_bus_3; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_11_io_i_data_bus2_0; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_11_io_i_data_bus2_1; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_11_io_i_data_bus2_2; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_11_io_i_data_bus2_3; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_11_io_o_adder_0; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_11_io_o_adder_1; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_11_io_o_adder_2; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_11_io_i_mux_bus_0; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_11_io_i_mux_bus_1; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_11_io_i_mux_bus_2; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_11_io_i_mux_bus_3; // @[FlexDPU.scala 110:47]
  wire  flexdpecom4_12_clock; // @[FlexDPU.scala 110:47]
  wire  flexdpecom4_12_reset; // @[FlexDPU.scala 110:47]
  wire  flexdpecom4_12_io_i_data_valid; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_12_io_i_data_bus_0; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_12_io_i_data_bus_1; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_12_io_i_data_bus_2; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_12_io_i_data_bus_3; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_12_io_i_data_bus2_0; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_12_io_i_data_bus2_1; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_12_io_i_data_bus2_2; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_12_io_i_data_bus2_3; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_12_io_o_adder_0; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_12_io_o_adder_1; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_12_io_o_adder_2; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_12_io_i_mux_bus_0; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_12_io_i_mux_bus_1; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_12_io_i_mux_bus_2; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_12_io_i_mux_bus_3; // @[FlexDPU.scala 110:47]
  wire  flexdpecom4_13_clock; // @[FlexDPU.scala 110:47]
  wire  flexdpecom4_13_reset; // @[FlexDPU.scala 110:47]
  wire  flexdpecom4_13_io_i_data_valid; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_13_io_i_data_bus_0; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_13_io_i_data_bus_1; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_13_io_i_data_bus_2; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_13_io_i_data_bus_3; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_13_io_i_data_bus2_0; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_13_io_i_data_bus2_1; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_13_io_i_data_bus2_2; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_13_io_i_data_bus2_3; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_13_io_o_adder_0; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_13_io_o_adder_1; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_13_io_o_adder_2; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_13_io_i_mux_bus_0; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_13_io_i_mux_bus_1; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_13_io_i_mux_bus_2; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_13_io_i_mux_bus_3; // @[FlexDPU.scala 110:47]
  wire  flexdpecom4_14_clock; // @[FlexDPU.scala 110:47]
  wire  flexdpecom4_14_reset; // @[FlexDPU.scala 110:47]
  wire  flexdpecom4_14_io_i_data_valid; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_14_io_i_data_bus_0; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_14_io_i_data_bus_1; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_14_io_i_data_bus_2; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_14_io_i_data_bus_3; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_14_io_i_data_bus2_0; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_14_io_i_data_bus2_1; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_14_io_i_data_bus2_2; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_14_io_i_data_bus2_3; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_14_io_o_adder_0; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_14_io_o_adder_1; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_14_io_o_adder_2; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_14_io_i_mux_bus_0; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_14_io_i_mux_bus_1; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_14_io_i_mux_bus_2; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_14_io_i_mux_bus_3; // @[FlexDPU.scala 110:47]
  wire  flexdpecom4_15_clock; // @[FlexDPU.scala 110:47]
  wire  flexdpecom4_15_reset; // @[FlexDPU.scala 110:47]
  wire  flexdpecom4_15_io_i_data_valid; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_15_io_i_data_bus_0; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_15_io_i_data_bus_1; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_15_io_i_data_bus_2; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_15_io_i_data_bus_3; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_15_io_i_data_bus2_0; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_15_io_i_data_bus2_1; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_15_io_i_data_bus2_2; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_15_io_i_data_bus2_3; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_15_io_o_adder_0; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_15_io_o_adder_1; // @[FlexDPU.scala 110:47]
  wire [15:0] flexdpecom4_15_io_o_adder_2; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_15_io_i_mux_bus_0; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_15_io_i_mux_bus_1; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_15_io_i_mux_bus_2; // @[FlexDPU.scala 110:47]
  wire [3:0] flexdpecom4_15_io_i_mux_bus_3; // @[FlexDPU.scala 110:47]
  reg [31:0] used_FlexDPE_0; // @[FlexDPU.scala 19:27]
  reg [31:0] used_FlexDPE_1; // @[FlexDPU.scala 19:27]
  wire [31:0] equalDistribution = io_CalFDE / 2'h2; // @[FlexDPU.scala 21:39]
  wire [31:0] _GEN_0 = io_CalFDE % 32'h2; // @[FlexDPU.scala 22:43]
  wire [1:0] remainingDistribution = _GEN_0[1:0]; // @[FlexDPU.scala 22:43]
  wire [31:0] _used_FlexDPE_0_T_2 = equalDistribution + 32'h1; // @[FlexDPU.scala 25:73]
  reg [31:0] iloop; // @[FlexDPU.scala 33:24]
  reg [31:0] jloop; // @[FlexDPU.scala 34:24]
  reg  Statvalid; // @[FlexDPU.scala 35:28]
  wire  _Statvalid_T_1 = jloop == 32'h7; // @[FlexDPU.scala 37:61]
  wire  _Statvalid_T_2 = iloop == 32'h7 & jloop == 32'h7; // @[FlexDPU.scala 37:51]
  wire [31:0] _iloop_T_1 = iloop + 32'h1; // @[FlexDPU.scala 44:24]
  wire [31:0] _jloop_T_1 = jloop + 32'h1; // @[FlexDPU.scala 48:24]
  reg [31:0] PF1_Stream_Col_0; // @[FlexDPU.scala 61:33]
  reg [31:0] PF1_Stream_Col_1; // @[FlexDPU.scala 61:33]
  reg [31:0] PF1_Stream_Col_2; // @[FlexDPU.scala 61:33]
  reg [31:0] PF1_Stream_Col_3; // @[FlexDPU.scala 61:33]
  reg [31:0] PF1_Stream_Col_4; // @[FlexDPU.scala 61:33]
  reg [31:0] PF1_Stream_Col_5; // @[FlexDPU.scala 61:33]
  reg [31:0] PF1_Stream_Col_6; // @[FlexDPU.scala 61:33]
  reg [31:0] PF1_Stream_Col_7; // @[FlexDPU.scala 61:33]
  reg [31:0] ModuleIndex; // @[FlexDPU.scala 62:30]
  wire [31:0] _ModuleIndex_T_1 = ModuleIndex + 32'h1; // @[FlexDPU.scala 154:40]
  wire  PF_0_PF_Valid = PathFinder_io_PF_Valid; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] _GEN_263 = 3'h1 == ModuleIndex[2:0] ? io_Streaming_matrix_0_1 : io_Streaming_matrix_0_0; // @[FlexDPU.scala 164:{31,31}]
  wire [15:0] _GEN_264 = 3'h2 == ModuleIndex[2:0] ? io_Streaming_matrix_0_2 : _GEN_263; // @[FlexDPU.scala 164:{31,31}]
  wire [15:0] _GEN_265 = 3'h3 == ModuleIndex[2:0] ? io_Streaming_matrix_0_3 : _GEN_264; // @[FlexDPU.scala 164:{31,31}]
  wire [15:0] _GEN_266 = 3'h4 == ModuleIndex[2:0] ? io_Streaming_matrix_0_4 : _GEN_265; // @[FlexDPU.scala 164:{31,31}]
  wire [15:0] _GEN_267 = 3'h5 == ModuleIndex[2:0] ? io_Streaming_matrix_0_5 : _GEN_266; // @[FlexDPU.scala 164:{31,31}]
  wire [15:0] _GEN_268 = 3'h6 == ModuleIndex[2:0] ? io_Streaming_matrix_0_6 : _GEN_267; // @[FlexDPU.scala 164:{31,31}]
  wire [15:0] _GEN_269 = 3'h7 == ModuleIndex[2:0] ? io_Streaming_matrix_0_7 : _GEN_268; // @[FlexDPU.scala 164:{31,31}]
  wire [15:0] _GEN_271 = 3'h1 == ModuleIndex[2:0] ? io_Streaming_matrix_1_1 : io_Streaming_matrix_1_0; // @[FlexDPU.scala 164:{31,31}]
  wire [15:0] _GEN_272 = 3'h2 == ModuleIndex[2:0] ? io_Streaming_matrix_1_2 : _GEN_271; // @[FlexDPU.scala 164:{31,31}]
  wire [15:0] _GEN_273 = 3'h3 == ModuleIndex[2:0] ? io_Streaming_matrix_1_3 : _GEN_272; // @[FlexDPU.scala 164:{31,31}]
  wire [15:0] _GEN_274 = 3'h4 == ModuleIndex[2:0] ? io_Streaming_matrix_1_4 : _GEN_273; // @[FlexDPU.scala 164:{31,31}]
  wire [15:0] _GEN_275 = 3'h5 == ModuleIndex[2:0] ? io_Streaming_matrix_1_5 : _GEN_274; // @[FlexDPU.scala 164:{31,31}]
  wire [15:0] _GEN_276 = 3'h6 == ModuleIndex[2:0] ? io_Streaming_matrix_1_6 : _GEN_275; // @[FlexDPU.scala 164:{31,31}]
  wire [15:0] _GEN_277 = 3'h7 == ModuleIndex[2:0] ? io_Streaming_matrix_1_7 : _GEN_276; // @[FlexDPU.scala 164:{31,31}]
  wire [15:0] _GEN_279 = 3'h1 == ModuleIndex[2:0] ? io_Streaming_matrix_2_1 : io_Streaming_matrix_2_0; // @[FlexDPU.scala 164:{31,31}]
  wire [15:0] _GEN_280 = 3'h2 == ModuleIndex[2:0] ? io_Streaming_matrix_2_2 : _GEN_279; // @[FlexDPU.scala 164:{31,31}]
  wire [15:0] _GEN_281 = 3'h3 == ModuleIndex[2:0] ? io_Streaming_matrix_2_3 : _GEN_280; // @[FlexDPU.scala 164:{31,31}]
  wire [15:0] _GEN_282 = 3'h4 == ModuleIndex[2:0] ? io_Streaming_matrix_2_4 : _GEN_281; // @[FlexDPU.scala 164:{31,31}]
  wire [15:0] _GEN_283 = 3'h5 == ModuleIndex[2:0] ? io_Streaming_matrix_2_5 : _GEN_282; // @[FlexDPU.scala 164:{31,31}]
  wire [15:0] _GEN_284 = 3'h6 == ModuleIndex[2:0] ? io_Streaming_matrix_2_6 : _GEN_283; // @[FlexDPU.scala 164:{31,31}]
  wire [15:0] _GEN_285 = 3'h7 == ModuleIndex[2:0] ? io_Streaming_matrix_2_7 : _GEN_284; // @[FlexDPU.scala 164:{31,31}]
  wire [15:0] _GEN_287 = 3'h1 == ModuleIndex[2:0] ? io_Streaming_matrix_3_1 : io_Streaming_matrix_3_0; // @[FlexDPU.scala 164:{31,31}]
  wire [15:0] _GEN_288 = 3'h2 == ModuleIndex[2:0] ? io_Streaming_matrix_3_2 : _GEN_287; // @[FlexDPU.scala 164:{31,31}]
  wire [15:0] _GEN_289 = 3'h3 == ModuleIndex[2:0] ? io_Streaming_matrix_3_3 : _GEN_288; // @[FlexDPU.scala 164:{31,31}]
  wire [15:0] _GEN_290 = 3'h4 == ModuleIndex[2:0] ? io_Streaming_matrix_3_4 : _GEN_289; // @[FlexDPU.scala 164:{31,31}]
  wire [15:0] _GEN_291 = 3'h5 == ModuleIndex[2:0] ? io_Streaming_matrix_3_5 : _GEN_290; // @[FlexDPU.scala 164:{31,31}]
  wire [15:0] _GEN_292 = 3'h6 == ModuleIndex[2:0] ? io_Streaming_matrix_3_6 : _GEN_291; // @[FlexDPU.scala 164:{31,31}]
  wire [15:0] _GEN_293 = 3'h7 == ModuleIndex[2:0] ? io_Streaming_matrix_3_7 : _GEN_292; // @[FlexDPU.scala 164:{31,31}]
  wire [15:0] _GEN_295 = 3'h1 == ModuleIndex[2:0] ? io_Streaming_matrix_4_1 : io_Streaming_matrix_4_0; // @[FlexDPU.scala 164:{31,31}]
  wire [15:0] _GEN_296 = 3'h2 == ModuleIndex[2:0] ? io_Streaming_matrix_4_2 : _GEN_295; // @[FlexDPU.scala 164:{31,31}]
  wire [15:0] _GEN_297 = 3'h3 == ModuleIndex[2:0] ? io_Streaming_matrix_4_3 : _GEN_296; // @[FlexDPU.scala 164:{31,31}]
  wire [15:0] _GEN_298 = 3'h4 == ModuleIndex[2:0] ? io_Streaming_matrix_4_4 : _GEN_297; // @[FlexDPU.scala 164:{31,31}]
  wire [15:0] _GEN_299 = 3'h5 == ModuleIndex[2:0] ? io_Streaming_matrix_4_5 : _GEN_298; // @[FlexDPU.scala 164:{31,31}]
  wire [15:0] _GEN_300 = 3'h6 == ModuleIndex[2:0] ? io_Streaming_matrix_4_6 : _GEN_299; // @[FlexDPU.scala 164:{31,31}]
  wire [15:0] _GEN_301 = 3'h7 == ModuleIndex[2:0] ? io_Streaming_matrix_4_7 : _GEN_300; // @[FlexDPU.scala 164:{31,31}]
  wire [15:0] _GEN_303 = 3'h1 == ModuleIndex[2:0] ? io_Streaming_matrix_5_1 : io_Streaming_matrix_5_0; // @[FlexDPU.scala 164:{31,31}]
  wire [15:0] _GEN_304 = 3'h2 == ModuleIndex[2:0] ? io_Streaming_matrix_5_2 : _GEN_303; // @[FlexDPU.scala 164:{31,31}]
  wire [15:0] _GEN_305 = 3'h3 == ModuleIndex[2:0] ? io_Streaming_matrix_5_3 : _GEN_304; // @[FlexDPU.scala 164:{31,31}]
  wire [15:0] _GEN_306 = 3'h4 == ModuleIndex[2:0] ? io_Streaming_matrix_5_4 : _GEN_305; // @[FlexDPU.scala 164:{31,31}]
  wire [15:0] _GEN_307 = 3'h5 == ModuleIndex[2:0] ? io_Streaming_matrix_5_5 : _GEN_306; // @[FlexDPU.scala 164:{31,31}]
  wire [15:0] _GEN_308 = 3'h6 == ModuleIndex[2:0] ? io_Streaming_matrix_5_6 : _GEN_307; // @[FlexDPU.scala 164:{31,31}]
  wire [15:0] _GEN_309 = 3'h7 == ModuleIndex[2:0] ? io_Streaming_matrix_5_7 : _GEN_308; // @[FlexDPU.scala 164:{31,31}]
  wire [15:0] _GEN_311 = 3'h1 == ModuleIndex[2:0] ? io_Streaming_matrix_6_1 : io_Streaming_matrix_6_0; // @[FlexDPU.scala 164:{31,31}]
  wire [15:0] _GEN_312 = 3'h2 == ModuleIndex[2:0] ? io_Streaming_matrix_6_2 : _GEN_311; // @[FlexDPU.scala 164:{31,31}]
  wire [15:0] _GEN_313 = 3'h3 == ModuleIndex[2:0] ? io_Streaming_matrix_6_3 : _GEN_312; // @[FlexDPU.scala 164:{31,31}]
  wire [15:0] _GEN_314 = 3'h4 == ModuleIndex[2:0] ? io_Streaming_matrix_6_4 : _GEN_313; // @[FlexDPU.scala 164:{31,31}]
  wire [15:0] _GEN_315 = 3'h5 == ModuleIndex[2:0] ? io_Streaming_matrix_6_5 : _GEN_314; // @[FlexDPU.scala 164:{31,31}]
  wire [15:0] _GEN_316 = 3'h6 == ModuleIndex[2:0] ? io_Streaming_matrix_6_6 : _GEN_315; // @[FlexDPU.scala 164:{31,31}]
  wire [15:0] _GEN_317 = 3'h7 == ModuleIndex[2:0] ? io_Streaming_matrix_6_7 : _GEN_316; // @[FlexDPU.scala 164:{31,31}]
  wire [15:0] _GEN_319 = 3'h1 == ModuleIndex[2:0] ? io_Streaming_matrix_7_1 : io_Streaming_matrix_7_0; // @[FlexDPU.scala 164:{31,31}]
  wire [15:0] _GEN_320 = 3'h2 == ModuleIndex[2:0] ? io_Streaming_matrix_7_2 : _GEN_319; // @[FlexDPU.scala 164:{31,31}]
  wire [15:0] _GEN_321 = 3'h3 == ModuleIndex[2:0] ? io_Streaming_matrix_7_3 : _GEN_320; // @[FlexDPU.scala 164:{31,31}]
  wire [15:0] _GEN_322 = 3'h4 == ModuleIndex[2:0] ? io_Streaming_matrix_7_4 : _GEN_321; // @[FlexDPU.scala 164:{31,31}]
  wire [15:0] _GEN_323 = 3'h5 == ModuleIndex[2:0] ? io_Streaming_matrix_7_5 : _GEN_322; // @[FlexDPU.scala 164:{31,31}]
  wire [15:0] _GEN_324 = 3'h6 == ModuleIndex[2:0] ? io_Streaming_matrix_7_6 : _GEN_323; // @[FlexDPU.scala 164:{31,31}]
  wire [15:0] _GEN_325 = 3'h7 == ModuleIndex[2:0] ? io_Streaming_matrix_7_7 : _GEN_324; // @[FlexDPU.scala 164:{31,31}]
  wire [31:0] _GEN_392 = Statvalid ? PF1_Stream_Col_0 : 32'h0; // @[FlexDPU.scala 98:20 104:32 84:32]
  wire [31:0] _GEN_393 = Statvalid ? PF1_Stream_Col_1 : 32'h0; // @[FlexDPU.scala 98:20 104:32 84:32]
  wire [31:0] _GEN_394 = Statvalid ? PF1_Stream_Col_2 : 32'h0; // @[FlexDPU.scala 98:20 104:32 84:32]
  wire [31:0] _GEN_395 = Statvalid ? PF1_Stream_Col_3 : 32'h0; // @[FlexDPU.scala 98:20 104:32 84:32]
  wire [31:0] _GEN_396 = Statvalid ? PF1_Stream_Col_4 : 32'h0; // @[FlexDPU.scala 98:20 104:32 84:32]
  wire [31:0] _GEN_397 = Statvalid ? PF1_Stream_Col_5 : 32'h0; // @[FlexDPU.scala 98:20 104:32 84:32]
  wire [31:0] _GEN_398 = Statvalid ? PF1_Stream_Col_6 : 32'h0; // @[FlexDPU.scala 98:20 104:32 84:32]
  wire [31:0] _GEN_399 = Statvalid ? PF1_Stream_Col_7 : 32'h0; // @[FlexDPU.scala 98:20 104:32 84:32]
  wire [1:0] _GEN_729 = Statvalid ? 2'h2 : 2'h0; // @[FlexDPU.scala 98:20 103:21 83:21]
  wire [1:0] _GEN_802 = Statvalid ? 2'h3 : 2'h0; // @[FlexDPU.scala 98:20 103:21 83:21]
  wire [2:0] _GEN_875 = Statvalid ? 3'h4 : 3'h0; // @[FlexDPU.scala 98:20 103:21 83:21]
  wire [2:0] _GEN_948 = Statvalid ? 3'h5 : 3'h0; // @[FlexDPU.scala 98:20 103:21 83:21]
  wire [2:0] _GEN_1021 = Statvalid ? 3'h6 : 3'h0; // @[FlexDPU.scala 98:20 103:21 83:21]
  wire [2:0] _GEN_1094 = Statvalid ? 3'h7 : 3'h0; // @[FlexDPU.scala 98:20 103:21 83:21]
  wire [3:0] _GEN_1167 = Statvalid ? 4'h8 : 4'h0; // @[FlexDPU.scala 98:20 103:21 83:21]
  wire [3:0] _GEN_1240 = Statvalid ? 4'h9 : 4'h0; // @[FlexDPU.scala 98:20 103:21 83:21]
  wire [3:0] _GEN_1313 = Statvalid ? 4'ha : 4'h0; // @[FlexDPU.scala 98:20 103:21 83:21]
  wire [3:0] _GEN_1386 = Statvalid ? 4'hb : 4'h0; // @[FlexDPU.scala 98:20 103:21 83:21]
  wire [3:0] _GEN_1459 = Statvalid ? 4'hc : 4'h0; // @[FlexDPU.scala 98:20 103:21 83:21]
  wire [3:0] _GEN_1532 = Statvalid ? 4'hd : 4'h0; // @[FlexDPU.scala 98:20 103:21 83:21]
  wire [3:0] _GEN_1605 = Statvalid ? 4'he : 4'h0; // @[FlexDPU.scala 98:20 103:21 83:21]
  wire [3:0] _GEN_1678 = Statvalid ? 4'hf : 4'h0; // @[FlexDPU.scala 98:20 103:21 83:21]
  wire [15:0] FDPE_0_o_adder_0 = flexdpecom4_io_o_adder_0; // @[FlexDPU.scala 110:{27,27}]
  wire [15:0] FDPE_0_o_adder_1 = flexdpecom4_io_o_adder_1; // @[FlexDPU.scala 110:{27,27}]
  wire [15:0] FDPE_0_o_adder_2 = flexdpecom4_io_o_adder_2; // @[FlexDPU.scala 110:{27,27}]
  wire [15:0] FDPE_1_o_adder_0 = flexdpecom4_1_io_o_adder_0; // @[FlexDPU.scala 110:{27,27}]
  wire [15:0] FDPE_1_o_adder_1 = flexdpecom4_1_io_o_adder_1; // @[FlexDPU.scala 110:{27,27}]
  wire [15:0] FDPE_1_o_adder_2 = flexdpecom4_1_io_o_adder_2; // @[FlexDPU.scala 110:{27,27}]
  wire [15:0] FDPE_2_o_adder_0 = flexdpecom4_2_io_o_adder_0; // @[FlexDPU.scala 110:{27,27}]
  wire [15:0] FDPE_2_o_adder_1 = flexdpecom4_2_io_o_adder_1; // @[FlexDPU.scala 110:{27,27}]
  wire [15:0] FDPE_2_o_adder_2 = flexdpecom4_2_io_o_adder_2; // @[FlexDPU.scala 110:{27,27}]
  wire [15:0] FDPE_3_o_adder_0 = flexdpecom4_3_io_o_adder_0; // @[FlexDPU.scala 110:{27,27}]
  wire [15:0] FDPE_3_o_adder_1 = flexdpecom4_3_io_o_adder_1; // @[FlexDPU.scala 110:{27,27}]
  wire [15:0] FDPE_3_o_adder_2 = flexdpecom4_3_io_o_adder_2; // @[FlexDPU.scala 110:{27,27}]
  wire [15:0] FDPE_4_o_adder_0 = flexdpecom4_4_io_o_adder_0; // @[FlexDPU.scala 110:{27,27}]
  wire [15:0] FDPE_4_o_adder_1 = flexdpecom4_4_io_o_adder_1; // @[FlexDPU.scala 110:{27,27}]
  wire [15:0] FDPE_4_o_adder_2 = flexdpecom4_4_io_o_adder_2; // @[FlexDPU.scala 110:{27,27}]
  wire [15:0] FDPE_5_o_adder_0 = flexdpecom4_5_io_o_adder_0; // @[FlexDPU.scala 110:{27,27}]
  wire [15:0] FDPE_5_o_adder_1 = flexdpecom4_5_io_o_adder_1; // @[FlexDPU.scala 110:{27,27}]
  wire [15:0] FDPE_5_o_adder_2 = flexdpecom4_5_io_o_adder_2; // @[FlexDPU.scala 110:{27,27}]
  wire [15:0] FDPE_6_o_adder_0 = flexdpecom4_6_io_o_adder_0; // @[FlexDPU.scala 110:{27,27}]
  wire [15:0] FDPE_6_o_adder_1 = flexdpecom4_6_io_o_adder_1; // @[FlexDPU.scala 110:{27,27}]
  wire [15:0] FDPE_6_o_adder_2 = flexdpecom4_6_io_o_adder_2; // @[FlexDPU.scala 110:{27,27}]
  wire [15:0] FDPE_7_o_adder_0 = flexdpecom4_7_io_o_adder_0; // @[FlexDPU.scala 110:{27,27}]
  wire [15:0] FDPE_7_o_adder_1 = flexdpecom4_7_io_o_adder_1; // @[FlexDPU.scala 110:{27,27}]
  wire [15:0] FDPE_7_o_adder_2 = flexdpecom4_7_io_o_adder_2; // @[FlexDPU.scala 110:{27,27}]
  wire [15:0] FDPE_8_o_adder_0 = flexdpecom4_8_io_o_adder_0; // @[FlexDPU.scala 110:{27,27}]
  wire [15:0] FDPE_8_o_adder_1 = flexdpecom4_8_io_o_adder_1; // @[FlexDPU.scala 110:{27,27}]
  wire [15:0] FDPE_8_o_adder_2 = flexdpecom4_8_io_o_adder_2; // @[FlexDPU.scala 110:{27,27}]
  wire [15:0] FDPE_9_o_adder_0 = flexdpecom4_9_io_o_adder_0; // @[FlexDPU.scala 110:{27,27}]
  wire [15:0] FDPE_9_o_adder_1 = flexdpecom4_9_io_o_adder_1; // @[FlexDPU.scala 110:{27,27}]
  wire [15:0] FDPE_9_o_adder_2 = flexdpecom4_9_io_o_adder_2; // @[FlexDPU.scala 110:{27,27}]
  wire [15:0] FDPE_10_o_adder_0 = flexdpecom4_10_io_o_adder_0; // @[FlexDPU.scala 110:{27,27}]
  wire [15:0] FDPE_10_o_adder_1 = flexdpecom4_10_io_o_adder_1; // @[FlexDPU.scala 110:{27,27}]
  wire [15:0] FDPE_10_o_adder_2 = flexdpecom4_10_io_o_adder_2; // @[FlexDPU.scala 110:{27,27}]
  wire [15:0] FDPE_11_o_adder_0 = flexdpecom4_11_io_o_adder_0; // @[FlexDPU.scala 110:{27,27}]
  wire [15:0] FDPE_11_o_adder_1 = flexdpecom4_11_io_o_adder_1; // @[FlexDPU.scala 110:{27,27}]
  wire [15:0] FDPE_11_o_adder_2 = flexdpecom4_11_io_o_adder_2; // @[FlexDPU.scala 110:{27,27}]
  wire [15:0] FDPE_12_o_adder_0 = flexdpecom4_12_io_o_adder_0; // @[FlexDPU.scala 110:{27,27}]
  wire [15:0] FDPE_12_o_adder_1 = flexdpecom4_12_io_o_adder_1; // @[FlexDPU.scala 110:{27,27}]
  wire [15:0] FDPE_12_o_adder_2 = flexdpecom4_12_io_o_adder_2; // @[FlexDPU.scala 110:{27,27}]
  wire [15:0] FDPE_13_o_adder_0 = flexdpecom4_13_io_o_adder_0; // @[FlexDPU.scala 110:{27,27}]
  wire [15:0] FDPE_13_o_adder_1 = flexdpecom4_13_io_o_adder_1; // @[FlexDPU.scala 110:{27,27}]
  wire [15:0] FDPE_13_o_adder_2 = flexdpecom4_13_io_o_adder_2; // @[FlexDPU.scala 110:{27,27}]
  wire [15:0] FDPE_14_o_adder_0 = flexdpecom4_14_io_o_adder_0; // @[FlexDPU.scala 110:{27,27}]
  wire [15:0] FDPE_14_o_adder_1 = flexdpecom4_14_io_o_adder_1; // @[FlexDPU.scala 110:{27,27}]
  wire [15:0] FDPE_14_o_adder_2 = flexdpecom4_14_io_o_adder_2; // @[FlexDPU.scala 110:{27,27}]
  wire [15:0] FDPE_15_o_adder_0 = flexdpecom4_15_io_o_adder_0; // @[FlexDPU.scala 110:{27,27}]
  wire [15:0] FDPE_15_o_adder_1 = flexdpecom4_15_io_o_adder_1; // @[FlexDPU.scala 110:{27,27}]
  wire [15:0] FDPE_15_o_adder_2 = flexdpecom4_15_io_o_adder_2; // @[FlexDPU.scala 110:{27,27}]
  PathFinder PathFinder ( // @[FlexDPU.scala 77:41]
    .clock(PathFinder_clock),
    .reset(PathFinder_reset),
    .io_Stationary_matrix_0_0(PathFinder_io_Stationary_matrix_0_0),
    .io_Stationary_matrix_0_1(PathFinder_io_Stationary_matrix_0_1),
    .io_Stationary_matrix_0_2(PathFinder_io_Stationary_matrix_0_2),
    .io_Stationary_matrix_0_3(PathFinder_io_Stationary_matrix_0_3),
    .io_Stationary_matrix_0_4(PathFinder_io_Stationary_matrix_0_4),
    .io_Stationary_matrix_0_5(PathFinder_io_Stationary_matrix_0_5),
    .io_Stationary_matrix_0_6(PathFinder_io_Stationary_matrix_0_6),
    .io_Stationary_matrix_0_7(PathFinder_io_Stationary_matrix_0_7),
    .io_Stationary_matrix_1_0(PathFinder_io_Stationary_matrix_1_0),
    .io_Stationary_matrix_1_1(PathFinder_io_Stationary_matrix_1_1),
    .io_Stationary_matrix_1_2(PathFinder_io_Stationary_matrix_1_2),
    .io_Stationary_matrix_1_3(PathFinder_io_Stationary_matrix_1_3),
    .io_Stationary_matrix_1_4(PathFinder_io_Stationary_matrix_1_4),
    .io_Stationary_matrix_1_5(PathFinder_io_Stationary_matrix_1_5),
    .io_Stationary_matrix_1_6(PathFinder_io_Stationary_matrix_1_6),
    .io_Stationary_matrix_1_7(PathFinder_io_Stationary_matrix_1_7),
    .io_Stationary_matrix_2_0(PathFinder_io_Stationary_matrix_2_0),
    .io_Stationary_matrix_2_1(PathFinder_io_Stationary_matrix_2_1),
    .io_Stationary_matrix_2_2(PathFinder_io_Stationary_matrix_2_2),
    .io_Stationary_matrix_2_3(PathFinder_io_Stationary_matrix_2_3),
    .io_Stationary_matrix_2_4(PathFinder_io_Stationary_matrix_2_4),
    .io_Stationary_matrix_2_5(PathFinder_io_Stationary_matrix_2_5),
    .io_Stationary_matrix_2_6(PathFinder_io_Stationary_matrix_2_6),
    .io_Stationary_matrix_2_7(PathFinder_io_Stationary_matrix_2_7),
    .io_Stationary_matrix_3_0(PathFinder_io_Stationary_matrix_3_0),
    .io_Stationary_matrix_3_1(PathFinder_io_Stationary_matrix_3_1),
    .io_Stationary_matrix_3_2(PathFinder_io_Stationary_matrix_3_2),
    .io_Stationary_matrix_3_3(PathFinder_io_Stationary_matrix_3_3),
    .io_Stationary_matrix_3_4(PathFinder_io_Stationary_matrix_3_4),
    .io_Stationary_matrix_3_5(PathFinder_io_Stationary_matrix_3_5),
    .io_Stationary_matrix_3_6(PathFinder_io_Stationary_matrix_3_6),
    .io_Stationary_matrix_3_7(PathFinder_io_Stationary_matrix_3_7),
    .io_Stationary_matrix_4_0(PathFinder_io_Stationary_matrix_4_0),
    .io_Stationary_matrix_4_1(PathFinder_io_Stationary_matrix_4_1),
    .io_Stationary_matrix_4_2(PathFinder_io_Stationary_matrix_4_2),
    .io_Stationary_matrix_4_3(PathFinder_io_Stationary_matrix_4_3),
    .io_Stationary_matrix_4_4(PathFinder_io_Stationary_matrix_4_4),
    .io_Stationary_matrix_4_5(PathFinder_io_Stationary_matrix_4_5),
    .io_Stationary_matrix_4_6(PathFinder_io_Stationary_matrix_4_6),
    .io_Stationary_matrix_4_7(PathFinder_io_Stationary_matrix_4_7),
    .io_Stationary_matrix_5_0(PathFinder_io_Stationary_matrix_5_0),
    .io_Stationary_matrix_5_1(PathFinder_io_Stationary_matrix_5_1),
    .io_Stationary_matrix_5_2(PathFinder_io_Stationary_matrix_5_2),
    .io_Stationary_matrix_5_3(PathFinder_io_Stationary_matrix_5_3),
    .io_Stationary_matrix_5_4(PathFinder_io_Stationary_matrix_5_4),
    .io_Stationary_matrix_5_5(PathFinder_io_Stationary_matrix_5_5),
    .io_Stationary_matrix_5_6(PathFinder_io_Stationary_matrix_5_6),
    .io_Stationary_matrix_5_7(PathFinder_io_Stationary_matrix_5_7),
    .io_Stationary_matrix_6_0(PathFinder_io_Stationary_matrix_6_0),
    .io_Stationary_matrix_6_1(PathFinder_io_Stationary_matrix_6_1),
    .io_Stationary_matrix_6_2(PathFinder_io_Stationary_matrix_6_2),
    .io_Stationary_matrix_6_3(PathFinder_io_Stationary_matrix_6_3),
    .io_Stationary_matrix_6_4(PathFinder_io_Stationary_matrix_6_4),
    .io_Stationary_matrix_6_5(PathFinder_io_Stationary_matrix_6_5),
    .io_Stationary_matrix_6_6(PathFinder_io_Stationary_matrix_6_6),
    .io_Stationary_matrix_6_7(PathFinder_io_Stationary_matrix_6_7),
    .io_Stationary_matrix_7_0(PathFinder_io_Stationary_matrix_7_0),
    .io_Stationary_matrix_7_1(PathFinder_io_Stationary_matrix_7_1),
    .io_Stationary_matrix_7_2(PathFinder_io_Stationary_matrix_7_2),
    .io_Stationary_matrix_7_3(PathFinder_io_Stationary_matrix_7_3),
    .io_Stationary_matrix_7_4(PathFinder_io_Stationary_matrix_7_4),
    .io_Stationary_matrix_7_5(PathFinder_io_Stationary_matrix_7_5),
    .io_Stationary_matrix_7_6(PathFinder_io_Stationary_matrix_7_6),
    .io_Stationary_matrix_7_7(PathFinder_io_Stationary_matrix_7_7),
    .io_Streaming_matrix_0(PathFinder_io_Streaming_matrix_0),
    .io_Streaming_matrix_1(PathFinder_io_Streaming_matrix_1),
    .io_Streaming_matrix_2(PathFinder_io_Streaming_matrix_2),
    .io_Streaming_matrix_3(PathFinder_io_Streaming_matrix_3),
    .io_Streaming_matrix_4(PathFinder_io_Streaming_matrix_4),
    .io_Streaming_matrix_5(PathFinder_io_Streaming_matrix_5),
    .io_Streaming_matrix_6(PathFinder_io_Streaming_matrix_6),
    .io_Streaming_matrix_7(PathFinder_io_Streaming_matrix_7),
    .io_i_mux_bus_0(PathFinder_io_i_mux_bus_0),
    .io_i_mux_bus_1(PathFinder_io_i_mux_bus_1),
    .io_i_mux_bus_2(PathFinder_io_i_mux_bus_2),
    .io_i_mux_bus_3(PathFinder_io_i_mux_bus_3),
    .io_Source_0(PathFinder_io_Source_0),
    .io_Source_1(PathFinder_io_Source_1),
    .io_Source_2(PathFinder_io_Source_2),
    .io_Source_3(PathFinder_io_Source_3),
    .io_destination_0(PathFinder_io_destination_0),
    .io_destination_1(PathFinder_io_destination_1),
    .io_destination_2(PathFinder_io_destination_2),
    .io_destination_3(PathFinder_io_destination_3),
    .io_PF_Valid(PathFinder_io_PF_Valid),
    .io_NoDPE(PathFinder_io_NoDPE),
    .io_DataValid(PathFinder_io_DataValid)
  );
  PathFinder PathFinder_1 ( // @[FlexDPU.scala 77:41]
    .clock(PathFinder_1_clock),
    .reset(PathFinder_1_reset),
    .io_Stationary_matrix_0_0(PathFinder_1_io_Stationary_matrix_0_0),
    .io_Stationary_matrix_0_1(PathFinder_1_io_Stationary_matrix_0_1),
    .io_Stationary_matrix_0_2(PathFinder_1_io_Stationary_matrix_0_2),
    .io_Stationary_matrix_0_3(PathFinder_1_io_Stationary_matrix_0_3),
    .io_Stationary_matrix_0_4(PathFinder_1_io_Stationary_matrix_0_4),
    .io_Stationary_matrix_0_5(PathFinder_1_io_Stationary_matrix_0_5),
    .io_Stationary_matrix_0_6(PathFinder_1_io_Stationary_matrix_0_6),
    .io_Stationary_matrix_0_7(PathFinder_1_io_Stationary_matrix_0_7),
    .io_Stationary_matrix_1_0(PathFinder_1_io_Stationary_matrix_1_0),
    .io_Stationary_matrix_1_1(PathFinder_1_io_Stationary_matrix_1_1),
    .io_Stationary_matrix_1_2(PathFinder_1_io_Stationary_matrix_1_2),
    .io_Stationary_matrix_1_3(PathFinder_1_io_Stationary_matrix_1_3),
    .io_Stationary_matrix_1_4(PathFinder_1_io_Stationary_matrix_1_4),
    .io_Stationary_matrix_1_5(PathFinder_1_io_Stationary_matrix_1_5),
    .io_Stationary_matrix_1_6(PathFinder_1_io_Stationary_matrix_1_6),
    .io_Stationary_matrix_1_7(PathFinder_1_io_Stationary_matrix_1_7),
    .io_Stationary_matrix_2_0(PathFinder_1_io_Stationary_matrix_2_0),
    .io_Stationary_matrix_2_1(PathFinder_1_io_Stationary_matrix_2_1),
    .io_Stationary_matrix_2_2(PathFinder_1_io_Stationary_matrix_2_2),
    .io_Stationary_matrix_2_3(PathFinder_1_io_Stationary_matrix_2_3),
    .io_Stationary_matrix_2_4(PathFinder_1_io_Stationary_matrix_2_4),
    .io_Stationary_matrix_2_5(PathFinder_1_io_Stationary_matrix_2_5),
    .io_Stationary_matrix_2_6(PathFinder_1_io_Stationary_matrix_2_6),
    .io_Stationary_matrix_2_7(PathFinder_1_io_Stationary_matrix_2_7),
    .io_Stationary_matrix_3_0(PathFinder_1_io_Stationary_matrix_3_0),
    .io_Stationary_matrix_3_1(PathFinder_1_io_Stationary_matrix_3_1),
    .io_Stationary_matrix_3_2(PathFinder_1_io_Stationary_matrix_3_2),
    .io_Stationary_matrix_3_3(PathFinder_1_io_Stationary_matrix_3_3),
    .io_Stationary_matrix_3_4(PathFinder_1_io_Stationary_matrix_3_4),
    .io_Stationary_matrix_3_5(PathFinder_1_io_Stationary_matrix_3_5),
    .io_Stationary_matrix_3_6(PathFinder_1_io_Stationary_matrix_3_6),
    .io_Stationary_matrix_3_7(PathFinder_1_io_Stationary_matrix_3_7),
    .io_Stationary_matrix_4_0(PathFinder_1_io_Stationary_matrix_4_0),
    .io_Stationary_matrix_4_1(PathFinder_1_io_Stationary_matrix_4_1),
    .io_Stationary_matrix_4_2(PathFinder_1_io_Stationary_matrix_4_2),
    .io_Stationary_matrix_4_3(PathFinder_1_io_Stationary_matrix_4_3),
    .io_Stationary_matrix_4_4(PathFinder_1_io_Stationary_matrix_4_4),
    .io_Stationary_matrix_4_5(PathFinder_1_io_Stationary_matrix_4_5),
    .io_Stationary_matrix_4_6(PathFinder_1_io_Stationary_matrix_4_6),
    .io_Stationary_matrix_4_7(PathFinder_1_io_Stationary_matrix_4_7),
    .io_Stationary_matrix_5_0(PathFinder_1_io_Stationary_matrix_5_0),
    .io_Stationary_matrix_5_1(PathFinder_1_io_Stationary_matrix_5_1),
    .io_Stationary_matrix_5_2(PathFinder_1_io_Stationary_matrix_5_2),
    .io_Stationary_matrix_5_3(PathFinder_1_io_Stationary_matrix_5_3),
    .io_Stationary_matrix_5_4(PathFinder_1_io_Stationary_matrix_5_4),
    .io_Stationary_matrix_5_5(PathFinder_1_io_Stationary_matrix_5_5),
    .io_Stationary_matrix_5_6(PathFinder_1_io_Stationary_matrix_5_6),
    .io_Stationary_matrix_5_7(PathFinder_1_io_Stationary_matrix_5_7),
    .io_Stationary_matrix_6_0(PathFinder_1_io_Stationary_matrix_6_0),
    .io_Stationary_matrix_6_1(PathFinder_1_io_Stationary_matrix_6_1),
    .io_Stationary_matrix_6_2(PathFinder_1_io_Stationary_matrix_6_2),
    .io_Stationary_matrix_6_3(PathFinder_1_io_Stationary_matrix_6_3),
    .io_Stationary_matrix_6_4(PathFinder_1_io_Stationary_matrix_6_4),
    .io_Stationary_matrix_6_5(PathFinder_1_io_Stationary_matrix_6_5),
    .io_Stationary_matrix_6_6(PathFinder_1_io_Stationary_matrix_6_6),
    .io_Stationary_matrix_6_7(PathFinder_1_io_Stationary_matrix_6_7),
    .io_Stationary_matrix_7_0(PathFinder_1_io_Stationary_matrix_7_0),
    .io_Stationary_matrix_7_1(PathFinder_1_io_Stationary_matrix_7_1),
    .io_Stationary_matrix_7_2(PathFinder_1_io_Stationary_matrix_7_2),
    .io_Stationary_matrix_7_3(PathFinder_1_io_Stationary_matrix_7_3),
    .io_Stationary_matrix_7_4(PathFinder_1_io_Stationary_matrix_7_4),
    .io_Stationary_matrix_7_5(PathFinder_1_io_Stationary_matrix_7_5),
    .io_Stationary_matrix_7_6(PathFinder_1_io_Stationary_matrix_7_6),
    .io_Stationary_matrix_7_7(PathFinder_1_io_Stationary_matrix_7_7),
    .io_Streaming_matrix_0(PathFinder_1_io_Streaming_matrix_0),
    .io_Streaming_matrix_1(PathFinder_1_io_Streaming_matrix_1),
    .io_Streaming_matrix_2(PathFinder_1_io_Streaming_matrix_2),
    .io_Streaming_matrix_3(PathFinder_1_io_Streaming_matrix_3),
    .io_Streaming_matrix_4(PathFinder_1_io_Streaming_matrix_4),
    .io_Streaming_matrix_5(PathFinder_1_io_Streaming_matrix_5),
    .io_Streaming_matrix_6(PathFinder_1_io_Streaming_matrix_6),
    .io_Streaming_matrix_7(PathFinder_1_io_Streaming_matrix_7),
    .io_i_mux_bus_0(PathFinder_1_io_i_mux_bus_0),
    .io_i_mux_bus_1(PathFinder_1_io_i_mux_bus_1),
    .io_i_mux_bus_2(PathFinder_1_io_i_mux_bus_2),
    .io_i_mux_bus_3(PathFinder_1_io_i_mux_bus_3),
    .io_Source_0(PathFinder_1_io_Source_0),
    .io_Source_1(PathFinder_1_io_Source_1),
    .io_Source_2(PathFinder_1_io_Source_2),
    .io_Source_3(PathFinder_1_io_Source_3),
    .io_destination_0(PathFinder_1_io_destination_0),
    .io_destination_1(PathFinder_1_io_destination_1),
    .io_destination_2(PathFinder_1_io_destination_2),
    .io_destination_3(PathFinder_1_io_destination_3),
    .io_PF_Valid(PathFinder_1_io_PF_Valid),
    .io_NoDPE(PathFinder_1_io_NoDPE),
    .io_DataValid(PathFinder_1_io_DataValid)
  );
  PathFinder PathFinder_2 ( // @[FlexDPU.scala 77:41]
    .clock(PathFinder_2_clock),
    .reset(PathFinder_2_reset),
    .io_Stationary_matrix_0_0(PathFinder_2_io_Stationary_matrix_0_0),
    .io_Stationary_matrix_0_1(PathFinder_2_io_Stationary_matrix_0_1),
    .io_Stationary_matrix_0_2(PathFinder_2_io_Stationary_matrix_0_2),
    .io_Stationary_matrix_0_3(PathFinder_2_io_Stationary_matrix_0_3),
    .io_Stationary_matrix_0_4(PathFinder_2_io_Stationary_matrix_0_4),
    .io_Stationary_matrix_0_5(PathFinder_2_io_Stationary_matrix_0_5),
    .io_Stationary_matrix_0_6(PathFinder_2_io_Stationary_matrix_0_6),
    .io_Stationary_matrix_0_7(PathFinder_2_io_Stationary_matrix_0_7),
    .io_Stationary_matrix_1_0(PathFinder_2_io_Stationary_matrix_1_0),
    .io_Stationary_matrix_1_1(PathFinder_2_io_Stationary_matrix_1_1),
    .io_Stationary_matrix_1_2(PathFinder_2_io_Stationary_matrix_1_2),
    .io_Stationary_matrix_1_3(PathFinder_2_io_Stationary_matrix_1_3),
    .io_Stationary_matrix_1_4(PathFinder_2_io_Stationary_matrix_1_4),
    .io_Stationary_matrix_1_5(PathFinder_2_io_Stationary_matrix_1_5),
    .io_Stationary_matrix_1_6(PathFinder_2_io_Stationary_matrix_1_6),
    .io_Stationary_matrix_1_7(PathFinder_2_io_Stationary_matrix_1_7),
    .io_Stationary_matrix_2_0(PathFinder_2_io_Stationary_matrix_2_0),
    .io_Stationary_matrix_2_1(PathFinder_2_io_Stationary_matrix_2_1),
    .io_Stationary_matrix_2_2(PathFinder_2_io_Stationary_matrix_2_2),
    .io_Stationary_matrix_2_3(PathFinder_2_io_Stationary_matrix_2_3),
    .io_Stationary_matrix_2_4(PathFinder_2_io_Stationary_matrix_2_4),
    .io_Stationary_matrix_2_5(PathFinder_2_io_Stationary_matrix_2_5),
    .io_Stationary_matrix_2_6(PathFinder_2_io_Stationary_matrix_2_6),
    .io_Stationary_matrix_2_7(PathFinder_2_io_Stationary_matrix_2_7),
    .io_Stationary_matrix_3_0(PathFinder_2_io_Stationary_matrix_3_0),
    .io_Stationary_matrix_3_1(PathFinder_2_io_Stationary_matrix_3_1),
    .io_Stationary_matrix_3_2(PathFinder_2_io_Stationary_matrix_3_2),
    .io_Stationary_matrix_3_3(PathFinder_2_io_Stationary_matrix_3_3),
    .io_Stationary_matrix_3_4(PathFinder_2_io_Stationary_matrix_3_4),
    .io_Stationary_matrix_3_5(PathFinder_2_io_Stationary_matrix_3_5),
    .io_Stationary_matrix_3_6(PathFinder_2_io_Stationary_matrix_3_6),
    .io_Stationary_matrix_3_7(PathFinder_2_io_Stationary_matrix_3_7),
    .io_Stationary_matrix_4_0(PathFinder_2_io_Stationary_matrix_4_0),
    .io_Stationary_matrix_4_1(PathFinder_2_io_Stationary_matrix_4_1),
    .io_Stationary_matrix_4_2(PathFinder_2_io_Stationary_matrix_4_2),
    .io_Stationary_matrix_4_3(PathFinder_2_io_Stationary_matrix_4_3),
    .io_Stationary_matrix_4_4(PathFinder_2_io_Stationary_matrix_4_4),
    .io_Stationary_matrix_4_5(PathFinder_2_io_Stationary_matrix_4_5),
    .io_Stationary_matrix_4_6(PathFinder_2_io_Stationary_matrix_4_6),
    .io_Stationary_matrix_4_7(PathFinder_2_io_Stationary_matrix_4_7),
    .io_Stationary_matrix_5_0(PathFinder_2_io_Stationary_matrix_5_0),
    .io_Stationary_matrix_5_1(PathFinder_2_io_Stationary_matrix_5_1),
    .io_Stationary_matrix_5_2(PathFinder_2_io_Stationary_matrix_5_2),
    .io_Stationary_matrix_5_3(PathFinder_2_io_Stationary_matrix_5_3),
    .io_Stationary_matrix_5_4(PathFinder_2_io_Stationary_matrix_5_4),
    .io_Stationary_matrix_5_5(PathFinder_2_io_Stationary_matrix_5_5),
    .io_Stationary_matrix_5_6(PathFinder_2_io_Stationary_matrix_5_6),
    .io_Stationary_matrix_5_7(PathFinder_2_io_Stationary_matrix_5_7),
    .io_Stationary_matrix_6_0(PathFinder_2_io_Stationary_matrix_6_0),
    .io_Stationary_matrix_6_1(PathFinder_2_io_Stationary_matrix_6_1),
    .io_Stationary_matrix_6_2(PathFinder_2_io_Stationary_matrix_6_2),
    .io_Stationary_matrix_6_3(PathFinder_2_io_Stationary_matrix_6_3),
    .io_Stationary_matrix_6_4(PathFinder_2_io_Stationary_matrix_6_4),
    .io_Stationary_matrix_6_5(PathFinder_2_io_Stationary_matrix_6_5),
    .io_Stationary_matrix_6_6(PathFinder_2_io_Stationary_matrix_6_6),
    .io_Stationary_matrix_6_7(PathFinder_2_io_Stationary_matrix_6_7),
    .io_Stationary_matrix_7_0(PathFinder_2_io_Stationary_matrix_7_0),
    .io_Stationary_matrix_7_1(PathFinder_2_io_Stationary_matrix_7_1),
    .io_Stationary_matrix_7_2(PathFinder_2_io_Stationary_matrix_7_2),
    .io_Stationary_matrix_7_3(PathFinder_2_io_Stationary_matrix_7_3),
    .io_Stationary_matrix_7_4(PathFinder_2_io_Stationary_matrix_7_4),
    .io_Stationary_matrix_7_5(PathFinder_2_io_Stationary_matrix_7_5),
    .io_Stationary_matrix_7_6(PathFinder_2_io_Stationary_matrix_7_6),
    .io_Stationary_matrix_7_7(PathFinder_2_io_Stationary_matrix_7_7),
    .io_Streaming_matrix_0(PathFinder_2_io_Streaming_matrix_0),
    .io_Streaming_matrix_1(PathFinder_2_io_Streaming_matrix_1),
    .io_Streaming_matrix_2(PathFinder_2_io_Streaming_matrix_2),
    .io_Streaming_matrix_3(PathFinder_2_io_Streaming_matrix_3),
    .io_Streaming_matrix_4(PathFinder_2_io_Streaming_matrix_4),
    .io_Streaming_matrix_5(PathFinder_2_io_Streaming_matrix_5),
    .io_Streaming_matrix_6(PathFinder_2_io_Streaming_matrix_6),
    .io_Streaming_matrix_7(PathFinder_2_io_Streaming_matrix_7),
    .io_i_mux_bus_0(PathFinder_2_io_i_mux_bus_0),
    .io_i_mux_bus_1(PathFinder_2_io_i_mux_bus_1),
    .io_i_mux_bus_2(PathFinder_2_io_i_mux_bus_2),
    .io_i_mux_bus_3(PathFinder_2_io_i_mux_bus_3),
    .io_Source_0(PathFinder_2_io_Source_0),
    .io_Source_1(PathFinder_2_io_Source_1),
    .io_Source_2(PathFinder_2_io_Source_2),
    .io_Source_3(PathFinder_2_io_Source_3),
    .io_destination_0(PathFinder_2_io_destination_0),
    .io_destination_1(PathFinder_2_io_destination_1),
    .io_destination_2(PathFinder_2_io_destination_2),
    .io_destination_3(PathFinder_2_io_destination_3),
    .io_PF_Valid(PathFinder_2_io_PF_Valid),
    .io_NoDPE(PathFinder_2_io_NoDPE),
    .io_DataValid(PathFinder_2_io_DataValid)
  );
  PathFinder PathFinder_3 ( // @[FlexDPU.scala 77:41]
    .clock(PathFinder_3_clock),
    .reset(PathFinder_3_reset),
    .io_Stationary_matrix_0_0(PathFinder_3_io_Stationary_matrix_0_0),
    .io_Stationary_matrix_0_1(PathFinder_3_io_Stationary_matrix_0_1),
    .io_Stationary_matrix_0_2(PathFinder_3_io_Stationary_matrix_0_2),
    .io_Stationary_matrix_0_3(PathFinder_3_io_Stationary_matrix_0_3),
    .io_Stationary_matrix_0_4(PathFinder_3_io_Stationary_matrix_0_4),
    .io_Stationary_matrix_0_5(PathFinder_3_io_Stationary_matrix_0_5),
    .io_Stationary_matrix_0_6(PathFinder_3_io_Stationary_matrix_0_6),
    .io_Stationary_matrix_0_7(PathFinder_3_io_Stationary_matrix_0_7),
    .io_Stationary_matrix_1_0(PathFinder_3_io_Stationary_matrix_1_0),
    .io_Stationary_matrix_1_1(PathFinder_3_io_Stationary_matrix_1_1),
    .io_Stationary_matrix_1_2(PathFinder_3_io_Stationary_matrix_1_2),
    .io_Stationary_matrix_1_3(PathFinder_3_io_Stationary_matrix_1_3),
    .io_Stationary_matrix_1_4(PathFinder_3_io_Stationary_matrix_1_4),
    .io_Stationary_matrix_1_5(PathFinder_3_io_Stationary_matrix_1_5),
    .io_Stationary_matrix_1_6(PathFinder_3_io_Stationary_matrix_1_6),
    .io_Stationary_matrix_1_7(PathFinder_3_io_Stationary_matrix_1_7),
    .io_Stationary_matrix_2_0(PathFinder_3_io_Stationary_matrix_2_0),
    .io_Stationary_matrix_2_1(PathFinder_3_io_Stationary_matrix_2_1),
    .io_Stationary_matrix_2_2(PathFinder_3_io_Stationary_matrix_2_2),
    .io_Stationary_matrix_2_3(PathFinder_3_io_Stationary_matrix_2_3),
    .io_Stationary_matrix_2_4(PathFinder_3_io_Stationary_matrix_2_4),
    .io_Stationary_matrix_2_5(PathFinder_3_io_Stationary_matrix_2_5),
    .io_Stationary_matrix_2_6(PathFinder_3_io_Stationary_matrix_2_6),
    .io_Stationary_matrix_2_7(PathFinder_3_io_Stationary_matrix_2_7),
    .io_Stationary_matrix_3_0(PathFinder_3_io_Stationary_matrix_3_0),
    .io_Stationary_matrix_3_1(PathFinder_3_io_Stationary_matrix_3_1),
    .io_Stationary_matrix_3_2(PathFinder_3_io_Stationary_matrix_3_2),
    .io_Stationary_matrix_3_3(PathFinder_3_io_Stationary_matrix_3_3),
    .io_Stationary_matrix_3_4(PathFinder_3_io_Stationary_matrix_3_4),
    .io_Stationary_matrix_3_5(PathFinder_3_io_Stationary_matrix_3_5),
    .io_Stationary_matrix_3_6(PathFinder_3_io_Stationary_matrix_3_6),
    .io_Stationary_matrix_3_7(PathFinder_3_io_Stationary_matrix_3_7),
    .io_Stationary_matrix_4_0(PathFinder_3_io_Stationary_matrix_4_0),
    .io_Stationary_matrix_4_1(PathFinder_3_io_Stationary_matrix_4_1),
    .io_Stationary_matrix_4_2(PathFinder_3_io_Stationary_matrix_4_2),
    .io_Stationary_matrix_4_3(PathFinder_3_io_Stationary_matrix_4_3),
    .io_Stationary_matrix_4_4(PathFinder_3_io_Stationary_matrix_4_4),
    .io_Stationary_matrix_4_5(PathFinder_3_io_Stationary_matrix_4_5),
    .io_Stationary_matrix_4_6(PathFinder_3_io_Stationary_matrix_4_6),
    .io_Stationary_matrix_4_7(PathFinder_3_io_Stationary_matrix_4_7),
    .io_Stationary_matrix_5_0(PathFinder_3_io_Stationary_matrix_5_0),
    .io_Stationary_matrix_5_1(PathFinder_3_io_Stationary_matrix_5_1),
    .io_Stationary_matrix_5_2(PathFinder_3_io_Stationary_matrix_5_2),
    .io_Stationary_matrix_5_3(PathFinder_3_io_Stationary_matrix_5_3),
    .io_Stationary_matrix_5_4(PathFinder_3_io_Stationary_matrix_5_4),
    .io_Stationary_matrix_5_5(PathFinder_3_io_Stationary_matrix_5_5),
    .io_Stationary_matrix_5_6(PathFinder_3_io_Stationary_matrix_5_6),
    .io_Stationary_matrix_5_7(PathFinder_3_io_Stationary_matrix_5_7),
    .io_Stationary_matrix_6_0(PathFinder_3_io_Stationary_matrix_6_0),
    .io_Stationary_matrix_6_1(PathFinder_3_io_Stationary_matrix_6_1),
    .io_Stationary_matrix_6_2(PathFinder_3_io_Stationary_matrix_6_2),
    .io_Stationary_matrix_6_3(PathFinder_3_io_Stationary_matrix_6_3),
    .io_Stationary_matrix_6_4(PathFinder_3_io_Stationary_matrix_6_4),
    .io_Stationary_matrix_6_5(PathFinder_3_io_Stationary_matrix_6_5),
    .io_Stationary_matrix_6_6(PathFinder_3_io_Stationary_matrix_6_6),
    .io_Stationary_matrix_6_7(PathFinder_3_io_Stationary_matrix_6_7),
    .io_Stationary_matrix_7_0(PathFinder_3_io_Stationary_matrix_7_0),
    .io_Stationary_matrix_7_1(PathFinder_3_io_Stationary_matrix_7_1),
    .io_Stationary_matrix_7_2(PathFinder_3_io_Stationary_matrix_7_2),
    .io_Stationary_matrix_7_3(PathFinder_3_io_Stationary_matrix_7_3),
    .io_Stationary_matrix_7_4(PathFinder_3_io_Stationary_matrix_7_4),
    .io_Stationary_matrix_7_5(PathFinder_3_io_Stationary_matrix_7_5),
    .io_Stationary_matrix_7_6(PathFinder_3_io_Stationary_matrix_7_6),
    .io_Stationary_matrix_7_7(PathFinder_3_io_Stationary_matrix_7_7),
    .io_Streaming_matrix_0(PathFinder_3_io_Streaming_matrix_0),
    .io_Streaming_matrix_1(PathFinder_3_io_Streaming_matrix_1),
    .io_Streaming_matrix_2(PathFinder_3_io_Streaming_matrix_2),
    .io_Streaming_matrix_3(PathFinder_3_io_Streaming_matrix_3),
    .io_Streaming_matrix_4(PathFinder_3_io_Streaming_matrix_4),
    .io_Streaming_matrix_5(PathFinder_3_io_Streaming_matrix_5),
    .io_Streaming_matrix_6(PathFinder_3_io_Streaming_matrix_6),
    .io_Streaming_matrix_7(PathFinder_3_io_Streaming_matrix_7),
    .io_i_mux_bus_0(PathFinder_3_io_i_mux_bus_0),
    .io_i_mux_bus_1(PathFinder_3_io_i_mux_bus_1),
    .io_i_mux_bus_2(PathFinder_3_io_i_mux_bus_2),
    .io_i_mux_bus_3(PathFinder_3_io_i_mux_bus_3),
    .io_Source_0(PathFinder_3_io_Source_0),
    .io_Source_1(PathFinder_3_io_Source_1),
    .io_Source_2(PathFinder_3_io_Source_2),
    .io_Source_3(PathFinder_3_io_Source_3),
    .io_destination_0(PathFinder_3_io_destination_0),
    .io_destination_1(PathFinder_3_io_destination_1),
    .io_destination_2(PathFinder_3_io_destination_2),
    .io_destination_3(PathFinder_3_io_destination_3),
    .io_PF_Valid(PathFinder_3_io_PF_Valid),
    .io_NoDPE(PathFinder_3_io_NoDPE),
    .io_DataValid(PathFinder_3_io_DataValid)
  );
  PathFinder PathFinder_4 ( // @[FlexDPU.scala 77:41]
    .clock(PathFinder_4_clock),
    .reset(PathFinder_4_reset),
    .io_Stationary_matrix_0_0(PathFinder_4_io_Stationary_matrix_0_0),
    .io_Stationary_matrix_0_1(PathFinder_4_io_Stationary_matrix_0_1),
    .io_Stationary_matrix_0_2(PathFinder_4_io_Stationary_matrix_0_2),
    .io_Stationary_matrix_0_3(PathFinder_4_io_Stationary_matrix_0_3),
    .io_Stationary_matrix_0_4(PathFinder_4_io_Stationary_matrix_0_4),
    .io_Stationary_matrix_0_5(PathFinder_4_io_Stationary_matrix_0_5),
    .io_Stationary_matrix_0_6(PathFinder_4_io_Stationary_matrix_0_6),
    .io_Stationary_matrix_0_7(PathFinder_4_io_Stationary_matrix_0_7),
    .io_Stationary_matrix_1_0(PathFinder_4_io_Stationary_matrix_1_0),
    .io_Stationary_matrix_1_1(PathFinder_4_io_Stationary_matrix_1_1),
    .io_Stationary_matrix_1_2(PathFinder_4_io_Stationary_matrix_1_2),
    .io_Stationary_matrix_1_3(PathFinder_4_io_Stationary_matrix_1_3),
    .io_Stationary_matrix_1_4(PathFinder_4_io_Stationary_matrix_1_4),
    .io_Stationary_matrix_1_5(PathFinder_4_io_Stationary_matrix_1_5),
    .io_Stationary_matrix_1_6(PathFinder_4_io_Stationary_matrix_1_6),
    .io_Stationary_matrix_1_7(PathFinder_4_io_Stationary_matrix_1_7),
    .io_Stationary_matrix_2_0(PathFinder_4_io_Stationary_matrix_2_0),
    .io_Stationary_matrix_2_1(PathFinder_4_io_Stationary_matrix_2_1),
    .io_Stationary_matrix_2_2(PathFinder_4_io_Stationary_matrix_2_2),
    .io_Stationary_matrix_2_3(PathFinder_4_io_Stationary_matrix_2_3),
    .io_Stationary_matrix_2_4(PathFinder_4_io_Stationary_matrix_2_4),
    .io_Stationary_matrix_2_5(PathFinder_4_io_Stationary_matrix_2_5),
    .io_Stationary_matrix_2_6(PathFinder_4_io_Stationary_matrix_2_6),
    .io_Stationary_matrix_2_7(PathFinder_4_io_Stationary_matrix_2_7),
    .io_Stationary_matrix_3_0(PathFinder_4_io_Stationary_matrix_3_0),
    .io_Stationary_matrix_3_1(PathFinder_4_io_Stationary_matrix_3_1),
    .io_Stationary_matrix_3_2(PathFinder_4_io_Stationary_matrix_3_2),
    .io_Stationary_matrix_3_3(PathFinder_4_io_Stationary_matrix_3_3),
    .io_Stationary_matrix_3_4(PathFinder_4_io_Stationary_matrix_3_4),
    .io_Stationary_matrix_3_5(PathFinder_4_io_Stationary_matrix_3_5),
    .io_Stationary_matrix_3_6(PathFinder_4_io_Stationary_matrix_3_6),
    .io_Stationary_matrix_3_7(PathFinder_4_io_Stationary_matrix_3_7),
    .io_Stationary_matrix_4_0(PathFinder_4_io_Stationary_matrix_4_0),
    .io_Stationary_matrix_4_1(PathFinder_4_io_Stationary_matrix_4_1),
    .io_Stationary_matrix_4_2(PathFinder_4_io_Stationary_matrix_4_2),
    .io_Stationary_matrix_4_3(PathFinder_4_io_Stationary_matrix_4_3),
    .io_Stationary_matrix_4_4(PathFinder_4_io_Stationary_matrix_4_4),
    .io_Stationary_matrix_4_5(PathFinder_4_io_Stationary_matrix_4_5),
    .io_Stationary_matrix_4_6(PathFinder_4_io_Stationary_matrix_4_6),
    .io_Stationary_matrix_4_7(PathFinder_4_io_Stationary_matrix_4_7),
    .io_Stationary_matrix_5_0(PathFinder_4_io_Stationary_matrix_5_0),
    .io_Stationary_matrix_5_1(PathFinder_4_io_Stationary_matrix_5_1),
    .io_Stationary_matrix_5_2(PathFinder_4_io_Stationary_matrix_5_2),
    .io_Stationary_matrix_5_3(PathFinder_4_io_Stationary_matrix_5_3),
    .io_Stationary_matrix_5_4(PathFinder_4_io_Stationary_matrix_5_4),
    .io_Stationary_matrix_5_5(PathFinder_4_io_Stationary_matrix_5_5),
    .io_Stationary_matrix_5_6(PathFinder_4_io_Stationary_matrix_5_6),
    .io_Stationary_matrix_5_7(PathFinder_4_io_Stationary_matrix_5_7),
    .io_Stationary_matrix_6_0(PathFinder_4_io_Stationary_matrix_6_0),
    .io_Stationary_matrix_6_1(PathFinder_4_io_Stationary_matrix_6_1),
    .io_Stationary_matrix_6_2(PathFinder_4_io_Stationary_matrix_6_2),
    .io_Stationary_matrix_6_3(PathFinder_4_io_Stationary_matrix_6_3),
    .io_Stationary_matrix_6_4(PathFinder_4_io_Stationary_matrix_6_4),
    .io_Stationary_matrix_6_5(PathFinder_4_io_Stationary_matrix_6_5),
    .io_Stationary_matrix_6_6(PathFinder_4_io_Stationary_matrix_6_6),
    .io_Stationary_matrix_6_7(PathFinder_4_io_Stationary_matrix_6_7),
    .io_Stationary_matrix_7_0(PathFinder_4_io_Stationary_matrix_7_0),
    .io_Stationary_matrix_7_1(PathFinder_4_io_Stationary_matrix_7_1),
    .io_Stationary_matrix_7_2(PathFinder_4_io_Stationary_matrix_7_2),
    .io_Stationary_matrix_7_3(PathFinder_4_io_Stationary_matrix_7_3),
    .io_Stationary_matrix_7_4(PathFinder_4_io_Stationary_matrix_7_4),
    .io_Stationary_matrix_7_5(PathFinder_4_io_Stationary_matrix_7_5),
    .io_Stationary_matrix_7_6(PathFinder_4_io_Stationary_matrix_7_6),
    .io_Stationary_matrix_7_7(PathFinder_4_io_Stationary_matrix_7_7),
    .io_Streaming_matrix_0(PathFinder_4_io_Streaming_matrix_0),
    .io_Streaming_matrix_1(PathFinder_4_io_Streaming_matrix_1),
    .io_Streaming_matrix_2(PathFinder_4_io_Streaming_matrix_2),
    .io_Streaming_matrix_3(PathFinder_4_io_Streaming_matrix_3),
    .io_Streaming_matrix_4(PathFinder_4_io_Streaming_matrix_4),
    .io_Streaming_matrix_5(PathFinder_4_io_Streaming_matrix_5),
    .io_Streaming_matrix_6(PathFinder_4_io_Streaming_matrix_6),
    .io_Streaming_matrix_7(PathFinder_4_io_Streaming_matrix_7),
    .io_i_mux_bus_0(PathFinder_4_io_i_mux_bus_0),
    .io_i_mux_bus_1(PathFinder_4_io_i_mux_bus_1),
    .io_i_mux_bus_2(PathFinder_4_io_i_mux_bus_2),
    .io_i_mux_bus_3(PathFinder_4_io_i_mux_bus_3),
    .io_Source_0(PathFinder_4_io_Source_0),
    .io_Source_1(PathFinder_4_io_Source_1),
    .io_Source_2(PathFinder_4_io_Source_2),
    .io_Source_3(PathFinder_4_io_Source_3),
    .io_destination_0(PathFinder_4_io_destination_0),
    .io_destination_1(PathFinder_4_io_destination_1),
    .io_destination_2(PathFinder_4_io_destination_2),
    .io_destination_3(PathFinder_4_io_destination_3),
    .io_PF_Valid(PathFinder_4_io_PF_Valid),
    .io_NoDPE(PathFinder_4_io_NoDPE),
    .io_DataValid(PathFinder_4_io_DataValid)
  );
  PathFinder PathFinder_5 ( // @[FlexDPU.scala 77:41]
    .clock(PathFinder_5_clock),
    .reset(PathFinder_5_reset),
    .io_Stationary_matrix_0_0(PathFinder_5_io_Stationary_matrix_0_0),
    .io_Stationary_matrix_0_1(PathFinder_5_io_Stationary_matrix_0_1),
    .io_Stationary_matrix_0_2(PathFinder_5_io_Stationary_matrix_0_2),
    .io_Stationary_matrix_0_3(PathFinder_5_io_Stationary_matrix_0_3),
    .io_Stationary_matrix_0_4(PathFinder_5_io_Stationary_matrix_0_4),
    .io_Stationary_matrix_0_5(PathFinder_5_io_Stationary_matrix_0_5),
    .io_Stationary_matrix_0_6(PathFinder_5_io_Stationary_matrix_0_6),
    .io_Stationary_matrix_0_7(PathFinder_5_io_Stationary_matrix_0_7),
    .io_Stationary_matrix_1_0(PathFinder_5_io_Stationary_matrix_1_0),
    .io_Stationary_matrix_1_1(PathFinder_5_io_Stationary_matrix_1_1),
    .io_Stationary_matrix_1_2(PathFinder_5_io_Stationary_matrix_1_2),
    .io_Stationary_matrix_1_3(PathFinder_5_io_Stationary_matrix_1_3),
    .io_Stationary_matrix_1_4(PathFinder_5_io_Stationary_matrix_1_4),
    .io_Stationary_matrix_1_5(PathFinder_5_io_Stationary_matrix_1_5),
    .io_Stationary_matrix_1_6(PathFinder_5_io_Stationary_matrix_1_6),
    .io_Stationary_matrix_1_7(PathFinder_5_io_Stationary_matrix_1_7),
    .io_Stationary_matrix_2_0(PathFinder_5_io_Stationary_matrix_2_0),
    .io_Stationary_matrix_2_1(PathFinder_5_io_Stationary_matrix_2_1),
    .io_Stationary_matrix_2_2(PathFinder_5_io_Stationary_matrix_2_2),
    .io_Stationary_matrix_2_3(PathFinder_5_io_Stationary_matrix_2_3),
    .io_Stationary_matrix_2_4(PathFinder_5_io_Stationary_matrix_2_4),
    .io_Stationary_matrix_2_5(PathFinder_5_io_Stationary_matrix_2_5),
    .io_Stationary_matrix_2_6(PathFinder_5_io_Stationary_matrix_2_6),
    .io_Stationary_matrix_2_7(PathFinder_5_io_Stationary_matrix_2_7),
    .io_Stationary_matrix_3_0(PathFinder_5_io_Stationary_matrix_3_0),
    .io_Stationary_matrix_3_1(PathFinder_5_io_Stationary_matrix_3_1),
    .io_Stationary_matrix_3_2(PathFinder_5_io_Stationary_matrix_3_2),
    .io_Stationary_matrix_3_3(PathFinder_5_io_Stationary_matrix_3_3),
    .io_Stationary_matrix_3_4(PathFinder_5_io_Stationary_matrix_3_4),
    .io_Stationary_matrix_3_5(PathFinder_5_io_Stationary_matrix_3_5),
    .io_Stationary_matrix_3_6(PathFinder_5_io_Stationary_matrix_3_6),
    .io_Stationary_matrix_3_7(PathFinder_5_io_Stationary_matrix_3_7),
    .io_Stationary_matrix_4_0(PathFinder_5_io_Stationary_matrix_4_0),
    .io_Stationary_matrix_4_1(PathFinder_5_io_Stationary_matrix_4_1),
    .io_Stationary_matrix_4_2(PathFinder_5_io_Stationary_matrix_4_2),
    .io_Stationary_matrix_4_3(PathFinder_5_io_Stationary_matrix_4_3),
    .io_Stationary_matrix_4_4(PathFinder_5_io_Stationary_matrix_4_4),
    .io_Stationary_matrix_4_5(PathFinder_5_io_Stationary_matrix_4_5),
    .io_Stationary_matrix_4_6(PathFinder_5_io_Stationary_matrix_4_6),
    .io_Stationary_matrix_4_7(PathFinder_5_io_Stationary_matrix_4_7),
    .io_Stationary_matrix_5_0(PathFinder_5_io_Stationary_matrix_5_0),
    .io_Stationary_matrix_5_1(PathFinder_5_io_Stationary_matrix_5_1),
    .io_Stationary_matrix_5_2(PathFinder_5_io_Stationary_matrix_5_2),
    .io_Stationary_matrix_5_3(PathFinder_5_io_Stationary_matrix_5_3),
    .io_Stationary_matrix_5_4(PathFinder_5_io_Stationary_matrix_5_4),
    .io_Stationary_matrix_5_5(PathFinder_5_io_Stationary_matrix_5_5),
    .io_Stationary_matrix_5_6(PathFinder_5_io_Stationary_matrix_5_6),
    .io_Stationary_matrix_5_7(PathFinder_5_io_Stationary_matrix_5_7),
    .io_Stationary_matrix_6_0(PathFinder_5_io_Stationary_matrix_6_0),
    .io_Stationary_matrix_6_1(PathFinder_5_io_Stationary_matrix_6_1),
    .io_Stationary_matrix_6_2(PathFinder_5_io_Stationary_matrix_6_2),
    .io_Stationary_matrix_6_3(PathFinder_5_io_Stationary_matrix_6_3),
    .io_Stationary_matrix_6_4(PathFinder_5_io_Stationary_matrix_6_4),
    .io_Stationary_matrix_6_5(PathFinder_5_io_Stationary_matrix_6_5),
    .io_Stationary_matrix_6_6(PathFinder_5_io_Stationary_matrix_6_6),
    .io_Stationary_matrix_6_7(PathFinder_5_io_Stationary_matrix_6_7),
    .io_Stationary_matrix_7_0(PathFinder_5_io_Stationary_matrix_7_0),
    .io_Stationary_matrix_7_1(PathFinder_5_io_Stationary_matrix_7_1),
    .io_Stationary_matrix_7_2(PathFinder_5_io_Stationary_matrix_7_2),
    .io_Stationary_matrix_7_3(PathFinder_5_io_Stationary_matrix_7_3),
    .io_Stationary_matrix_7_4(PathFinder_5_io_Stationary_matrix_7_4),
    .io_Stationary_matrix_7_5(PathFinder_5_io_Stationary_matrix_7_5),
    .io_Stationary_matrix_7_6(PathFinder_5_io_Stationary_matrix_7_6),
    .io_Stationary_matrix_7_7(PathFinder_5_io_Stationary_matrix_7_7),
    .io_Streaming_matrix_0(PathFinder_5_io_Streaming_matrix_0),
    .io_Streaming_matrix_1(PathFinder_5_io_Streaming_matrix_1),
    .io_Streaming_matrix_2(PathFinder_5_io_Streaming_matrix_2),
    .io_Streaming_matrix_3(PathFinder_5_io_Streaming_matrix_3),
    .io_Streaming_matrix_4(PathFinder_5_io_Streaming_matrix_4),
    .io_Streaming_matrix_5(PathFinder_5_io_Streaming_matrix_5),
    .io_Streaming_matrix_6(PathFinder_5_io_Streaming_matrix_6),
    .io_Streaming_matrix_7(PathFinder_5_io_Streaming_matrix_7),
    .io_i_mux_bus_0(PathFinder_5_io_i_mux_bus_0),
    .io_i_mux_bus_1(PathFinder_5_io_i_mux_bus_1),
    .io_i_mux_bus_2(PathFinder_5_io_i_mux_bus_2),
    .io_i_mux_bus_3(PathFinder_5_io_i_mux_bus_3),
    .io_Source_0(PathFinder_5_io_Source_0),
    .io_Source_1(PathFinder_5_io_Source_1),
    .io_Source_2(PathFinder_5_io_Source_2),
    .io_Source_3(PathFinder_5_io_Source_3),
    .io_destination_0(PathFinder_5_io_destination_0),
    .io_destination_1(PathFinder_5_io_destination_1),
    .io_destination_2(PathFinder_5_io_destination_2),
    .io_destination_3(PathFinder_5_io_destination_3),
    .io_PF_Valid(PathFinder_5_io_PF_Valid),
    .io_NoDPE(PathFinder_5_io_NoDPE),
    .io_DataValid(PathFinder_5_io_DataValid)
  );
  PathFinder PathFinder_6 ( // @[FlexDPU.scala 77:41]
    .clock(PathFinder_6_clock),
    .reset(PathFinder_6_reset),
    .io_Stationary_matrix_0_0(PathFinder_6_io_Stationary_matrix_0_0),
    .io_Stationary_matrix_0_1(PathFinder_6_io_Stationary_matrix_0_1),
    .io_Stationary_matrix_0_2(PathFinder_6_io_Stationary_matrix_0_2),
    .io_Stationary_matrix_0_3(PathFinder_6_io_Stationary_matrix_0_3),
    .io_Stationary_matrix_0_4(PathFinder_6_io_Stationary_matrix_0_4),
    .io_Stationary_matrix_0_5(PathFinder_6_io_Stationary_matrix_0_5),
    .io_Stationary_matrix_0_6(PathFinder_6_io_Stationary_matrix_0_6),
    .io_Stationary_matrix_0_7(PathFinder_6_io_Stationary_matrix_0_7),
    .io_Stationary_matrix_1_0(PathFinder_6_io_Stationary_matrix_1_0),
    .io_Stationary_matrix_1_1(PathFinder_6_io_Stationary_matrix_1_1),
    .io_Stationary_matrix_1_2(PathFinder_6_io_Stationary_matrix_1_2),
    .io_Stationary_matrix_1_3(PathFinder_6_io_Stationary_matrix_1_3),
    .io_Stationary_matrix_1_4(PathFinder_6_io_Stationary_matrix_1_4),
    .io_Stationary_matrix_1_5(PathFinder_6_io_Stationary_matrix_1_5),
    .io_Stationary_matrix_1_6(PathFinder_6_io_Stationary_matrix_1_6),
    .io_Stationary_matrix_1_7(PathFinder_6_io_Stationary_matrix_1_7),
    .io_Stationary_matrix_2_0(PathFinder_6_io_Stationary_matrix_2_0),
    .io_Stationary_matrix_2_1(PathFinder_6_io_Stationary_matrix_2_1),
    .io_Stationary_matrix_2_2(PathFinder_6_io_Stationary_matrix_2_2),
    .io_Stationary_matrix_2_3(PathFinder_6_io_Stationary_matrix_2_3),
    .io_Stationary_matrix_2_4(PathFinder_6_io_Stationary_matrix_2_4),
    .io_Stationary_matrix_2_5(PathFinder_6_io_Stationary_matrix_2_5),
    .io_Stationary_matrix_2_6(PathFinder_6_io_Stationary_matrix_2_6),
    .io_Stationary_matrix_2_7(PathFinder_6_io_Stationary_matrix_2_7),
    .io_Stationary_matrix_3_0(PathFinder_6_io_Stationary_matrix_3_0),
    .io_Stationary_matrix_3_1(PathFinder_6_io_Stationary_matrix_3_1),
    .io_Stationary_matrix_3_2(PathFinder_6_io_Stationary_matrix_3_2),
    .io_Stationary_matrix_3_3(PathFinder_6_io_Stationary_matrix_3_3),
    .io_Stationary_matrix_3_4(PathFinder_6_io_Stationary_matrix_3_4),
    .io_Stationary_matrix_3_5(PathFinder_6_io_Stationary_matrix_3_5),
    .io_Stationary_matrix_3_6(PathFinder_6_io_Stationary_matrix_3_6),
    .io_Stationary_matrix_3_7(PathFinder_6_io_Stationary_matrix_3_7),
    .io_Stationary_matrix_4_0(PathFinder_6_io_Stationary_matrix_4_0),
    .io_Stationary_matrix_4_1(PathFinder_6_io_Stationary_matrix_4_1),
    .io_Stationary_matrix_4_2(PathFinder_6_io_Stationary_matrix_4_2),
    .io_Stationary_matrix_4_3(PathFinder_6_io_Stationary_matrix_4_3),
    .io_Stationary_matrix_4_4(PathFinder_6_io_Stationary_matrix_4_4),
    .io_Stationary_matrix_4_5(PathFinder_6_io_Stationary_matrix_4_5),
    .io_Stationary_matrix_4_6(PathFinder_6_io_Stationary_matrix_4_6),
    .io_Stationary_matrix_4_7(PathFinder_6_io_Stationary_matrix_4_7),
    .io_Stationary_matrix_5_0(PathFinder_6_io_Stationary_matrix_5_0),
    .io_Stationary_matrix_5_1(PathFinder_6_io_Stationary_matrix_5_1),
    .io_Stationary_matrix_5_2(PathFinder_6_io_Stationary_matrix_5_2),
    .io_Stationary_matrix_5_3(PathFinder_6_io_Stationary_matrix_5_3),
    .io_Stationary_matrix_5_4(PathFinder_6_io_Stationary_matrix_5_4),
    .io_Stationary_matrix_5_5(PathFinder_6_io_Stationary_matrix_5_5),
    .io_Stationary_matrix_5_6(PathFinder_6_io_Stationary_matrix_5_6),
    .io_Stationary_matrix_5_7(PathFinder_6_io_Stationary_matrix_5_7),
    .io_Stationary_matrix_6_0(PathFinder_6_io_Stationary_matrix_6_0),
    .io_Stationary_matrix_6_1(PathFinder_6_io_Stationary_matrix_6_1),
    .io_Stationary_matrix_6_2(PathFinder_6_io_Stationary_matrix_6_2),
    .io_Stationary_matrix_6_3(PathFinder_6_io_Stationary_matrix_6_3),
    .io_Stationary_matrix_6_4(PathFinder_6_io_Stationary_matrix_6_4),
    .io_Stationary_matrix_6_5(PathFinder_6_io_Stationary_matrix_6_5),
    .io_Stationary_matrix_6_6(PathFinder_6_io_Stationary_matrix_6_6),
    .io_Stationary_matrix_6_7(PathFinder_6_io_Stationary_matrix_6_7),
    .io_Stationary_matrix_7_0(PathFinder_6_io_Stationary_matrix_7_0),
    .io_Stationary_matrix_7_1(PathFinder_6_io_Stationary_matrix_7_1),
    .io_Stationary_matrix_7_2(PathFinder_6_io_Stationary_matrix_7_2),
    .io_Stationary_matrix_7_3(PathFinder_6_io_Stationary_matrix_7_3),
    .io_Stationary_matrix_7_4(PathFinder_6_io_Stationary_matrix_7_4),
    .io_Stationary_matrix_7_5(PathFinder_6_io_Stationary_matrix_7_5),
    .io_Stationary_matrix_7_6(PathFinder_6_io_Stationary_matrix_7_6),
    .io_Stationary_matrix_7_7(PathFinder_6_io_Stationary_matrix_7_7),
    .io_Streaming_matrix_0(PathFinder_6_io_Streaming_matrix_0),
    .io_Streaming_matrix_1(PathFinder_6_io_Streaming_matrix_1),
    .io_Streaming_matrix_2(PathFinder_6_io_Streaming_matrix_2),
    .io_Streaming_matrix_3(PathFinder_6_io_Streaming_matrix_3),
    .io_Streaming_matrix_4(PathFinder_6_io_Streaming_matrix_4),
    .io_Streaming_matrix_5(PathFinder_6_io_Streaming_matrix_5),
    .io_Streaming_matrix_6(PathFinder_6_io_Streaming_matrix_6),
    .io_Streaming_matrix_7(PathFinder_6_io_Streaming_matrix_7),
    .io_i_mux_bus_0(PathFinder_6_io_i_mux_bus_0),
    .io_i_mux_bus_1(PathFinder_6_io_i_mux_bus_1),
    .io_i_mux_bus_2(PathFinder_6_io_i_mux_bus_2),
    .io_i_mux_bus_3(PathFinder_6_io_i_mux_bus_3),
    .io_Source_0(PathFinder_6_io_Source_0),
    .io_Source_1(PathFinder_6_io_Source_1),
    .io_Source_2(PathFinder_6_io_Source_2),
    .io_Source_3(PathFinder_6_io_Source_3),
    .io_destination_0(PathFinder_6_io_destination_0),
    .io_destination_1(PathFinder_6_io_destination_1),
    .io_destination_2(PathFinder_6_io_destination_2),
    .io_destination_3(PathFinder_6_io_destination_3),
    .io_PF_Valid(PathFinder_6_io_PF_Valid),
    .io_NoDPE(PathFinder_6_io_NoDPE),
    .io_DataValid(PathFinder_6_io_DataValid)
  );
  PathFinder PathFinder_7 ( // @[FlexDPU.scala 77:41]
    .clock(PathFinder_7_clock),
    .reset(PathFinder_7_reset),
    .io_Stationary_matrix_0_0(PathFinder_7_io_Stationary_matrix_0_0),
    .io_Stationary_matrix_0_1(PathFinder_7_io_Stationary_matrix_0_1),
    .io_Stationary_matrix_0_2(PathFinder_7_io_Stationary_matrix_0_2),
    .io_Stationary_matrix_0_3(PathFinder_7_io_Stationary_matrix_0_3),
    .io_Stationary_matrix_0_4(PathFinder_7_io_Stationary_matrix_0_4),
    .io_Stationary_matrix_0_5(PathFinder_7_io_Stationary_matrix_0_5),
    .io_Stationary_matrix_0_6(PathFinder_7_io_Stationary_matrix_0_6),
    .io_Stationary_matrix_0_7(PathFinder_7_io_Stationary_matrix_0_7),
    .io_Stationary_matrix_1_0(PathFinder_7_io_Stationary_matrix_1_0),
    .io_Stationary_matrix_1_1(PathFinder_7_io_Stationary_matrix_1_1),
    .io_Stationary_matrix_1_2(PathFinder_7_io_Stationary_matrix_1_2),
    .io_Stationary_matrix_1_3(PathFinder_7_io_Stationary_matrix_1_3),
    .io_Stationary_matrix_1_4(PathFinder_7_io_Stationary_matrix_1_4),
    .io_Stationary_matrix_1_5(PathFinder_7_io_Stationary_matrix_1_5),
    .io_Stationary_matrix_1_6(PathFinder_7_io_Stationary_matrix_1_6),
    .io_Stationary_matrix_1_7(PathFinder_7_io_Stationary_matrix_1_7),
    .io_Stationary_matrix_2_0(PathFinder_7_io_Stationary_matrix_2_0),
    .io_Stationary_matrix_2_1(PathFinder_7_io_Stationary_matrix_2_1),
    .io_Stationary_matrix_2_2(PathFinder_7_io_Stationary_matrix_2_2),
    .io_Stationary_matrix_2_3(PathFinder_7_io_Stationary_matrix_2_3),
    .io_Stationary_matrix_2_4(PathFinder_7_io_Stationary_matrix_2_4),
    .io_Stationary_matrix_2_5(PathFinder_7_io_Stationary_matrix_2_5),
    .io_Stationary_matrix_2_6(PathFinder_7_io_Stationary_matrix_2_6),
    .io_Stationary_matrix_2_7(PathFinder_7_io_Stationary_matrix_2_7),
    .io_Stationary_matrix_3_0(PathFinder_7_io_Stationary_matrix_3_0),
    .io_Stationary_matrix_3_1(PathFinder_7_io_Stationary_matrix_3_1),
    .io_Stationary_matrix_3_2(PathFinder_7_io_Stationary_matrix_3_2),
    .io_Stationary_matrix_3_3(PathFinder_7_io_Stationary_matrix_3_3),
    .io_Stationary_matrix_3_4(PathFinder_7_io_Stationary_matrix_3_4),
    .io_Stationary_matrix_3_5(PathFinder_7_io_Stationary_matrix_3_5),
    .io_Stationary_matrix_3_6(PathFinder_7_io_Stationary_matrix_3_6),
    .io_Stationary_matrix_3_7(PathFinder_7_io_Stationary_matrix_3_7),
    .io_Stationary_matrix_4_0(PathFinder_7_io_Stationary_matrix_4_0),
    .io_Stationary_matrix_4_1(PathFinder_7_io_Stationary_matrix_4_1),
    .io_Stationary_matrix_4_2(PathFinder_7_io_Stationary_matrix_4_2),
    .io_Stationary_matrix_4_3(PathFinder_7_io_Stationary_matrix_4_3),
    .io_Stationary_matrix_4_4(PathFinder_7_io_Stationary_matrix_4_4),
    .io_Stationary_matrix_4_5(PathFinder_7_io_Stationary_matrix_4_5),
    .io_Stationary_matrix_4_6(PathFinder_7_io_Stationary_matrix_4_6),
    .io_Stationary_matrix_4_7(PathFinder_7_io_Stationary_matrix_4_7),
    .io_Stationary_matrix_5_0(PathFinder_7_io_Stationary_matrix_5_0),
    .io_Stationary_matrix_5_1(PathFinder_7_io_Stationary_matrix_5_1),
    .io_Stationary_matrix_5_2(PathFinder_7_io_Stationary_matrix_5_2),
    .io_Stationary_matrix_5_3(PathFinder_7_io_Stationary_matrix_5_3),
    .io_Stationary_matrix_5_4(PathFinder_7_io_Stationary_matrix_5_4),
    .io_Stationary_matrix_5_5(PathFinder_7_io_Stationary_matrix_5_5),
    .io_Stationary_matrix_5_6(PathFinder_7_io_Stationary_matrix_5_6),
    .io_Stationary_matrix_5_7(PathFinder_7_io_Stationary_matrix_5_7),
    .io_Stationary_matrix_6_0(PathFinder_7_io_Stationary_matrix_6_0),
    .io_Stationary_matrix_6_1(PathFinder_7_io_Stationary_matrix_6_1),
    .io_Stationary_matrix_6_2(PathFinder_7_io_Stationary_matrix_6_2),
    .io_Stationary_matrix_6_3(PathFinder_7_io_Stationary_matrix_6_3),
    .io_Stationary_matrix_6_4(PathFinder_7_io_Stationary_matrix_6_4),
    .io_Stationary_matrix_6_5(PathFinder_7_io_Stationary_matrix_6_5),
    .io_Stationary_matrix_6_6(PathFinder_7_io_Stationary_matrix_6_6),
    .io_Stationary_matrix_6_7(PathFinder_7_io_Stationary_matrix_6_7),
    .io_Stationary_matrix_7_0(PathFinder_7_io_Stationary_matrix_7_0),
    .io_Stationary_matrix_7_1(PathFinder_7_io_Stationary_matrix_7_1),
    .io_Stationary_matrix_7_2(PathFinder_7_io_Stationary_matrix_7_2),
    .io_Stationary_matrix_7_3(PathFinder_7_io_Stationary_matrix_7_3),
    .io_Stationary_matrix_7_4(PathFinder_7_io_Stationary_matrix_7_4),
    .io_Stationary_matrix_7_5(PathFinder_7_io_Stationary_matrix_7_5),
    .io_Stationary_matrix_7_6(PathFinder_7_io_Stationary_matrix_7_6),
    .io_Stationary_matrix_7_7(PathFinder_7_io_Stationary_matrix_7_7),
    .io_Streaming_matrix_0(PathFinder_7_io_Streaming_matrix_0),
    .io_Streaming_matrix_1(PathFinder_7_io_Streaming_matrix_1),
    .io_Streaming_matrix_2(PathFinder_7_io_Streaming_matrix_2),
    .io_Streaming_matrix_3(PathFinder_7_io_Streaming_matrix_3),
    .io_Streaming_matrix_4(PathFinder_7_io_Streaming_matrix_4),
    .io_Streaming_matrix_5(PathFinder_7_io_Streaming_matrix_5),
    .io_Streaming_matrix_6(PathFinder_7_io_Streaming_matrix_6),
    .io_Streaming_matrix_7(PathFinder_7_io_Streaming_matrix_7),
    .io_i_mux_bus_0(PathFinder_7_io_i_mux_bus_0),
    .io_i_mux_bus_1(PathFinder_7_io_i_mux_bus_1),
    .io_i_mux_bus_2(PathFinder_7_io_i_mux_bus_2),
    .io_i_mux_bus_3(PathFinder_7_io_i_mux_bus_3),
    .io_Source_0(PathFinder_7_io_Source_0),
    .io_Source_1(PathFinder_7_io_Source_1),
    .io_Source_2(PathFinder_7_io_Source_2),
    .io_Source_3(PathFinder_7_io_Source_3),
    .io_destination_0(PathFinder_7_io_destination_0),
    .io_destination_1(PathFinder_7_io_destination_1),
    .io_destination_2(PathFinder_7_io_destination_2),
    .io_destination_3(PathFinder_7_io_destination_3),
    .io_PF_Valid(PathFinder_7_io_PF_Valid),
    .io_NoDPE(PathFinder_7_io_NoDPE),
    .io_DataValid(PathFinder_7_io_DataValid)
  );
  PathFinder PathFinder_8 ( // @[FlexDPU.scala 77:41]
    .clock(PathFinder_8_clock),
    .reset(PathFinder_8_reset),
    .io_Stationary_matrix_0_0(PathFinder_8_io_Stationary_matrix_0_0),
    .io_Stationary_matrix_0_1(PathFinder_8_io_Stationary_matrix_0_1),
    .io_Stationary_matrix_0_2(PathFinder_8_io_Stationary_matrix_0_2),
    .io_Stationary_matrix_0_3(PathFinder_8_io_Stationary_matrix_0_3),
    .io_Stationary_matrix_0_4(PathFinder_8_io_Stationary_matrix_0_4),
    .io_Stationary_matrix_0_5(PathFinder_8_io_Stationary_matrix_0_5),
    .io_Stationary_matrix_0_6(PathFinder_8_io_Stationary_matrix_0_6),
    .io_Stationary_matrix_0_7(PathFinder_8_io_Stationary_matrix_0_7),
    .io_Stationary_matrix_1_0(PathFinder_8_io_Stationary_matrix_1_0),
    .io_Stationary_matrix_1_1(PathFinder_8_io_Stationary_matrix_1_1),
    .io_Stationary_matrix_1_2(PathFinder_8_io_Stationary_matrix_1_2),
    .io_Stationary_matrix_1_3(PathFinder_8_io_Stationary_matrix_1_3),
    .io_Stationary_matrix_1_4(PathFinder_8_io_Stationary_matrix_1_4),
    .io_Stationary_matrix_1_5(PathFinder_8_io_Stationary_matrix_1_5),
    .io_Stationary_matrix_1_6(PathFinder_8_io_Stationary_matrix_1_6),
    .io_Stationary_matrix_1_7(PathFinder_8_io_Stationary_matrix_1_7),
    .io_Stationary_matrix_2_0(PathFinder_8_io_Stationary_matrix_2_0),
    .io_Stationary_matrix_2_1(PathFinder_8_io_Stationary_matrix_2_1),
    .io_Stationary_matrix_2_2(PathFinder_8_io_Stationary_matrix_2_2),
    .io_Stationary_matrix_2_3(PathFinder_8_io_Stationary_matrix_2_3),
    .io_Stationary_matrix_2_4(PathFinder_8_io_Stationary_matrix_2_4),
    .io_Stationary_matrix_2_5(PathFinder_8_io_Stationary_matrix_2_5),
    .io_Stationary_matrix_2_6(PathFinder_8_io_Stationary_matrix_2_6),
    .io_Stationary_matrix_2_7(PathFinder_8_io_Stationary_matrix_2_7),
    .io_Stationary_matrix_3_0(PathFinder_8_io_Stationary_matrix_3_0),
    .io_Stationary_matrix_3_1(PathFinder_8_io_Stationary_matrix_3_1),
    .io_Stationary_matrix_3_2(PathFinder_8_io_Stationary_matrix_3_2),
    .io_Stationary_matrix_3_3(PathFinder_8_io_Stationary_matrix_3_3),
    .io_Stationary_matrix_3_4(PathFinder_8_io_Stationary_matrix_3_4),
    .io_Stationary_matrix_3_5(PathFinder_8_io_Stationary_matrix_3_5),
    .io_Stationary_matrix_3_6(PathFinder_8_io_Stationary_matrix_3_6),
    .io_Stationary_matrix_3_7(PathFinder_8_io_Stationary_matrix_3_7),
    .io_Stationary_matrix_4_0(PathFinder_8_io_Stationary_matrix_4_0),
    .io_Stationary_matrix_4_1(PathFinder_8_io_Stationary_matrix_4_1),
    .io_Stationary_matrix_4_2(PathFinder_8_io_Stationary_matrix_4_2),
    .io_Stationary_matrix_4_3(PathFinder_8_io_Stationary_matrix_4_3),
    .io_Stationary_matrix_4_4(PathFinder_8_io_Stationary_matrix_4_4),
    .io_Stationary_matrix_4_5(PathFinder_8_io_Stationary_matrix_4_5),
    .io_Stationary_matrix_4_6(PathFinder_8_io_Stationary_matrix_4_6),
    .io_Stationary_matrix_4_7(PathFinder_8_io_Stationary_matrix_4_7),
    .io_Stationary_matrix_5_0(PathFinder_8_io_Stationary_matrix_5_0),
    .io_Stationary_matrix_5_1(PathFinder_8_io_Stationary_matrix_5_1),
    .io_Stationary_matrix_5_2(PathFinder_8_io_Stationary_matrix_5_2),
    .io_Stationary_matrix_5_3(PathFinder_8_io_Stationary_matrix_5_3),
    .io_Stationary_matrix_5_4(PathFinder_8_io_Stationary_matrix_5_4),
    .io_Stationary_matrix_5_5(PathFinder_8_io_Stationary_matrix_5_5),
    .io_Stationary_matrix_5_6(PathFinder_8_io_Stationary_matrix_5_6),
    .io_Stationary_matrix_5_7(PathFinder_8_io_Stationary_matrix_5_7),
    .io_Stationary_matrix_6_0(PathFinder_8_io_Stationary_matrix_6_0),
    .io_Stationary_matrix_6_1(PathFinder_8_io_Stationary_matrix_6_1),
    .io_Stationary_matrix_6_2(PathFinder_8_io_Stationary_matrix_6_2),
    .io_Stationary_matrix_6_3(PathFinder_8_io_Stationary_matrix_6_3),
    .io_Stationary_matrix_6_4(PathFinder_8_io_Stationary_matrix_6_4),
    .io_Stationary_matrix_6_5(PathFinder_8_io_Stationary_matrix_6_5),
    .io_Stationary_matrix_6_6(PathFinder_8_io_Stationary_matrix_6_6),
    .io_Stationary_matrix_6_7(PathFinder_8_io_Stationary_matrix_6_7),
    .io_Stationary_matrix_7_0(PathFinder_8_io_Stationary_matrix_7_0),
    .io_Stationary_matrix_7_1(PathFinder_8_io_Stationary_matrix_7_1),
    .io_Stationary_matrix_7_2(PathFinder_8_io_Stationary_matrix_7_2),
    .io_Stationary_matrix_7_3(PathFinder_8_io_Stationary_matrix_7_3),
    .io_Stationary_matrix_7_4(PathFinder_8_io_Stationary_matrix_7_4),
    .io_Stationary_matrix_7_5(PathFinder_8_io_Stationary_matrix_7_5),
    .io_Stationary_matrix_7_6(PathFinder_8_io_Stationary_matrix_7_6),
    .io_Stationary_matrix_7_7(PathFinder_8_io_Stationary_matrix_7_7),
    .io_Streaming_matrix_0(PathFinder_8_io_Streaming_matrix_0),
    .io_Streaming_matrix_1(PathFinder_8_io_Streaming_matrix_1),
    .io_Streaming_matrix_2(PathFinder_8_io_Streaming_matrix_2),
    .io_Streaming_matrix_3(PathFinder_8_io_Streaming_matrix_3),
    .io_Streaming_matrix_4(PathFinder_8_io_Streaming_matrix_4),
    .io_Streaming_matrix_5(PathFinder_8_io_Streaming_matrix_5),
    .io_Streaming_matrix_6(PathFinder_8_io_Streaming_matrix_6),
    .io_Streaming_matrix_7(PathFinder_8_io_Streaming_matrix_7),
    .io_i_mux_bus_0(PathFinder_8_io_i_mux_bus_0),
    .io_i_mux_bus_1(PathFinder_8_io_i_mux_bus_1),
    .io_i_mux_bus_2(PathFinder_8_io_i_mux_bus_2),
    .io_i_mux_bus_3(PathFinder_8_io_i_mux_bus_3),
    .io_Source_0(PathFinder_8_io_Source_0),
    .io_Source_1(PathFinder_8_io_Source_1),
    .io_Source_2(PathFinder_8_io_Source_2),
    .io_Source_3(PathFinder_8_io_Source_3),
    .io_destination_0(PathFinder_8_io_destination_0),
    .io_destination_1(PathFinder_8_io_destination_1),
    .io_destination_2(PathFinder_8_io_destination_2),
    .io_destination_3(PathFinder_8_io_destination_3),
    .io_PF_Valid(PathFinder_8_io_PF_Valid),
    .io_NoDPE(PathFinder_8_io_NoDPE),
    .io_DataValid(PathFinder_8_io_DataValid)
  );
  PathFinder PathFinder_9 ( // @[FlexDPU.scala 77:41]
    .clock(PathFinder_9_clock),
    .reset(PathFinder_9_reset),
    .io_Stationary_matrix_0_0(PathFinder_9_io_Stationary_matrix_0_0),
    .io_Stationary_matrix_0_1(PathFinder_9_io_Stationary_matrix_0_1),
    .io_Stationary_matrix_0_2(PathFinder_9_io_Stationary_matrix_0_2),
    .io_Stationary_matrix_0_3(PathFinder_9_io_Stationary_matrix_0_3),
    .io_Stationary_matrix_0_4(PathFinder_9_io_Stationary_matrix_0_4),
    .io_Stationary_matrix_0_5(PathFinder_9_io_Stationary_matrix_0_5),
    .io_Stationary_matrix_0_6(PathFinder_9_io_Stationary_matrix_0_6),
    .io_Stationary_matrix_0_7(PathFinder_9_io_Stationary_matrix_0_7),
    .io_Stationary_matrix_1_0(PathFinder_9_io_Stationary_matrix_1_0),
    .io_Stationary_matrix_1_1(PathFinder_9_io_Stationary_matrix_1_1),
    .io_Stationary_matrix_1_2(PathFinder_9_io_Stationary_matrix_1_2),
    .io_Stationary_matrix_1_3(PathFinder_9_io_Stationary_matrix_1_3),
    .io_Stationary_matrix_1_4(PathFinder_9_io_Stationary_matrix_1_4),
    .io_Stationary_matrix_1_5(PathFinder_9_io_Stationary_matrix_1_5),
    .io_Stationary_matrix_1_6(PathFinder_9_io_Stationary_matrix_1_6),
    .io_Stationary_matrix_1_7(PathFinder_9_io_Stationary_matrix_1_7),
    .io_Stationary_matrix_2_0(PathFinder_9_io_Stationary_matrix_2_0),
    .io_Stationary_matrix_2_1(PathFinder_9_io_Stationary_matrix_2_1),
    .io_Stationary_matrix_2_2(PathFinder_9_io_Stationary_matrix_2_2),
    .io_Stationary_matrix_2_3(PathFinder_9_io_Stationary_matrix_2_3),
    .io_Stationary_matrix_2_4(PathFinder_9_io_Stationary_matrix_2_4),
    .io_Stationary_matrix_2_5(PathFinder_9_io_Stationary_matrix_2_5),
    .io_Stationary_matrix_2_6(PathFinder_9_io_Stationary_matrix_2_6),
    .io_Stationary_matrix_2_7(PathFinder_9_io_Stationary_matrix_2_7),
    .io_Stationary_matrix_3_0(PathFinder_9_io_Stationary_matrix_3_0),
    .io_Stationary_matrix_3_1(PathFinder_9_io_Stationary_matrix_3_1),
    .io_Stationary_matrix_3_2(PathFinder_9_io_Stationary_matrix_3_2),
    .io_Stationary_matrix_3_3(PathFinder_9_io_Stationary_matrix_3_3),
    .io_Stationary_matrix_3_4(PathFinder_9_io_Stationary_matrix_3_4),
    .io_Stationary_matrix_3_5(PathFinder_9_io_Stationary_matrix_3_5),
    .io_Stationary_matrix_3_6(PathFinder_9_io_Stationary_matrix_3_6),
    .io_Stationary_matrix_3_7(PathFinder_9_io_Stationary_matrix_3_7),
    .io_Stationary_matrix_4_0(PathFinder_9_io_Stationary_matrix_4_0),
    .io_Stationary_matrix_4_1(PathFinder_9_io_Stationary_matrix_4_1),
    .io_Stationary_matrix_4_2(PathFinder_9_io_Stationary_matrix_4_2),
    .io_Stationary_matrix_4_3(PathFinder_9_io_Stationary_matrix_4_3),
    .io_Stationary_matrix_4_4(PathFinder_9_io_Stationary_matrix_4_4),
    .io_Stationary_matrix_4_5(PathFinder_9_io_Stationary_matrix_4_5),
    .io_Stationary_matrix_4_6(PathFinder_9_io_Stationary_matrix_4_6),
    .io_Stationary_matrix_4_7(PathFinder_9_io_Stationary_matrix_4_7),
    .io_Stationary_matrix_5_0(PathFinder_9_io_Stationary_matrix_5_0),
    .io_Stationary_matrix_5_1(PathFinder_9_io_Stationary_matrix_5_1),
    .io_Stationary_matrix_5_2(PathFinder_9_io_Stationary_matrix_5_2),
    .io_Stationary_matrix_5_3(PathFinder_9_io_Stationary_matrix_5_3),
    .io_Stationary_matrix_5_4(PathFinder_9_io_Stationary_matrix_5_4),
    .io_Stationary_matrix_5_5(PathFinder_9_io_Stationary_matrix_5_5),
    .io_Stationary_matrix_5_6(PathFinder_9_io_Stationary_matrix_5_6),
    .io_Stationary_matrix_5_7(PathFinder_9_io_Stationary_matrix_5_7),
    .io_Stationary_matrix_6_0(PathFinder_9_io_Stationary_matrix_6_0),
    .io_Stationary_matrix_6_1(PathFinder_9_io_Stationary_matrix_6_1),
    .io_Stationary_matrix_6_2(PathFinder_9_io_Stationary_matrix_6_2),
    .io_Stationary_matrix_6_3(PathFinder_9_io_Stationary_matrix_6_3),
    .io_Stationary_matrix_6_4(PathFinder_9_io_Stationary_matrix_6_4),
    .io_Stationary_matrix_6_5(PathFinder_9_io_Stationary_matrix_6_5),
    .io_Stationary_matrix_6_6(PathFinder_9_io_Stationary_matrix_6_6),
    .io_Stationary_matrix_6_7(PathFinder_9_io_Stationary_matrix_6_7),
    .io_Stationary_matrix_7_0(PathFinder_9_io_Stationary_matrix_7_0),
    .io_Stationary_matrix_7_1(PathFinder_9_io_Stationary_matrix_7_1),
    .io_Stationary_matrix_7_2(PathFinder_9_io_Stationary_matrix_7_2),
    .io_Stationary_matrix_7_3(PathFinder_9_io_Stationary_matrix_7_3),
    .io_Stationary_matrix_7_4(PathFinder_9_io_Stationary_matrix_7_4),
    .io_Stationary_matrix_7_5(PathFinder_9_io_Stationary_matrix_7_5),
    .io_Stationary_matrix_7_6(PathFinder_9_io_Stationary_matrix_7_6),
    .io_Stationary_matrix_7_7(PathFinder_9_io_Stationary_matrix_7_7),
    .io_Streaming_matrix_0(PathFinder_9_io_Streaming_matrix_0),
    .io_Streaming_matrix_1(PathFinder_9_io_Streaming_matrix_1),
    .io_Streaming_matrix_2(PathFinder_9_io_Streaming_matrix_2),
    .io_Streaming_matrix_3(PathFinder_9_io_Streaming_matrix_3),
    .io_Streaming_matrix_4(PathFinder_9_io_Streaming_matrix_4),
    .io_Streaming_matrix_5(PathFinder_9_io_Streaming_matrix_5),
    .io_Streaming_matrix_6(PathFinder_9_io_Streaming_matrix_6),
    .io_Streaming_matrix_7(PathFinder_9_io_Streaming_matrix_7),
    .io_i_mux_bus_0(PathFinder_9_io_i_mux_bus_0),
    .io_i_mux_bus_1(PathFinder_9_io_i_mux_bus_1),
    .io_i_mux_bus_2(PathFinder_9_io_i_mux_bus_2),
    .io_i_mux_bus_3(PathFinder_9_io_i_mux_bus_3),
    .io_Source_0(PathFinder_9_io_Source_0),
    .io_Source_1(PathFinder_9_io_Source_1),
    .io_Source_2(PathFinder_9_io_Source_2),
    .io_Source_3(PathFinder_9_io_Source_3),
    .io_destination_0(PathFinder_9_io_destination_0),
    .io_destination_1(PathFinder_9_io_destination_1),
    .io_destination_2(PathFinder_9_io_destination_2),
    .io_destination_3(PathFinder_9_io_destination_3),
    .io_PF_Valid(PathFinder_9_io_PF_Valid),
    .io_NoDPE(PathFinder_9_io_NoDPE),
    .io_DataValid(PathFinder_9_io_DataValid)
  );
  PathFinder PathFinder_10 ( // @[FlexDPU.scala 77:41]
    .clock(PathFinder_10_clock),
    .reset(PathFinder_10_reset),
    .io_Stationary_matrix_0_0(PathFinder_10_io_Stationary_matrix_0_0),
    .io_Stationary_matrix_0_1(PathFinder_10_io_Stationary_matrix_0_1),
    .io_Stationary_matrix_0_2(PathFinder_10_io_Stationary_matrix_0_2),
    .io_Stationary_matrix_0_3(PathFinder_10_io_Stationary_matrix_0_3),
    .io_Stationary_matrix_0_4(PathFinder_10_io_Stationary_matrix_0_4),
    .io_Stationary_matrix_0_5(PathFinder_10_io_Stationary_matrix_0_5),
    .io_Stationary_matrix_0_6(PathFinder_10_io_Stationary_matrix_0_6),
    .io_Stationary_matrix_0_7(PathFinder_10_io_Stationary_matrix_0_7),
    .io_Stationary_matrix_1_0(PathFinder_10_io_Stationary_matrix_1_0),
    .io_Stationary_matrix_1_1(PathFinder_10_io_Stationary_matrix_1_1),
    .io_Stationary_matrix_1_2(PathFinder_10_io_Stationary_matrix_1_2),
    .io_Stationary_matrix_1_3(PathFinder_10_io_Stationary_matrix_1_3),
    .io_Stationary_matrix_1_4(PathFinder_10_io_Stationary_matrix_1_4),
    .io_Stationary_matrix_1_5(PathFinder_10_io_Stationary_matrix_1_5),
    .io_Stationary_matrix_1_6(PathFinder_10_io_Stationary_matrix_1_6),
    .io_Stationary_matrix_1_7(PathFinder_10_io_Stationary_matrix_1_7),
    .io_Stationary_matrix_2_0(PathFinder_10_io_Stationary_matrix_2_0),
    .io_Stationary_matrix_2_1(PathFinder_10_io_Stationary_matrix_2_1),
    .io_Stationary_matrix_2_2(PathFinder_10_io_Stationary_matrix_2_2),
    .io_Stationary_matrix_2_3(PathFinder_10_io_Stationary_matrix_2_3),
    .io_Stationary_matrix_2_4(PathFinder_10_io_Stationary_matrix_2_4),
    .io_Stationary_matrix_2_5(PathFinder_10_io_Stationary_matrix_2_5),
    .io_Stationary_matrix_2_6(PathFinder_10_io_Stationary_matrix_2_6),
    .io_Stationary_matrix_2_7(PathFinder_10_io_Stationary_matrix_2_7),
    .io_Stationary_matrix_3_0(PathFinder_10_io_Stationary_matrix_3_0),
    .io_Stationary_matrix_3_1(PathFinder_10_io_Stationary_matrix_3_1),
    .io_Stationary_matrix_3_2(PathFinder_10_io_Stationary_matrix_3_2),
    .io_Stationary_matrix_3_3(PathFinder_10_io_Stationary_matrix_3_3),
    .io_Stationary_matrix_3_4(PathFinder_10_io_Stationary_matrix_3_4),
    .io_Stationary_matrix_3_5(PathFinder_10_io_Stationary_matrix_3_5),
    .io_Stationary_matrix_3_6(PathFinder_10_io_Stationary_matrix_3_6),
    .io_Stationary_matrix_3_7(PathFinder_10_io_Stationary_matrix_3_7),
    .io_Stationary_matrix_4_0(PathFinder_10_io_Stationary_matrix_4_0),
    .io_Stationary_matrix_4_1(PathFinder_10_io_Stationary_matrix_4_1),
    .io_Stationary_matrix_4_2(PathFinder_10_io_Stationary_matrix_4_2),
    .io_Stationary_matrix_4_3(PathFinder_10_io_Stationary_matrix_4_3),
    .io_Stationary_matrix_4_4(PathFinder_10_io_Stationary_matrix_4_4),
    .io_Stationary_matrix_4_5(PathFinder_10_io_Stationary_matrix_4_5),
    .io_Stationary_matrix_4_6(PathFinder_10_io_Stationary_matrix_4_6),
    .io_Stationary_matrix_4_7(PathFinder_10_io_Stationary_matrix_4_7),
    .io_Stationary_matrix_5_0(PathFinder_10_io_Stationary_matrix_5_0),
    .io_Stationary_matrix_5_1(PathFinder_10_io_Stationary_matrix_5_1),
    .io_Stationary_matrix_5_2(PathFinder_10_io_Stationary_matrix_5_2),
    .io_Stationary_matrix_5_3(PathFinder_10_io_Stationary_matrix_5_3),
    .io_Stationary_matrix_5_4(PathFinder_10_io_Stationary_matrix_5_4),
    .io_Stationary_matrix_5_5(PathFinder_10_io_Stationary_matrix_5_5),
    .io_Stationary_matrix_5_6(PathFinder_10_io_Stationary_matrix_5_6),
    .io_Stationary_matrix_5_7(PathFinder_10_io_Stationary_matrix_5_7),
    .io_Stationary_matrix_6_0(PathFinder_10_io_Stationary_matrix_6_0),
    .io_Stationary_matrix_6_1(PathFinder_10_io_Stationary_matrix_6_1),
    .io_Stationary_matrix_6_2(PathFinder_10_io_Stationary_matrix_6_2),
    .io_Stationary_matrix_6_3(PathFinder_10_io_Stationary_matrix_6_3),
    .io_Stationary_matrix_6_4(PathFinder_10_io_Stationary_matrix_6_4),
    .io_Stationary_matrix_6_5(PathFinder_10_io_Stationary_matrix_6_5),
    .io_Stationary_matrix_6_6(PathFinder_10_io_Stationary_matrix_6_6),
    .io_Stationary_matrix_6_7(PathFinder_10_io_Stationary_matrix_6_7),
    .io_Stationary_matrix_7_0(PathFinder_10_io_Stationary_matrix_7_0),
    .io_Stationary_matrix_7_1(PathFinder_10_io_Stationary_matrix_7_1),
    .io_Stationary_matrix_7_2(PathFinder_10_io_Stationary_matrix_7_2),
    .io_Stationary_matrix_7_3(PathFinder_10_io_Stationary_matrix_7_3),
    .io_Stationary_matrix_7_4(PathFinder_10_io_Stationary_matrix_7_4),
    .io_Stationary_matrix_7_5(PathFinder_10_io_Stationary_matrix_7_5),
    .io_Stationary_matrix_7_6(PathFinder_10_io_Stationary_matrix_7_6),
    .io_Stationary_matrix_7_7(PathFinder_10_io_Stationary_matrix_7_7),
    .io_Streaming_matrix_0(PathFinder_10_io_Streaming_matrix_0),
    .io_Streaming_matrix_1(PathFinder_10_io_Streaming_matrix_1),
    .io_Streaming_matrix_2(PathFinder_10_io_Streaming_matrix_2),
    .io_Streaming_matrix_3(PathFinder_10_io_Streaming_matrix_3),
    .io_Streaming_matrix_4(PathFinder_10_io_Streaming_matrix_4),
    .io_Streaming_matrix_5(PathFinder_10_io_Streaming_matrix_5),
    .io_Streaming_matrix_6(PathFinder_10_io_Streaming_matrix_6),
    .io_Streaming_matrix_7(PathFinder_10_io_Streaming_matrix_7),
    .io_i_mux_bus_0(PathFinder_10_io_i_mux_bus_0),
    .io_i_mux_bus_1(PathFinder_10_io_i_mux_bus_1),
    .io_i_mux_bus_2(PathFinder_10_io_i_mux_bus_2),
    .io_i_mux_bus_3(PathFinder_10_io_i_mux_bus_3),
    .io_Source_0(PathFinder_10_io_Source_0),
    .io_Source_1(PathFinder_10_io_Source_1),
    .io_Source_2(PathFinder_10_io_Source_2),
    .io_Source_3(PathFinder_10_io_Source_3),
    .io_destination_0(PathFinder_10_io_destination_0),
    .io_destination_1(PathFinder_10_io_destination_1),
    .io_destination_2(PathFinder_10_io_destination_2),
    .io_destination_3(PathFinder_10_io_destination_3),
    .io_PF_Valid(PathFinder_10_io_PF_Valid),
    .io_NoDPE(PathFinder_10_io_NoDPE),
    .io_DataValid(PathFinder_10_io_DataValid)
  );
  PathFinder PathFinder_11 ( // @[FlexDPU.scala 77:41]
    .clock(PathFinder_11_clock),
    .reset(PathFinder_11_reset),
    .io_Stationary_matrix_0_0(PathFinder_11_io_Stationary_matrix_0_0),
    .io_Stationary_matrix_0_1(PathFinder_11_io_Stationary_matrix_0_1),
    .io_Stationary_matrix_0_2(PathFinder_11_io_Stationary_matrix_0_2),
    .io_Stationary_matrix_0_3(PathFinder_11_io_Stationary_matrix_0_3),
    .io_Stationary_matrix_0_4(PathFinder_11_io_Stationary_matrix_0_4),
    .io_Stationary_matrix_0_5(PathFinder_11_io_Stationary_matrix_0_5),
    .io_Stationary_matrix_0_6(PathFinder_11_io_Stationary_matrix_0_6),
    .io_Stationary_matrix_0_7(PathFinder_11_io_Stationary_matrix_0_7),
    .io_Stationary_matrix_1_0(PathFinder_11_io_Stationary_matrix_1_0),
    .io_Stationary_matrix_1_1(PathFinder_11_io_Stationary_matrix_1_1),
    .io_Stationary_matrix_1_2(PathFinder_11_io_Stationary_matrix_1_2),
    .io_Stationary_matrix_1_3(PathFinder_11_io_Stationary_matrix_1_3),
    .io_Stationary_matrix_1_4(PathFinder_11_io_Stationary_matrix_1_4),
    .io_Stationary_matrix_1_5(PathFinder_11_io_Stationary_matrix_1_5),
    .io_Stationary_matrix_1_6(PathFinder_11_io_Stationary_matrix_1_6),
    .io_Stationary_matrix_1_7(PathFinder_11_io_Stationary_matrix_1_7),
    .io_Stationary_matrix_2_0(PathFinder_11_io_Stationary_matrix_2_0),
    .io_Stationary_matrix_2_1(PathFinder_11_io_Stationary_matrix_2_1),
    .io_Stationary_matrix_2_2(PathFinder_11_io_Stationary_matrix_2_2),
    .io_Stationary_matrix_2_3(PathFinder_11_io_Stationary_matrix_2_3),
    .io_Stationary_matrix_2_4(PathFinder_11_io_Stationary_matrix_2_4),
    .io_Stationary_matrix_2_5(PathFinder_11_io_Stationary_matrix_2_5),
    .io_Stationary_matrix_2_6(PathFinder_11_io_Stationary_matrix_2_6),
    .io_Stationary_matrix_2_7(PathFinder_11_io_Stationary_matrix_2_7),
    .io_Stationary_matrix_3_0(PathFinder_11_io_Stationary_matrix_3_0),
    .io_Stationary_matrix_3_1(PathFinder_11_io_Stationary_matrix_3_1),
    .io_Stationary_matrix_3_2(PathFinder_11_io_Stationary_matrix_3_2),
    .io_Stationary_matrix_3_3(PathFinder_11_io_Stationary_matrix_3_3),
    .io_Stationary_matrix_3_4(PathFinder_11_io_Stationary_matrix_3_4),
    .io_Stationary_matrix_3_5(PathFinder_11_io_Stationary_matrix_3_5),
    .io_Stationary_matrix_3_6(PathFinder_11_io_Stationary_matrix_3_6),
    .io_Stationary_matrix_3_7(PathFinder_11_io_Stationary_matrix_3_7),
    .io_Stationary_matrix_4_0(PathFinder_11_io_Stationary_matrix_4_0),
    .io_Stationary_matrix_4_1(PathFinder_11_io_Stationary_matrix_4_1),
    .io_Stationary_matrix_4_2(PathFinder_11_io_Stationary_matrix_4_2),
    .io_Stationary_matrix_4_3(PathFinder_11_io_Stationary_matrix_4_3),
    .io_Stationary_matrix_4_4(PathFinder_11_io_Stationary_matrix_4_4),
    .io_Stationary_matrix_4_5(PathFinder_11_io_Stationary_matrix_4_5),
    .io_Stationary_matrix_4_6(PathFinder_11_io_Stationary_matrix_4_6),
    .io_Stationary_matrix_4_7(PathFinder_11_io_Stationary_matrix_4_7),
    .io_Stationary_matrix_5_0(PathFinder_11_io_Stationary_matrix_5_0),
    .io_Stationary_matrix_5_1(PathFinder_11_io_Stationary_matrix_5_1),
    .io_Stationary_matrix_5_2(PathFinder_11_io_Stationary_matrix_5_2),
    .io_Stationary_matrix_5_3(PathFinder_11_io_Stationary_matrix_5_3),
    .io_Stationary_matrix_5_4(PathFinder_11_io_Stationary_matrix_5_4),
    .io_Stationary_matrix_5_5(PathFinder_11_io_Stationary_matrix_5_5),
    .io_Stationary_matrix_5_6(PathFinder_11_io_Stationary_matrix_5_6),
    .io_Stationary_matrix_5_7(PathFinder_11_io_Stationary_matrix_5_7),
    .io_Stationary_matrix_6_0(PathFinder_11_io_Stationary_matrix_6_0),
    .io_Stationary_matrix_6_1(PathFinder_11_io_Stationary_matrix_6_1),
    .io_Stationary_matrix_6_2(PathFinder_11_io_Stationary_matrix_6_2),
    .io_Stationary_matrix_6_3(PathFinder_11_io_Stationary_matrix_6_3),
    .io_Stationary_matrix_6_4(PathFinder_11_io_Stationary_matrix_6_4),
    .io_Stationary_matrix_6_5(PathFinder_11_io_Stationary_matrix_6_5),
    .io_Stationary_matrix_6_6(PathFinder_11_io_Stationary_matrix_6_6),
    .io_Stationary_matrix_6_7(PathFinder_11_io_Stationary_matrix_6_7),
    .io_Stationary_matrix_7_0(PathFinder_11_io_Stationary_matrix_7_0),
    .io_Stationary_matrix_7_1(PathFinder_11_io_Stationary_matrix_7_1),
    .io_Stationary_matrix_7_2(PathFinder_11_io_Stationary_matrix_7_2),
    .io_Stationary_matrix_7_3(PathFinder_11_io_Stationary_matrix_7_3),
    .io_Stationary_matrix_7_4(PathFinder_11_io_Stationary_matrix_7_4),
    .io_Stationary_matrix_7_5(PathFinder_11_io_Stationary_matrix_7_5),
    .io_Stationary_matrix_7_6(PathFinder_11_io_Stationary_matrix_7_6),
    .io_Stationary_matrix_7_7(PathFinder_11_io_Stationary_matrix_7_7),
    .io_Streaming_matrix_0(PathFinder_11_io_Streaming_matrix_0),
    .io_Streaming_matrix_1(PathFinder_11_io_Streaming_matrix_1),
    .io_Streaming_matrix_2(PathFinder_11_io_Streaming_matrix_2),
    .io_Streaming_matrix_3(PathFinder_11_io_Streaming_matrix_3),
    .io_Streaming_matrix_4(PathFinder_11_io_Streaming_matrix_4),
    .io_Streaming_matrix_5(PathFinder_11_io_Streaming_matrix_5),
    .io_Streaming_matrix_6(PathFinder_11_io_Streaming_matrix_6),
    .io_Streaming_matrix_7(PathFinder_11_io_Streaming_matrix_7),
    .io_i_mux_bus_0(PathFinder_11_io_i_mux_bus_0),
    .io_i_mux_bus_1(PathFinder_11_io_i_mux_bus_1),
    .io_i_mux_bus_2(PathFinder_11_io_i_mux_bus_2),
    .io_i_mux_bus_3(PathFinder_11_io_i_mux_bus_3),
    .io_Source_0(PathFinder_11_io_Source_0),
    .io_Source_1(PathFinder_11_io_Source_1),
    .io_Source_2(PathFinder_11_io_Source_2),
    .io_Source_3(PathFinder_11_io_Source_3),
    .io_destination_0(PathFinder_11_io_destination_0),
    .io_destination_1(PathFinder_11_io_destination_1),
    .io_destination_2(PathFinder_11_io_destination_2),
    .io_destination_3(PathFinder_11_io_destination_3),
    .io_PF_Valid(PathFinder_11_io_PF_Valid),
    .io_NoDPE(PathFinder_11_io_NoDPE),
    .io_DataValid(PathFinder_11_io_DataValid)
  );
  PathFinder PathFinder_12 ( // @[FlexDPU.scala 77:41]
    .clock(PathFinder_12_clock),
    .reset(PathFinder_12_reset),
    .io_Stationary_matrix_0_0(PathFinder_12_io_Stationary_matrix_0_0),
    .io_Stationary_matrix_0_1(PathFinder_12_io_Stationary_matrix_0_1),
    .io_Stationary_matrix_0_2(PathFinder_12_io_Stationary_matrix_0_2),
    .io_Stationary_matrix_0_3(PathFinder_12_io_Stationary_matrix_0_3),
    .io_Stationary_matrix_0_4(PathFinder_12_io_Stationary_matrix_0_4),
    .io_Stationary_matrix_0_5(PathFinder_12_io_Stationary_matrix_0_5),
    .io_Stationary_matrix_0_6(PathFinder_12_io_Stationary_matrix_0_6),
    .io_Stationary_matrix_0_7(PathFinder_12_io_Stationary_matrix_0_7),
    .io_Stationary_matrix_1_0(PathFinder_12_io_Stationary_matrix_1_0),
    .io_Stationary_matrix_1_1(PathFinder_12_io_Stationary_matrix_1_1),
    .io_Stationary_matrix_1_2(PathFinder_12_io_Stationary_matrix_1_2),
    .io_Stationary_matrix_1_3(PathFinder_12_io_Stationary_matrix_1_3),
    .io_Stationary_matrix_1_4(PathFinder_12_io_Stationary_matrix_1_4),
    .io_Stationary_matrix_1_5(PathFinder_12_io_Stationary_matrix_1_5),
    .io_Stationary_matrix_1_6(PathFinder_12_io_Stationary_matrix_1_6),
    .io_Stationary_matrix_1_7(PathFinder_12_io_Stationary_matrix_1_7),
    .io_Stationary_matrix_2_0(PathFinder_12_io_Stationary_matrix_2_0),
    .io_Stationary_matrix_2_1(PathFinder_12_io_Stationary_matrix_2_1),
    .io_Stationary_matrix_2_2(PathFinder_12_io_Stationary_matrix_2_2),
    .io_Stationary_matrix_2_3(PathFinder_12_io_Stationary_matrix_2_3),
    .io_Stationary_matrix_2_4(PathFinder_12_io_Stationary_matrix_2_4),
    .io_Stationary_matrix_2_5(PathFinder_12_io_Stationary_matrix_2_5),
    .io_Stationary_matrix_2_6(PathFinder_12_io_Stationary_matrix_2_6),
    .io_Stationary_matrix_2_7(PathFinder_12_io_Stationary_matrix_2_7),
    .io_Stationary_matrix_3_0(PathFinder_12_io_Stationary_matrix_3_0),
    .io_Stationary_matrix_3_1(PathFinder_12_io_Stationary_matrix_3_1),
    .io_Stationary_matrix_3_2(PathFinder_12_io_Stationary_matrix_3_2),
    .io_Stationary_matrix_3_3(PathFinder_12_io_Stationary_matrix_3_3),
    .io_Stationary_matrix_3_4(PathFinder_12_io_Stationary_matrix_3_4),
    .io_Stationary_matrix_3_5(PathFinder_12_io_Stationary_matrix_3_5),
    .io_Stationary_matrix_3_6(PathFinder_12_io_Stationary_matrix_3_6),
    .io_Stationary_matrix_3_7(PathFinder_12_io_Stationary_matrix_3_7),
    .io_Stationary_matrix_4_0(PathFinder_12_io_Stationary_matrix_4_0),
    .io_Stationary_matrix_4_1(PathFinder_12_io_Stationary_matrix_4_1),
    .io_Stationary_matrix_4_2(PathFinder_12_io_Stationary_matrix_4_2),
    .io_Stationary_matrix_4_3(PathFinder_12_io_Stationary_matrix_4_3),
    .io_Stationary_matrix_4_4(PathFinder_12_io_Stationary_matrix_4_4),
    .io_Stationary_matrix_4_5(PathFinder_12_io_Stationary_matrix_4_5),
    .io_Stationary_matrix_4_6(PathFinder_12_io_Stationary_matrix_4_6),
    .io_Stationary_matrix_4_7(PathFinder_12_io_Stationary_matrix_4_7),
    .io_Stationary_matrix_5_0(PathFinder_12_io_Stationary_matrix_5_0),
    .io_Stationary_matrix_5_1(PathFinder_12_io_Stationary_matrix_5_1),
    .io_Stationary_matrix_5_2(PathFinder_12_io_Stationary_matrix_5_2),
    .io_Stationary_matrix_5_3(PathFinder_12_io_Stationary_matrix_5_3),
    .io_Stationary_matrix_5_4(PathFinder_12_io_Stationary_matrix_5_4),
    .io_Stationary_matrix_5_5(PathFinder_12_io_Stationary_matrix_5_5),
    .io_Stationary_matrix_5_6(PathFinder_12_io_Stationary_matrix_5_6),
    .io_Stationary_matrix_5_7(PathFinder_12_io_Stationary_matrix_5_7),
    .io_Stationary_matrix_6_0(PathFinder_12_io_Stationary_matrix_6_0),
    .io_Stationary_matrix_6_1(PathFinder_12_io_Stationary_matrix_6_1),
    .io_Stationary_matrix_6_2(PathFinder_12_io_Stationary_matrix_6_2),
    .io_Stationary_matrix_6_3(PathFinder_12_io_Stationary_matrix_6_3),
    .io_Stationary_matrix_6_4(PathFinder_12_io_Stationary_matrix_6_4),
    .io_Stationary_matrix_6_5(PathFinder_12_io_Stationary_matrix_6_5),
    .io_Stationary_matrix_6_6(PathFinder_12_io_Stationary_matrix_6_6),
    .io_Stationary_matrix_6_7(PathFinder_12_io_Stationary_matrix_6_7),
    .io_Stationary_matrix_7_0(PathFinder_12_io_Stationary_matrix_7_0),
    .io_Stationary_matrix_7_1(PathFinder_12_io_Stationary_matrix_7_1),
    .io_Stationary_matrix_7_2(PathFinder_12_io_Stationary_matrix_7_2),
    .io_Stationary_matrix_7_3(PathFinder_12_io_Stationary_matrix_7_3),
    .io_Stationary_matrix_7_4(PathFinder_12_io_Stationary_matrix_7_4),
    .io_Stationary_matrix_7_5(PathFinder_12_io_Stationary_matrix_7_5),
    .io_Stationary_matrix_7_6(PathFinder_12_io_Stationary_matrix_7_6),
    .io_Stationary_matrix_7_7(PathFinder_12_io_Stationary_matrix_7_7),
    .io_Streaming_matrix_0(PathFinder_12_io_Streaming_matrix_0),
    .io_Streaming_matrix_1(PathFinder_12_io_Streaming_matrix_1),
    .io_Streaming_matrix_2(PathFinder_12_io_Streaming_matrix_2),
    .io_Streaming_matrix_3(PathFinder_12_io_Streaming_matrix_3),
    .io_Streaming_matrix_4(PathFinder_12_io_Streaming_matrix_4),
    .io_Streaming_matrix_5(PathFinder_12_io_Streaming_matrix_5),
    .io_Streaming_matrix_6(PathFinder_12_io_Streaming_matrix_6),
    .io_Streaming_matrix_7(PathFinder_12_io_Streaming_matrix_7),
    .io_i_mux_bus_0(PathFinder_12_io_i_mux_bus_0),
    .io_i_mux_bus_1(PathFinder_12_io_i_mux_bus_1),
    .io_i_mux_bus_2(PathFinder_12_io_i_mux_bus_2),
    .io_i_mux_bus_3(PathFinder_12_io_i_mux_bus_3),
    .io_Source_0(PathFinder_12_io_Source_0),
    .io_Source_1(PathFinder_12_io_Source_1),
    .io_Source_2(PathFinder_12_io_Source_2),
    .io_Source_3(PathFinder_12_io_Source_3),
    .io_destination_0(PathFinder_12_io_destination_0),
    .io_destination_1(PathFinder_12_io_destination_1),
    .io_destination_2(PathFinder_12_io_destination_2),
    .io_destination_3(PathFinder_12_io_destination_3),
    .io_PF_Valid(PathFinder_12_io_PF_Valid),
    .io_NoDPE(PathFinder_12_io_NoDPE),
    .io_DataValid(PathFinder_12_io_DataValid)
  );
  PathFinder PathFinder_13 ( // @[FlexDPU.scala 77:41]
    .clock(PathFinder_13_clock),
    .reset(PathFinder_13_reset),
    .io_Stationary_matrix_0_0(PathFinder_13_io_Stationary_matrix_0_0),
    .io_Stationary_matrix_0_1(PathFinder_13_io_Stationary_matrix_0_1),
    .io_Stationary_matrix_0_2(PathFinder_13_io_Stationary_matrix_0_2),
    .io_Stationary_matrix_0_3(PathFinder_13_io_Stationary_matrix_0_3),
    .io_Stationary_matrix_0_4(PathFinder_13_io_Stationary_matrix_0_4),
    .io_Stationary_matrix_0_5(PathFinder_13_io_Stationary_matrix_0_5),
    .io_Stationary_matrix_0_6(PathFinder_13_io_Stationary_matrix_0_6),
    .io_Stationary_matrix_0_7(PathFinder_13_io_Stationary_matrix_0_7),
    .io_Stationary_matrix_1_0(PathFinder_13_io_Stationary_matrix_1_0),
    .io_Stationary_matrix_1_1(PathFinder_13_io_Stationary_matrix_1_1),
    .io_Stationary_matrix_1_2(PathFinder_13_io_Stationary_matrix_1_2),
    .io_Stationary_matrix_1_3(PathFinder_13_io_Stationary_matrix_1_3),
    .io_Stationary_matrix_1_4(PathFinder_13_io_Stationary_matrix_1_4),
    .io_Stationary_matrix_1_5(PathFinder_13_io_Stationary_matrix_1_5),
    .io_Stationary_matrix_1_6(PathFinder_13_io_Stationary_matrix_1_6),
    .io_Stationary_matrix_1_7(PathFinder_13_io_Stationary_matrix_1_7),
    .io_Stationary_matrix_2_0(PathFinder_13_io_Stationary_matrix_2_0),
    .io_Stationary_matrix_2_1(PathFinder_13_io_Stationary_matrix_2_1),
    .io_Stationary_matrix_2_2(PathFinder_13_io_Stationary_matrix_2_2),
    .io_Stationary_matrix_2_3(PathFinder_13_io_Stationary_matrix_2_3),
    .io_Stationary_matrix_2_4(PathFinder_13_io_Stationary_matrix_2_4),
    .io_Stationary_matrix_2_5(PathFinder_13_io_Stationary_matrix_2_5),
    .io_Stationary_matrix_2_6(PathFinder_13_io_Stationary_matrix_2_6),
    .io_Stationary_matrix_2_7(PathFinder_13_io_Stationary_matrix_2_7),
    .io_Stationary_matrix_3_0(PathFinder_13_io_Stationary_matrix_3_0),
    .io_Stationary_matrix_3_1(PathFinder_13_io_Stationary_matrix_3_1),
    .io_Stationary_matrix_3_2(PathFinder_13_io_Stationary_matrix_3_2),
    .io_Stationary_matrix_3_3(PathFinder_13_io_Stationary_matrix_3_3),
    .io_Stationary_matrix_3_4(PathFinder_13_io_Stationary_matrix_3_4),
    .io_Stationary_matrix_3_5(PathFinder_13_io_Stationary_matrix_3_5),
    .io_Stationary_matrix_3_6(PathFinder_13_io_Stationary_matrix_3_6),
    .io_Stationary_matrix_3_7(PathFinder_13_io_Stationary_matrix_3_7),
    .io_Stationary_matrix_4_0(PathFinder_13_io_Stationary_matrix_4_0),
    .io_Stationary_matrix_4_1(PathFinder_13_io_Stationary_matrix_4_1),
    .io_Stationary_matrix_4_2(PathFinder_13_io_Stationary_matrix_4_2),
    .io_Stationary_matrix_4_3(PathFinder_13_io_Stationary_matrix_4_3),
    .io_Stationary_matrix_4_4(PathFinder_13_io_Stationary_matrix_4_4),
    .io_Stationary_matrix_4_5(PathFinder_13_io_Stationary_matrix_4_5),
    .io_Stationary_matrix_4_6(PathFinder_13_io_Stationary_matrix_4_6),
    .io_Stationary_matrix_4_7(PathFinder_13_io_Stationary_matrix_4_7),
    .io_Stationary_matrix_5_0(PathFinder_13_io_Stationary_matrix_5_0),
    .io_Stationary_matrix_5_1(PathFinder_13_io_Stationary_matrix_5_1),
    .io_Stationary_matrix_5_2(PathFinder_13_io_Stationary_matrix_5_2),
    .io_Stationary_matrix_5_3(PathFinder_13_io_Stationary_matrix_5_3),
    .io_Stationary_matrix_5_4(PathFinder_13_io_Stationary_matrix_5_4),
    .io_Stationary_matrix_5_5(PathFinder_13_io_Stationary_matrix_5_5),
    .io_Stationary_matrix_5_6(PathFinder_13_io_Stationary_matrix_5_6),
    .io_Stationary_matrix_5_7(PathFinder_13_io_Stationary_matrix_5_7),
    .io_Stationary_matrix_6_0(PathFinder_13_io_Stationary_matrix_6_0),
    .io_Stationary_matrix_6_1(PathFinder_13_io_Stationary_matrix_6_1),
    .io_Stationary_matrix_6_2(PathFinder_13_io_Stationary_matrix_6_2),
    .io_Stationary_matrix_6_3(PathFinder_13_io_Stationary_matrix_6_3),
    .io_Stationary_matrix_6_4(PathFinder_13_io_Stationary_matrix_6_4),
    .io_Stationary_matrix_6_5(PathFinder_13_io_Stationary_matrix_6_5),
    .io_Stationary_matrix_6_6(PathFinder_13_io_Stationary_matrix_6_6),
    .io_Stationary_matrix_6_7(PathFinder_13_io_Stationary_matrix_6_7),
    .io_Stationary_matrix_7_0(PathFinder_13_io_Stationary_matrix_7_0),
    .io_Stationary_matrix_7_1(PathFinder_13_io_Stationary_matrix_7_1),
    .io_Stationary_matrix_7_2(PathFinder_13_io_Stationary_matrix_7_2),
    .io_Stationary_matrix_7_3(PathFinder_13_io_Stationary_matrix_7_3),
    .io_Stationary_matrix_7_4(PathFinder_13_io_Stationary_matrix_7_4),
    .io_Stationary_matrix_7_5(PathFinder_13_io_Stationary_matrix_7_5),
    .io_Stationary_matrix_7_6(PathFinder_13_io_Stationary_matrix_7_6),
    .io_Stationary_matrix_7_7(PathFinder_13_io_Stationary_matrix_7_7),
    .io_Streaming_matrix_0(PathFinder_13_io_Streaming_matrix_0),
    .io_Streaming_matrix_1(PathFinder_13_io_Streaming_matrix_1),
    .io_Streaming_matrix_2(PathFinder_13_io_Streaming_matrix_2),
    .io_Streaming_matrix_3(PathFinder_13_io_Streaming_matrix_3),
    .io_Streaming_matrix_4(PathFinder_13_io_Streaming_matrix_4),
    .io_Streaming_matrix_5(PathFinder_13_io_Streaming_matrix_5),
    .io_Streaming_matrix_6(PathFinder_13_io_Streaming_matrix_6),
    .io_Streaming_matrix_7(PathFinder_13_io_Streaming_matrix_7),
    .io_i_mux_bus_0(PathFinder_13_io_i_mux_bus_0),
    .io_i_mux_bus_1(PathFinder_13_io_i_mux_bus_1),
    .io_i_mux_bus_2(PathFinder_13_io_i_mux_bus_2),
    .io_i_mux_bus_3(PathFinder_13_io_i_mux_bus_3),
    .io_Source_0(PathFinder_13_io_Source_0),
    .io_Source_1(PathFinder_13_io_Source_1),
    .io_Source_2(PathFinder_13_io_Source_2),
    .io_Source_3(PathFinder_13_io_Source_3),
    .io_destination_0(PathFinder_13_io_destination_0),
    .io_destination_1(PathFinder_13_io_destination_1),
    .io_destination_2(PathFinder_13_io_destination_2),
    .io_destination_3(PathFinder_13_io_destination_3),
    .io_PF_Valid(PathFinder_13_io_PF_Valid),
    .io_NoDPE(PathFinder_13_io_NoDPE),
    .io_DataValid(PathFinder_13_io_DataValid)
  );
  PathFinder PathFinder_14 ( // @[FlexDPU.scala 77:41]
    .clock(PathFinder_14_clock),
    .reset(PathFinder_14_reset),
    .io_Stationary_matrix_0_0(PathFinder_14_io_Stationary_matrix_0_0),
    .io_Stationary_matrix_0_1(PathFinder_14_io_Stationary_matrix_0_1),
    .io_Stationary_matrix_0_2(PathFinder_14_io_Stationary_matrix_0_2),
    .io_Stationary_matrix_0_3(PathFinder_14_io_Stationary_matrix_0_3),
    .io_Stationary_matrix_0_4(PathFinder_14_io_Stationary_matrix_0_4),
    .io_Stationary_matrix_0_5(PathFinder_14_io_Stationary_matrix_0_5),
    .io_Stationary_matrix_0_6(PathFinder_14_io_Stationary_matrix_0_6),
    .io_Stationary_matrix_0_7(PathFinder_14_io_Stationary_matrix_0_7),
    .io_Stationary_matrix_1_0(PathFinder_14_io_Stationary_matrix_1_0),
    .io_Stationary_matrix_1_1(PathFinder_14_io_Stationary_matrix_1_1),
    .io_Stationary_matrix_1_2(PathFinder_14_io_Stationary_matrix_1_2),
    .io_Stationary_matrix_1_3(PathFinder_14_io_Stationary_matrix_1_3),
    .io_Stationary_matrix_1_4(PathFinder_14_io_Stationary_matrix_1_4),
    .io_Stationary_matrix_1_5(PathFinder_14_io_Stationary_matrix_1_5),
    .io_Stationary_matrix_1_6(PathFinder_14_io_Stationary_matrix_1_6),
    .io_Stationary_matrix_1_7(PathFinder_14_io_Stationary_matrix_1_7),
    .io_Stationary_matrix_2_0(PathFinder_14_io_Stationary_matrix_2_0),
    .io_Stationary_matrix_2_1(PathFinder_14_io_Stationary_matrix_2_1),
    .io_Stationary_matrix_2_2(PathFinder_14_io_Stationary_matrix_2_2),
    .io_Stationary_matrix_2_3(PathFinder_14_io_Stationary_matrix_2_3),
    .io_Stationary_matrix_2_4(PathFinder_14_io_Stationary_matrix_2_4),
    .io_Stationary_matrix_2_5(PathFinder_14_io_Stationary_matrix_2_5),
    .io_Stationary_matrix_2_6(PathFinder_14_io_Stationary_matrix_2_6),
    .io_Stationary_matrix_2_7(PathFinder_14_io_Stationary_matrix_2_7),
    .io_Stationary_matrix_3_0(PathFinder_14_io_Stationary_matrix_3_0),
    .io_Stationary_matrix_3_1(PathFinder_14_io_Stationary_matrix_3_1),
    .io_Stationary_matrix_3_2(PathFinder_14_io_Stationary_matrix_3_2),
    .io_Stationary_matrix_3_3(PathFinder_14_io_Stationary_matrix_3_3),
    .io_Stationary_matrix_3_4(PathFinder_14_io_Stationary_matrix_3_4),
    .io_Stationary_matrix_3_5(PathFinder_14_io_Stationary_matrix_3_5),
    .io_Stationary_matrix_3_6(PathFinder_14_io_Stationary_matrix_3_6),
    .io_Stationary_matrix_3_7(PathFinder_14_io_Stationary_matrix_3_7),
    .io_Stationary_matrix_4_0(PathFinder_14_io_Stationary_matrix_4_0),
    .io_Stationary_matrix_4_1(PathFinder_14_io_Stationary_matrix_4_1),
    .io_Stationary_matrix_4_2(PathFinder_14_io_Stationary_matrix_4_2),
    .io_Stationary_matrix_4_3(PathFinder_14_io_Stationary_matrix_4_3),
    .io_Stationary_matrix_4_4(PathFinder_14_io_Stationary_matrix_4_4),
    .io_Stationary_matrix_4_5(PathFinder_14_io_Stationary_matrix_4_5),
    .io_Stationary_matrix_4_6(PathFinder_14_io_Stationary_matrix_4_6),
    .io_Stationary_matrix_4_7(PathFinder_14_io_Stationary_matrix_4_7),
    .io_Stationary_matrix_5_0(PathFinder_14_io_Stationary_matrix_5_0),
    .io_Stationary_matrix_5_1(PathFinder_14_io_Stationary_matrix_5_1),
    .io_Stationary_matrix_5_2(PathFinder_14_io_Stationary_matrix_5_2),
    .io_Stationary_matrix_5_3(PathFinder_14_io_Stationary_matrix_5_3),
    .io_Stationary_matrix_5_4(PathFinder_14_io_Stationary_matrix_5_4),
    .io_Stationary_matrix_5_5(PathFinder_14_io_Stationary_matrix_5_5),
    .io_Stationary_matrix_5_6(PathFinder_14_io_Stationary_matrix_5_6),
    .io_Stationary_matrix_5_7(PathFinder_14_io_Stationary_matrix_5_7),
    .io_Stationary_matrix_6_0(PathFinder_14_io_Stationary_matrix_6_0),
    .io_Stationary_matrix_6_1(PathFinder_14_io_Stationary_matrix_6_1),
    .io_Stationary_matrix_6_2(PathFinder_14_io_Stationary_matrix_6_2),
    .io_Stationary_matrix_6_3(PathFinder_14_io_Stationary_matrix_6_3),
    .io_Stationary_matrix_6_4(PathFinder_14_io_Stationary_matrix_6_4),
    .io_Stationary_matrix_6_5(PathFinder_14_io_Stationary_matrix_6_5),
    .io_Stationary_matrix_6_6(PathFinder_14_io_Stationary_matrix_6_6),
    .io_Stationary_matrix_6_7(PathFinder_14_io_Stationary_matrix_6_7),
    .io_Stationary_matrix_7_0(PathFinder_14_io_Stationary_matrix_7_0),
    .io_Stationary_matrix_7_1(PathFinder_14_io_Stationary_matrix_7_1),
    .io_Stationary_matrix_7_2(PathFinder_14_io_Stationary_matrix_7_2),
    .io_Stationary_matrix_7_3(PathFinder_14_io_Stationary_matrix_7_3),
    .io_Stationary_matrix_7_4(PathFinder_14_io_Stationary_matrix_7_4),
    .io_Stationary_matrix_7_5(PathFinder_14_io_Stationary_matrix_7_5),
    .io_Stationary_matrix_7_6(PathFinder_14_io_Stationary_matrix_7_6),
    .io_Stationary_matrix_7_7(PathFinder_14_io_Stationary_matrix_7_7),
    .io_Streaming_matrix_0(PathFinder_14_io_Streaming_matrix_0),
    .io_Streaming_matrix_1(PathFinder_14_io_Streaming_matrix_1),
    .io_Streaming_matrix_2(PathFinder_14_io_Streaming_matrix_2),
    .io_Streaming_matrix_3(PathFinder_14_io_Streaming_matrix_3),
    .io_Streaming_matrix_4(PathFinder_14_io_Streaming_matrix_4),
    .io_Streaming_matrix_5(PathFinder_14_io_Streaming_matrix_5),
    .io_Streaming_matrix_6(PathFinder_14_io_Streaming_matrix_6),
    .io_Streaming_matrix_7(PathFinder_14_io_Streaming_matrix_7),
    .io_i_mux_bus_0(PathFinder_14_io_i_mux_bus_0),
    .io_i_mux_bus_1(PathFinder_14_io_i_mux_bus_1),
    .io_i_mux_bus_2(PathFinder_14_io_i_mux_bus_2),
    .io_i_mux_bus_3(PathFinder_14_io_i_mux_bus_3),
    .io_Source_0(PathFinder_14_io_Source_0),
    .io_Source_1(PathFinder_14_io_Source_1),
    .io_Source_2(PathFinder_14_io_Source_2),
    .io_Source_3(PathFinder_14_io_Source_3),
    .io_destination_0(PathFinder_14_io_destination_0),
    .io_destination_1(PathFinder_14_io_destination_1),
    .io_destination_2(PathFinder_14_io_destination_2),
    .io_destination_3(PathFinder_14_io_destination_3),
    .io_PF_Valid(PathFinder_14_io_PF_Valid),
    .io_NoDPE(PathFinder_14_io_NoDPE),
    .io_DataValid(PathFinder_14_io_DataValid)
  );
  PathFinder PathFinder_15 ( // @[FlexDPU.scala 77:41]
    .clock(PathFinder_15_clock),
    .reset(PathFinder_15_reset),
    .io_Stationary_matrix_0_0(PathFinder_15_io_Stationary_matrix_0_0),
    .io_Stationary_matrix_0_1(PathFinder_15_io_Stationary_matrix_0_1),
    .io_Stationary_matrix_0_2(PathFinder_15_io_Stationary_matrix_0_2),
    .io_Stationary_matrix_0_3(PathFinder_15_io_Stationary_matrix_0_3),
    .io_Stationary_matrix_0_4(PathFinder_15_io_Stationary_matrix_0_4),
    .io_Stationary_matrix_0_5(PathFinder_15_io_Stationary_matrix_0_5),
    .io_Stationary_matrix_0_6(PathFinder_15_io_Stationary_matrix_0_6),
    .io_Stationary_matrix_0_7(PathFinder_15_io_Stationary_matrix_0_7),
    .io_Stationary_matrix_1_0(PathFinder_15_io_Stationary_matrix_1_0),
    .io_Stationary_matrix_1_1(PathFinder_15_io_Stationary_matrix_1_1),
    .io_Stationary_matrix_1_2(PathFinder_15_io_Stationary_matrix_1_2),
    .io_Stationary_matrix_1_3(PathFinder_15_io_Stationary_matrix_1_3),
    .io_Stationary_matrix_1_4(PathFinder_15_io_Stationary_matrix_1_4),
    .io_Stationary_matrix_1_5(PathFinder_15_io_Stationary_matrix_1_5),
    .io_Stationary_matrix_1_6(PathFinder_15_io_Stationary_matrix_1_6),
    .io_Stationary_matrix_1_7(PathFinder_15_io_Stationary_matrix_1_7),
    .io_Stationary_matrix_2_0(PathFinder_15_io_Stationary_matrix_2_0),
    .io_Stationary_matrix_2_1(PathFinder_15_io_Stationary_matrix_2_1),
    .io_Stationary_matrix_2_2(PathFinder_15_io_Stationary_matrix_2_2),
    .io_Stationary_matrix_2_3(PathFinder_15_io_Stationary_matrix_2_3),
    .io_Stationary_matrix_2_4(PathFinder_15_io_Stationary_matrix_2_4),
    .io_Stationary_matrix_2_5(PathFinder_15_io_Stationary_matrix_2_5),
    .io_Stationary_matrix_2_6(PathFinder_15_io_Stationary_matrix_2_6),
    .io_Stationary_matrix_2_7(PathFinder_15_io_Stationary_matrix_2_7),
    .io_Stationary_matrix_3_0(PathFinder_15_io_Stationary_matrix_3_0),
    .io_Stationary_matrix_3_1(PathFinder_15_io_Stationary_matrix_3_1),
    .io_Stationary_matrix_3_2(PathFinder_15_io_Stationary_matrix_3_2),
    .io_Stationary_matrix_3_3(PathFinder_15_io_Stationary_matrix_3_3),
    .io_Stationary_matrix_3_4(PathFinder_15_io_Stationary_matrix_3_4),
    .io_Stationary_matrix_3_5(PathFinder_15_io_Stationary_matrix_3_5),
    .io_Stationary_matrix_3_6(PathFinder_15_io_Stationary_matrix_3_6),
    .io_Stationary_matrix_3_7(PathFinder_15_io_Stationary_matrix_3_7),
    .io_Stationary_matrix_4_0(PathFinder_15_io_Stationary_matrix_4_0),
    .io_Stationary_matrix_4_1(PathFinder_15_io_Stationary_matrix_4_1),
    .io_Stationary_matrix_4_2(PathFinder_15_io_Stationary_matrix_4_2),
    .io_Stationary_matrix_4_3(PathFinder_15_io_Stationary_matrix_4_3),
    .io_Stationary_matrix_4_4(PathFinder_15_io_Stationary_matrix_4_4),
    .io_Stationary_matrix_4_5(PathFinder_15_io_Stationary_matrix_4_5),
    .io_Stationary_matrix_4_6(PathFinder_15_io_Stationary_matrix_4_6),
    .io_Stationary_matrix_4_7(PathFinder_15_io_Stationary_matrix_4_7),
    .io_Stationary_matrix_5_0(PathFinder_15_io_Stationary_matrix_5_0),
    .io_Stationary_matrix_5_1(PathFinder_15_io_Stationary_matrix_5_1),
    .io_Stationary_matrix_5_2(PathFinder_15_io_Stationary_matrix_5_2),
    .io_Stationary_matrix_5_3(PathFinder_15_io_Stationary_matrix_5_3),
    .io_Stationary_matrix_5_4(PathFinder_15_io_Stationary_matrix_5_4),
    .io_Stationary_matrix_5_5(PathFinder_15_io_Stationary_matrix_5_5),
    .io_Stationary_matrix_5_6(PathFinder_15_io_Stationary_matrix_5_6),
    .io_Stationary_matrix_5_7(PathFinder_15_io_Stationary_matrix_5_7),
    .io_Stationary_matrix_6_0(PathFinder_15_io_Stationary_matrix_6_0),
    .io_Stationary_matrix_6_1(PathFinder_15_io_Stationary_matrix_6_1),
    .io_Stationary_matrix_6_2(PathFinder_15_io_Stationary_matrix_6_2),
    .io_Stationary_matrix_6_3(PathFinder_15_io_Stationary_matrix_6_3),
    .io_Stationary_matrix_6_4(PathFinder_15_io_Stationary_matrix_6_4),
    .io_Stationary_matrix_6_5(PathFinder_15_io_Stationary_matrix_6_5),
    .io_Stationary_matrix_6_6(PathFinder_15_io_Stationary_matrix_6_6),
    .io_Stationary_matrix_6_7(PathFinder_15_io_Stationary_matrix_6_7),
    .io_Stationary_matrix_7_0(PathFinder_15_io_Stationary_matrix_7_0),
    .io_Stationary_matrix_7_1(PathFinder_15_io_Stationary_matrix_7_1),
    .io_Stationary_matrix_7_2(PathFinder_15_io_Stationary_matrix_7_2),
    .io_Stationary_matrix_7_3(PathFinder_15_io_Stationary_matrix_7_3),
    .io_Stationary_matrix_7_4(PathFinder_15_io_Stationary_matrix_7_4),
    .io_Stationary_matrix_7_5(PathFinder_15_io_Stationary_matrix_7_5),
    .io_Stationary_matrix_7_6(PathFinder_15_io_Stationary_matrix_7_6),
    .io_Stationary_matrix_7_7(PathFinder_15_io_Stationary_matrix_7_7),
    .io_Streaming_matrix_0(PathFinder_15_io_Streaming_matrix_0),
    .io_Streaming_matrix_1(PathFinder_15_io_Streaming_matrix_1),
    .io_Streaming_matrix_2(PathFinder_15_io_Streaming_matrix_2),
    .io_Streaming_matrix_3(PathFinder_15_io_Streaming_matrix_3),
    .io_Streaming_matrix_4(PathFinder_15_io_Streaming_matrix_4),
    .io_Streaming_matrix_5(PathFinder_15_io_Streaming_matrix_5),
    .io_Streaming_matrix_6(PathFinder_15_io_Streaming_matrix_6),
    .io_Streaming_matrix_7(PathFinder_15_io_Streaming_matrix_7),
    .io_i_mux_bus_0(PathFinder_15_io_i_mux_bus_0),
    .io_i_mux_bus_1(PathFinder_15_io_i_mux_bus_1),
    .io_i_mux_bus_2(PathFinder_15_io_i_mux_bus_2),
    .io_i_mux_bus_3(PathFinder_15_io_i_mux_bus_3),
    .io_Source_0(PathFinder_15_io_Source_0),
    .io_Source_1(PathFinder_15_io_Source_1),
    .io_Source_2(PathFinder_15_io_Source_2),
    .io_Source_3(PathFinder_15_io_Source_3),
    .io_destination_0(PathFinder_15_io_destination_0),
    .io_destination_1(PathFinder_15_io_destination_1),
    .io_destination_2(PathFinder_15_io_destination_2),
    .io_destination_3(PathFinder_15_io_destination_3),
    .io_PF_Valid(PathFinder_15_io_PF_Valid),
    .io_NoDPE(PathFinder_15_io_NoDPE),
    .io_DataValid(PathFinder_15_io_DataValid)
  );
  flexdpecom4 flexdpecom4 ( // @[FlexDPU.scala 110:47]
    .clock(flexdpecom4_clock),
    .reset(flexdpecom4_reset),
    .io_i_data_valid(flexdpecom4_io_i_data_valid),
    .io_i_data_bus_0(flexdpecom4_io_i_data_bus_0),
    .io_i_data_bus_1(flexdpecom4_io_i_data_bus_1),
    .io_i_data_bus_2(flexdpecom4_io_i_data_bus_2),
    .io_i_data_bus_3(flexdpecom4_io_i_data_bus_3),
    .io_i_data_bus2_0(flexdpecom4_io_i_data_bus2_0),
    .io_i_data_bus2_1(flexdpecom4_io_i_data_bus2_1),
    .io_i_data_bus2_2(flexdpecom4_io_i_data_bus2_2),
    .io_i_data_bus2_3(flexdpecom4_io_i_data_bus2_3),
    .io_o_adder_0(flexdpecom4_io_o_adder_0),
    .io_o_adder_1(flexdpecom4_io_o_adder_1),
    .io_o_adder_2(flexdpecom4_io_o_adder_2),
    .io_i_mux_bus_0(flexdpecom4_io_i_mux_bus_0),
    .io_i_mux_bus_1(flexdpecom4_io_i_mux_bus_1),
    .io_i_mux_bus_2(flexdpecom4_io_i_mux_bus_2),
    .io_i_mux_bus_3(flexdpecom4_io_i_mux_bus_3)
  );
  flexdpecom4 flexdpecom4_1 ( // @[FlexDPU.scala 110:47]
    .clock(flexdpecom4_1_clock),
    .reset(flexdpecom4_1_reset),
    .io_i_data_valid(flexdpecom4_1_io_i_data_valid),
    .io_i_data_bus_0(flexdpecom4_1_io_i_data_bus_0),
    .io_i_data_bus_1(flexdpecom4_1_io_i_data_bus_1),
    .io_i_data_bus_2(flexdpecom4_1_io_i_data_bus_2),
    .io_i_data_bus_3(flexdpecom4_1_io_i_data_bus_3),
    .io_i_data_bus2_0(flexdpecom4_1_io_i_data_bus2_0),
    .io_i_data_bus2_1(flexdpecom4_1_io_i_data_bus2_1),
    .io_i_data_bus2_2(flexdpecom4_1_io_i_data_bus2_2),
    .io_i_data_bus2_3(flexdpecom4_1_io_i_data_bus2_3),
    .io_o_adder_0(flexdpecom4_1_io_o_adder_0),
    .io_o_adder_1(flexdpecom4_1_io_o_adder_1),
    .io_o_adder_2(flexdpecom4_1_io_o_adder_2),
    .io_i_mux_bus_0(flexdpecom4_1_io_i_mux_bus_0),
    .io_i_mux_bus_1(flexdpecom4_1_io_i_mux_bus_1),
    .io_i_mux_bus_2(flexdpecom4_1_io_i_mux_bus_2),
    .io_i_mux_bus_3(flexdpecom4_1_io_i_mux_bus_3)
  );
  flexdpecom4 flexdpecom4_2 ( // @[FlexDPU.scala 110:47]
    .clock(flexdpecom4_2_clock),
    .reset(flexdpecom4_2_reset),
    .io_i_data_valid(flexdpecom4_2_io_i_data_valid),
    .io_i_data_bus_0(flexdpecom4_2_io_i_data_bus_0),
    .io_i_data_bus_1(flexdpecom4_2_io_i_data_bus_1),
    .io_i_data_bus_2(flexdpecom4_2_io_i_data_bus_2),
    .io_i_data_bus_3(flexdpecom4_2_io_i_data_bus_3),
    .io_i_data_bus2_0(flexdpecom4_2_io_i_data_bus2_0),
    .io_i_data_bus2_1(flexdpecom4_2_io_i_data_bus2_1),
    .io_i_data_bus2_2(flexdpecom4_2_io_i_data_bus2_2),
    .io_i_data_bus2_3(flexdpecom4_2_io_i_data_bus2_3),
    .io_o_adder_0(flexdpecom4_2_io_o_adder_0),
    .io_o_adder_1(flexdpecom4_2_io_o_adder_1),
    .io_o_adder_2(flexdpecom4_2_io_o_adder_2),
    .io_i_mux_bus_0(flexdpecom4_2_io_i_mux_bus_0),
    .io_i_mux_bus_1(flexdpecom4_2_io_i_mux_bus_1),
    .io_i_mux_bus_2(flexdpecom4_2_io_i_mux_bus_2),
    .io_i_mux_bus_3(flexdpecom4_2_io_i_mux_bus_3)
  );
  flexdpecom4 flexdpecom4_3 ( // @[FlexDPU.scala 110:47]
    .clock(flexdpecom4_3_clock),
    .reset(flexdpecom4_3_reset),
    .io_i_data_valid(flexdpecom4_3_io_i_data_valid),
    .io_i_data_bus_0(flexdpecom4_3_io_i_data_bus_0),
    .io_i_data_bus_1(flexdpecom4_3_io_i_data_bus_1),
    .io_i_data_bus_2(flexdpecom4_3_io_i_data_bus_2),
    .io_i_data_bus_3(flexdpecom4_3_io_i_data_bus_3),
    .io_i_data_bus2_0(flexdpecom4_3_io_i_data_bus2_0),
    .io_i_data_bus2_1(flexdpecom4_3_io_i_data_bus2_1),
    .io_i_data_bus2_2(flexdpecom4_3_io_i_data_bus2_2),
    .io_i_data_bus2_3(flexdpecom4_3_io_i_data_bus2_3),
    .io_o_adder_0(flexdpecom4_3_io_o_adder_0),
    .io_o_adder_1(flexdpecom4_3_io_o_adder_1),
    .io_o_adder_2(flexdpecom4_3_io_o_adder_2),
    .io_i_mux_bus_0(flexdpecom4_3_io_i_mux_bus_0),
    .io_i_mux_bus_1(flexdpecom4_3_io_i_mux_bus_1),
    .io_i_mux_bus_2(flexdpecom4_3_io_i_mux_bus_2),
    .io_i_mux_bus_3(flexdpecom4_3_io_i_mux_bus_3)
  );
  flexdpecom4 flexdpecom4_4 ( // @[FlexDPU.scala 110:47]
    .clock(flexdpecom4_4_clock),
    .reset(flexdpecom4_4_reset),
    .io_i_data_valid(flexdpecom4_4_io_i_data_valid),
    .io_i_data_bus_0(flexdpecom4_4_io_i_data_bus_0),
    .io_i_data_bus_1(flexdpecom4_4_io_i_data_bus_1),
    .io_i_data_bus_2(flexdpecom4_4_io_i_data_bus_2),
    .io_i_data_bus_3(flexdpecom4_4_io_i_data_bus_3),
    .io_i_data_bus2_0(flexdpecom4_4_io_i_data_bus2_0),
    .io_i_data_bus2_1(flexdpecom4_4_io_i_data_bus2_1),
    .io_i_data_bus2_2(flexdpecom4_4_io_i_data_bus2_2),
    .io_i_data_bus2_3(flexdpecom4_4_io_i_data_bus2_3),
    .io_o_adder_0(flexdpecom4_4_io_o_adder_0),
    .io_o_adder_1(flexdpecom4_4_io_o_adder_1),
    .io_o_adder_2(flexdpecom4_4_io_o_adder_2),
    .io_i_mux_bus_0(flexdpecom4_4_io_i_mux_bus_0),
    .io_i_mux_bus_1(flexdpecom4_4_io_i_mux_bus_1),
    .io_i_mux_bus_2(flexdpecom4_4_io_i_mux_bus_2),
    .io_i_mux_bus_3(flexdpecom4_4_io_i_mux_bus_3)
  );
  flexdpecom4 flexdpecom4_5 ( // @[FlexDPU.scala 110:47]
    .clock(flexdpecom4_5_clock),
    .reset(flexdpecom4_5_reset),
    .io_i_data_valid(flexdpecom4_5_io_i_data_valid),
    .io_i_data_bus_0(flexdpecom4_5_io_i_data_bus_0),
    .io_i_data_bus_1(flexdpecom4_5_io_i_data_bus_1),
    .io_i_data_bus_2(flexdpecom4_5_io_i_data_bus_2),
    .io_i_data_bus_3(flexdpecom4_5_io_i_data_bus_3),
    .io_i_data_bus2_0(flexdpecom4_5_io_i_data_bus2_0),
    .io_i_data_bus2_1(flexdpecom4_5_io_i_data_bus2_1),
    .io_i_data_bus2_2(flexdpecom4_5_io_i_data_bus2_2),
    .io_i_data_bus2_3(flexdpecom4_5_io_i_data_bus2_3),
    .io_o_adder_0(flexdpecom4_5_io_o_adder_0),
    .io_o_adder_1(flexdpecom4_5_io_o_adder_1),
    .io_o_adder_2(flexdpecom4_5_io_o_adder_2),
    .io_i_mux_bus_0(flexdpecom4_5_io_i_mux_bus_0),
    .io_i_mux_bus_1(flexdpecom4_5_io_i_mux_bus_1),
    .io_i_mux_bus_2(flexdpecom4_5_io_i_mux_bus_2),
    .io_i_mux_bus_3(flexdpecom4_5_io_i_mux_bus_3)
  );
  flexdpecom4 flexdpecom4_6 ( // @[FlexDPU.scala 110:47]
    .clock(flexdpecom4_6_clock),
    .reset(flexdpecom4_6_reset),
    .io_i_data_valid(flexdpecom4_6_io_i_data_valid),
    .io_i_data_bus_0(flexdpecom4_6_io_i_data_bus_0),
    .io_i_data_bus_1(flexdpecom4_6_io_i_data_bus_1),
    .io_i_data_bus_2(flexdpecom4_6_io_i_data_bus_2),
    .io_i_data_bus_3(flexdpecom4_6_io_i_data_bus_3),
    .io_i_data_bus2_0(flexdpecom4_6_io_i_data_bus2_0),
    .io_i_data_bus2_1(flexdpecom4_6_io_i_data_bus2_1),
    .io_i_data_bus2_2(flexdpecom4_6_io_i_data_bus2_2),
    .io_i_data_bus2_3(flexdpecom4_6_io_i_data_bus2_3),
    .io_o_adder_0(flexdpecom4_6_io_o_adder_0),
    .io_o_adder_1(flexdpecom4_6_io_o_adder_1),
    .io_o_adder_2(flexdpecom4_6_io_o_adder_2),
    .io_i_mux_bus_0(flexdpecom4_6_io_i_mux_bus_0),
    .io_i_mux_bus_1(flexdpecom4_6_io_i_mux_bus_1),
    .io_i_mux_bus_2(flexdpecom4_6_io_i_mux_bus_2),
    .io_i_mux_bus_3(flexdpecom4_6_io_i_mux_bus_3)
  );
  flexdpecom4 flexdpecom4_7 ( // @[FlexDPU.scala 110:47]
    .clock(flexdpecom4_7_clock),
    .reset(flexdpecom4_7_reset),
    .io_i_data_valid(flexdpecom4_7_io_i_data_valid),
    .io_i_data_bus_0(flexdpecom4_7_io_i_data_bus_0),
    .io_i_data_bus_1(flexdpecom4_7_io_i_data_bus_1),
    .io_i_data_bus_2(flexdpecom4_7_io_i_data_bus_2),
    .io_i_data_bus_3(flexdpecom4_7_io_i_data_bus_3),
    .io_i_data_bus2_0(flexdpecom4_7_io_i_data_bus2_0),
    .io_i_data_bus2_1(flexdpecom4_7_io_i_data_bus2_1),
    .io_i_data_bus2_2(flexdpecom4_7_io_i_data_bus2_2),
    .io_i_data_bus2_3(flexdpecom4_7_io_i_data_bus2_3),
    .io_o_adder_0(flexdpecom4_7_io_o_adder_0),
    .io_o_adder_1(flexdpecom4_7_io_o_adder_1),
    .io_o_adder_2(flexdpecom4_7_io_o_adder_2),
    .io_i_mux_bus_0(flexdpecom4_7_io_i_mux_bus_0),
    .io_i_mux_bus_1(flexdpecom4_7_io_i_mux_bus_1),
    .io_i_mux_bus_2(flexdpecom4_7_io_i_mux_bus_2),
    .io_i_mux_bus_3(flexdpecom4_7_io_i_mux_bus_3)
  );
  flexdpecom4 flexdpecom4_8 ( // @[FlexDPU.scala 110:47]
    .clock(flexdpecom4_8_clock),
    .reset(flexdpecom4_8_reset),
    .io_i_data_valid(flexdpecom4_8_io_i_data_valid),
    .io_i_data_bus_0(flexdpecom4_8_io_i_data_bus_0),
    .io_i_data_bus_1(flexdpecom4_8_io_i_data_bus_1),
    .io_i_data_bus_2(flexdpecom4_8_io_i_data_bus_2),
    .io_i_data_bus_3(flexdpecom4_8_io_i_data_bus_3),
    .io_i_data_bus2_0(flexdpecom4_8_io_i_data_bus2_0),
    .io_i_data_bus2_1(flexdpecom4_8_io_i_data_bus2_1),
    .io_i_data_bus2_2(flexdpecom4_8_io_i_data_bus2_2),
    .io_i_data_bus2_3(flexdpecom4_8_io_i_data_bus2_3),
    .io_o_adder_0(flexdpecom4_8_io_o_adder_0),
    .io_o_adder_1(flexdpecom4_8_io_o_adder_1),
    .io_o_adder_2(flexdpecom4_8_io_o_adder_2),
    .io_i_mux_bus_0(flexdpecom4_8_io_i_mux_bus_0),
    .io_i_mux_bus_1(flexdpecom4_8_io_i_mux_bus_1),
    .io_i_mux_bus_2(flexdpecom4_8_io_i_mux_bus_2),
    .io_i_mux_bus_3(flexdpecom4_8_io_i_mux_bus_3)
  );
  flexdpecom4 flexdpecom4_9 ( // @[FlexDPU.scala 110:47]
    .clock(flexdpecom4_9_clock),
    .reset(flexdpecom4_9_reset),
    .io_i_data_valid(flexdpecom4_9_io_i_data_valid),
    .io_i_data_bus_0(flexdpecom4_9_io_i_data_bus_0),
    .io_i_data_bus_1(flexdpecom4_9_io_i_data_bus_1),
    .io_i_data_bus_2(flexdpecom4_9_io_i_data_bus_2),
    .io_i_data_bus_3(flexdpecom4_9_io_i_data_bus_3),
    .io_i_data_bus2_0(flexdpecom4_9_io_i_data_bus2_0),
    .io_i_data_bus2_1(flexdpecom4_9_io_i_data_bus2_1),
    .io_i_data_bus2_2(flexdpecom4_9_io_i_data_bus2_2),
    .io_i_data_bus2_3(flexdpecom4_9_io_i_data_bus2_3),
    .io_o_adder_0(flexdpecom4_9_io_o_adder_0),
    .io_o_adder_1(flexdpecom4_9_io_o_adder_1),
    .io_o_adder_2(flexdpecom4_9_io_o_adder_2),
    .io_i_mux_bus_0(flexdpecom4_9_io_i_mux_bus_0),
    .io_i_mux_bus_1(flexdpecom4_9_io_i_mux_bus_1),
    .io_i_mux_bus_2(flexdpecom4_9_io_i_mux_bus_2),
    .io_i_mux_bus_3(flexdpecom4_9_io_i_mux_bus_3)
  );
  flexdpecom4 flexdpecom4_10 ( // @[FlexDPU.scala 110:47]
    .clock(flexdpecom4_10_clock),
    .reset(flexdpecom4_10_reset),
    .io_i_data_valid(flexdpecom4_10_io_i_data_valid),
    .io_i_data_bus_0(flexdpecom4_10_io_i_data_bus_0),
    .io_i_data_bus_1(flexdpecom4_10_io_i_data_bus_1),
    .io_i_data_bus_2(flexdpecom4_10_io_i_data_bus_2),
    .io_i_data_bus_3(flexdpecom4_10_io_i_data_bus_3),
    .io_i_data_bus2_0(flexdpecom4_10_io_i_data_bus2_0),
    .io_i_data_bus2_1(flexdpecom4_10_io_i_data_bus2_1),
    .io_i_data_bus2_2(flexdpecom4_10_io_i_data_bus2_2),
    .io_i_data_bus2_3(flexdpecom4_10_io_i_data_bus2_3),
    .io_o_adder_0(flexdpecom4_10_io_o_adder_0),
    .io_o_adder_1(flexdpecom4_10_io_o_adder_1),
    .io_o_adder_2(flexdpecom4_10_io_o_adder_2),
    .io_i_mux_bus_0(flexdpecom4_10_io_i_mux_bus_0),
    .io_i_mux_bus_1(flexdpecom4_10_io_i_mux_bus_1),
    .io_i_mux_bus_2(flexdpecom4_10_io_i_mux_bus_2),
    .io_i_mux_bus_3(flexdpecom4_10_io_i_mux_bus_3)
  );
  flexdpecom4 flexdpecom4_11 ( // @[FlexDPU.scala 110:47]
    .clock(flexdpecom4_11_clock),
    .reset(flexdpecom4_11_reset),
    .io_i_data_valid(flexdpecom4_11_io_i_data_valid),
    .io_i_data_bus_0(flexdpecom4_11_io_i_data_bus_0),
    .io_i_data_bus_1(flexdpecom4_11_io_i_data_bus_1),
    .io_i_data_bus_2(flexdpecom4_11_io_i_data_bus_2),
    .io_i_data_bus_3(flexdpecom4_11_io_i_data_bus_3),
    .io_i_data_bus2_0(flexdpecom4_11_io_i_data_bus2_0),
    .io_i_data_bus2_1(flexdpecom4_11_io_i_data_bus2_1),
    .io_i_data_bus2_2(flexdpecom4_11_io_i_data_bus2_2),
    .io_i_data_bus2_3(flexdpecom4_11_io_i_data_bus2_3),
    .io_o_adder_0(flexdpecom4_11_io_o_adder_0),
    .io_o_adder_1(flexdpecom4_11_io_o_adder_1),
    .io_o_adder_2(flexdpecom4_11_io_o_adder_2),
    .io_i_mux_bus_0(flexdpecom4_11_io_i_mux_bus_0),
    .io_i_mux_bus_1(flexdpecom4_11_io_i_mux_bus_1),
    .io_i_mux_bus_2(flexdpecom4_11_io_i_mux_bus_2),
    .io_i_mux_bus_3(flexdpecom4_11_io_i_mux_bus_3)
  );
  flexdpecom4 flexdpecom4_12 ( // @[FlexDPU.scala 110:47]
    .clock(flexdpecom4_12_clock),
    .reset(flexdpecom4_12_reset),
    .io_i_data_valid(flexdpecom4_12_io_i_data_valid),
    .io_i_data_bus_0(flexdpecom4_12_io_i_data_bus_0),
    .io_i_data_bus_1(flexdpecom4_12_io_i_data_bus_1),
    .io_i_data_bus_2(flexdpecom4_12_io_i_data_bus_2),
    .io_i_data_bus_3(flexdpecom4_12_io_i_data_bus_3),
    .io_i_data_bus2_0(flexdpecom4_12_io_i_data_bus2_0),
    .io_i_data_bus2_1(flexdpecom4_12_io_i_data_bus2_1),
    .io_i_data_bus2_2(flexdpecom4_12_io_i_data_bus2_2),
    .io_i_data_bus2_3(flexdpecom4_12_io_i_data_bus2_3),
    .io_o_adder_0(flexdpecom4_12_io_o_adder_0),
    .io_o_adder_1(flexdpecom4_12_io_o_adder_1),
    .io_o_adder_2(flexdpecom4_12_io_o_adder_2),
    .io_i_mux_bus_0(flexdpecom4_12_io_i_mux_bus_0),
    .io_i_mux_bus_1(flexdpecom4_12_io_i_mux_bus_1),
    .io_i_mux_bus_2(flexdpecom4_12_io_i_mux_bus_2),
    .io_i_mux_bus_3(flexdpecom4_12_io_i_mux_bus_3)
  );
  flexdpecom4 flexdpecom4_13 ( // @[FlexDPU.scala 110:47]
    .clock(flexdpecom4_13_clock),
    .reset(flexdpecom4_13_reset),
    .io_i_data_valid(flexdpecom4_13_io_i_data_valid),
    .io_i_data_bus_0(flexdpecom4_13_io_i_data_bus_0),
    .io_i_data_bus_1(flexdpecom4_13_io_i_data_bus_1),
    .io_i_data_bus_2(flexdpecom4_13_io_i_data_bus_2),
    .io_i_data_bus_3(flexdpecom4_13_io_i_data_bus_3),
    .io_i_data_bus2_0(flexdpecom4_13_io_i_data_bus2_0),
    .io_i_data_bus2_1(flexdpecom4_13_io_i_data_bus2_1),
    .io_i_data_bus2_2(flexdpecom4_13_io_i_data_bus2_2),
    .io_i_data_bus2_3(flexdpecom4_13_io_i_data_bus2_3),
    .io_o_adder_0(flexdpecom4_13_io_o_adder_0),
    .io_o_adder_1(flexdpecom4_13_io_o_adder_1),
    .io_o_adder_2(flexdpecom4_13_io_o_adder_2),
    .io_i_mux_bus_0(flexdpecom4_13_io_i_mux_bus_0),
    .io_i_mux_bus_1(flexdpecom4_13_io_i_mux_bus_1),
    .io_i_mux_bus_2(flexdpecom4_13_io_i_mux_bus_2),
    .io_i_mux_bus_3(flexdpecom4_13_io_i_mux_bus_3)
  );
  flexdpecom4 flexdpecom4_14 ( // @[FlexDPU.scala 110:47]
    .clock(flexdpecom4_14_clock),
    .reset(flexdpecom4_14_reset),
    .io_i_data_valid(flexdpecom4_14_io_i_data_valid),
    .io_i_data_bus_0(flexdpecom4_14_io_i_data_bus_0),
    .io_i_data_bus_1(flexdpecom4_14_io_i_data_bus_1),
    .io_i_data_bus_2(flexdpecom4_14_io_i_data_bus_2),
    .io_i_data_bus_3(flexdpecom4_14_io_i_data_bus_3),
    .io_i_data_bus2_0(flexdpecom4_14_io_i_data_bus2_0),
    .io_i_data_bus2_1(flexdpecom4_14_io_i_data_bus2_1),
    .io_i_data_bus2_2(flexdpecom4_14_io_i_data_bus2_2),
    .io_i_data_bus2_3(flexdpecom4_14_io_i_data_bus2_3),
    .io_o_adder_0(flexdpecom4_14_io_o_adder_0),
    .io_o_adder_1(flexdpecom4_14_io_o_adder_1),
    .io_o_adder_2(flexdpecom4_14_io_o_adder_2),
    .io_i_mux_bus_0(flexdpecom4_14_io_i_mux_bus_0),
    .io_i_mux_bus_1(flexdpecom4_14_io_i_mux_bus_1),
    .io_i_mux_bus_2(flexdpecom4_14_io_i_mux_bus_2),
    .io_i_mux_bus_3(flexdpecom4_14_io_i_mux_bus_3)
  );
  flexdpecom4 flexdpecom4_15 ( // @[FlexDPU.scala 110:47]
    .clock(flexdpecom4_15_clock),
    .reset(flexdpecom4_15_reset),
    .io_i_data_valid(flexdpecom4_15_io_i_data_valid),
    .io_i_data_bus_0(flexdpecom4_15_io_i_data_bus_0),
    .io_i_data_bus_1(flexdpecom4_15_io_i_data_bus_1),
    .io_i_data_bus_2(flexdpecom4_15_io_i_data_bus_2),
    .io_i_data_bus_3(flexdpecom4_15_io_i_data_bus_3),
    .io_i_data_bus2_0(flexdpecom4_15_io_i_data_bus2_0),
    .io_i_data_bus2_1(flexdpecom4_15_io_i_data_bus2_1),
    .io_i_data_bus2_2(flexdpecom4_15_io_i_data_bus2_2),
    .io_i_data_bus2_3(flexdpecom4_15_io_i_data_bus2_3),
    .io_o_adder_0(flexdpecom4_15_io_o_adder_0),
    .io_o_adder_1(flexdpecom4_15_io_o_adder_1),
    .io_o_adder_2(flexdpecom4_15_io_o_adder_2),
    .io_i_mux_bus_0(flexdpecom4_15_io_i_mux_bus_0),
    .io_i_mux_bus_1(flexdpecom4_15_io_i_mux_bus_1),
    .io_i_mux_bus_2(flexdpecom4_15_io_i_mux_bus_2),
    .io_i_mux_bus_3(flexdpecom4_15_io_i_mux_bus_3)
  );
  assign io_output_0_0 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_0_1 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_0_2 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_0_3 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_0_4 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_0_5 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_0_6 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_0_7 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_1_0 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_1_1 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_1_2 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_1_3 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_1_4 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_1_5 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_1_6 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_1_7 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_2_0 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_2_1 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_2_2 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_2_3 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_2_4 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_2_5 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_2_6 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_2_7 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_3_0 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_3_1 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_3_2 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_3_3 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_3_4 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_3_5 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_3_6 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_3_7 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_4_0 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_4_1 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_4_2 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_4_3 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_4_4 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_4_5 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_4_6 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_4_7 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_5_0 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_5_1 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_5_2 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_5_3 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_5_4 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_5_5 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_5_6 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_5_7 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_6_0 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_6_1 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_6_2 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_6_3 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_6_4 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_6_5 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_6_6 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_6_7 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_7_0 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_7_1 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_7_2 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_7_3 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_7_4 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_7_5 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_7_6 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign io_output_7_7 = 16'h0; // @[FlexDPU.scala 18:{67,67}]
  assign PathFinder_clock = clock;
  assign PathFinder_reset = reset;
  assign PathFinder_io_Stationary_matrix_0_0 = Statvalid ? io_Stationary_matrix_0_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_0_1 = Statvalid ? io_Stationary_matrix_0_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_0_2 = Statvalid ? io_Stationary_matrix_0_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_0_3 = Statvalid ? io_Stationary_matrix_0_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_0_4 = Statvalid ? io_Stationary_matrix_0_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_0_5 = Statvalid ? io_Stationary_matrix_0_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_0_6 = Statvalid ? io_Stationary_matrix_0_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_0_7 = Statvalid ? io_Stationary_matrix_0_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_1_0 = Statvalid ? io_Stationary_matrix_1_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_1_1 = Statvalid ? io_Stationary_matrix_1_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_1_2 = Statvalid ? io_Stationary_matrix_1_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_1_3 = Statvalid ? io_Stationary_matrix_1_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_1_4 = Statvalid ? io_Stationary_matrix_1_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_1_5 = Statvalid ? io_Stationary_matrix_1_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_1_6 = Statvalid ? io_Stationary_matrix_1_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_1_7 = Statvalid ? io_Stationary_matrix_1_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_2_0 = Statvalid ? io_Stationary_matrix_2_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_2_1 = Statvalid ? io_Stationary_matrix_2_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_2_2 = Statvalid ? io_Stationary_matrix_2_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_2_3 = Statvalid ? io_Stationary_matrix_2_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_2_4 = Statvalid ? io_Stationary_matrix_2_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_2_5 = Statvalid ? io_Stationary_matrix_2_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_2_6 = Statvalid ? io_Stationary_matrix_2_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_2_7 = Statvalid ? io_Stationary_matrix_2_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_3_0 = Statvalid ? io_Stationary_matrix_3_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_3_1 = Statvalid ? io_Stationary_matrix_3_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_3_2 = Statvalid ? io_Stationary_matrix_3_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_3_3 = Statvalid ? io_Stationary_matrix_3_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_3_4 = Statvalid ? io_Stationary_matrix_3_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_3_5 = Statvalid ? io_Stationary_matrix_3_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_3_6 = Statvalid ? io_Stationary_matrix_3_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_3_7 = Statvalid ? io_Stationary_matrix_3_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_4_0 = Statvalid ? io_Stationary_matrix_4_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_4_1 = Statvalid ? io_Stationary_matrix_4_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_4_2 = Statvalid ? io_Stationary_matrix_4_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_4_3 = Statvalid ? io_Stationary_matrix_4_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_4_4 = Statvalid ? io_Stationary_matrix_4_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_4_5 = Statvalid ? io_Stationary_matrix_4_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_4_6 = Statvalid ? io_Stationary_matrix_4_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_4_7 = Statvalid ? io_Stationary_matrix_4_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_5_0 = Statvalid ? io_Stationary_matrix_5_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_5_1 = Statvalid ? io_Stationary_matrix_5_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_5_2 = Statvalid ? io_Stationary_matrix_5_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_5_3 = Statvalid ? io_Stationary_matrix_5_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_5_4 = Statvalid ? io_Stationary_matrix_5_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_5_5 = Statvalid ? io_Stationary_matrix_5_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_5_6 = Statvalid ? io_Stationary_matrix_5_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_5_7 = Statvalid ? io_Stationary_matrix_5_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_6_0 = Statvalid ? io_Stationary_matrix_6_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_6_1 = Statvalid ? io_Stationary_matrix_6_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_6_2 = Statvalid ? io_Stationary_matrix_6_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_6_3 = Statvalid ? io_Stationary_matrix_6_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_6_4 = Statvalid ? io_Stationary_matrix_6_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_6_5 = Statvalid ? io_Stationary_matrix_6_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_6_6 = Statvalid ? io_Stationary_matrix_6_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_6_7 = Statvalid ? io_Stationary_matrix_6_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_7_0 = Statvalid ? io_Stationary_matrix_7_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_7_1 = Statvalid ? io_Stationary_matrix_7_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_7_2 = Statvalid ? io_Stationary_matrix_7_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_7_3 = Statvalid ? io_Stationary_matrix_7_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_7_4 = Statvalid ? io_Stationary_matrix_7_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_7_5 = Statvalid ? io_Stationary_matrix_7_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_7_6 = Statvalid ? io_Stationary_matrix_7_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Stationary_matrix_7_7 = Statvalid ? io_Stationary_matrix_7_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_io_Streaming_matrix_0 = _GEN_392[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_io_Streaming_matrix_1 = _GEN_393[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_io_Streaming_matrix_2 = _GEN_394[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_io_Streaming_matrix_3 = _GEN_395[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_io_Streaming_matrix_4 = _GEN_396[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_io_Streaming_matrix_5 = _GEN_397[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_io_Streaming_matrix_6 = _GEN_398[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_io_Streaming_matrix_7 = _GEN_399[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_io_NoDPE = 32'h0; // @[FlexDPU.scala 77:21]
  assign PathFinder_io_DataValid = Statvalid; // @[FlexDPU.scala 98:20 101:25 81:25]
  assign PathFinder_1_clock = clock;
  assign PathFinder_1_reset = reset;
  assign PathFinder_1_io_Stationary_matrix_0_0 = Statvalid ? io_Stationary_matrix_0_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_0_1 = Statvalid ? io_Stationary_matrix_0_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_0_2 = Statvalid ? io_Stationary_matrix_0_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_0_3 = Statvalid ? io_Stationary_matrix_0_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_0_4 = Statvalid ? io_Stationary_matrix_0_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_0_5 = Statvalid ? io_Stationary_matrix_0_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_0_6 = Statvalid ? io_Stationary_matrix_0_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_0_7 = Statvalid ? io_Stationary_matrix_0_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_1_0 = Statvalid ? io_Stationary_matrix_1_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_1_1 = Statvalid ? io_Stationary_matrix_1_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_1_2 = Statvalid ? io_Stationary_matrix_1_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_1_3 = Statvalid ? io_Stationary_matrix_1_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_1_4 = Statvalid ? io_Stationary_matrix_1_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_1_5 = Statvalid ? io_Stationary_matrix_1_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_1_6 = Statvalid ? io_Stationary_matrix_1_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_1_7 = Statvalid ? io_Stationary_matrix_1_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_2_0 = Statvalid ? io_Stationary_matrix_2_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_2_1 = Statvalid ? io_Stationary_matrix_2_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_2_2 = Statvalid ? io_Stationary_matrix_2_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_2_3 = Statvalid ? io_Stationary_matrix_2_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_2_4 = Statvalid ? io_Stationary_matrix_2_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_2_5 = Statvalid ? io_Stationary_matrix_2_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_2_6 = Statvalid ? io_Stationary_matrix_2_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_2_7 = Statvalid ? io_Stationary_matrix_2_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_3_0 = Statvalid ? io_Stationary_matrix_3_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_3_1 = Statvalid ? io_Stationary_matrix_3_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_3_2 = Statvalid ? io_Stationary_matrix_3_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_3_3 = Statvalid ? io_Stationary_matrix_3_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_3_4 = Statvalid ? io_Stationary_matrix_3_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_3_5 = Statvalid ? io_Stationary_matrix_3_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_3_6 = Statvalid ? io_Stationary_matrix_3_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_3_7 = Statvalid ? io_Stationary_matrix_3_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_4_0 = Statvalid ? io_Stationary_matrix_4_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_4_1 = Statvalid ? io_Stationary_matrix_4_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_4_2 = Statvalid ? io_Stationary_matrix_4_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_4_3 = Statvalid ? io_Stationary_matrix_4_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_4_4 = Statvalid ? io_Stationary_matrix_4_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_4_5 = Statvalid ? io_Stationary_matrix_4_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_4_6 = Statvalid ? io_Stationary_matrix_4_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_4_7 = Statvalid ? io_Stationary_matrix_4_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_5_0 = Statvalid ? io_Stationary_matrix_5_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_5_1 = Statvalid ? io_Stationary_matrix_5_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_5_2 = Statvalid ? io_Stationary_matrix_5_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_5_3 = Statvalid ? io_Stationary_matrix_5_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_5_4 = Statvalid ? io_Stationary_matrix_5_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_5_5 = Statvalid ? io_Stationary_matrix_5_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_5_6 = Statvalid ? io_Stationary_matrix_5_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_5_7 = Statvalid ? io_Stationary_matrix_5_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_6_0 = Statvalid ? io_Stationary_matrix_6_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_6_1 = Statvalid ? io_Stationary_matrix_6_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_6_2 = Statvalid ? io_Stationary_matrix_6_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_6_3 = Statvalid ? io_Stationary_matrix_6_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_6_4 = Statvalid ? io_Stationary_matrix_6_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_6_5 = Statvalid ? io_Stationary_matrix_6_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_6_6 = Statvalid ? io_Stationary_matrix_6_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_6_7 = Statvalid ? io_Stationary_matrix_6_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_7_0 = Statvalid ? io_Stationary_matrix_7_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_7_1 = Statvalid ? io_Stationary_matrix_7_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_7_2 = Statvalid ? io_Stationary_matrix_7_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_7_3 = Statvalid ? io_Stationary_matrix_7_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_7_4 = Statvalid ? io_Stationary_matrix_7_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_7_5 = Statvalid ? io_Stationary_matrix_7_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_7_6 = Statvalid ? io_Stationary_matrix_7_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_7_7 = Statvalid ? io_Stationary_matrix_7_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_1_io_Streaming_matrix_0 = _GEN_392[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_1_io_Streaming_matrix_1 = _GEN_393[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_1_io_Streaming_matrix_2 = _GEN_394[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_1_io_Streaming_matrix_3 = _GEN_395[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_1_io_Streaming_matrix_4 = _GEN_396[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_1_io_Streaming_matrix_5 = _GEN_397[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_1_io_Streaming_matrix_6 = _GEN_398[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_1_io_Streaming_matrix_7 = _GEN_399[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_1_io_NoDPE = {{31'd0}, Statvalid}; // @[FlexDPU.scala 77:21]
  assign PathFinder_1_io_DataValid = Statvalid; // @[FlexDPU.scala 98:20 101:25 81:25]
  assign PathFinder_2_clock = clock;
  assign PathFinder_2_reset = reset;
  assign PathFinder_2_io_Stationary_matrix_0_0 = Statvalid ? io_Stationary_matrix_0_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_0_1 = Statvalid ? io_Stationary_matrix_0_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_0_2 = Statvalid ? io_Stationary_matrix_0_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_0_3 = Statvalid ? io_Stationary_matrix_0_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_0_4 = Statvalid ? io_Stationary_matrix_0_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_0_5 = Statvalid ? io_Stationary_matrix_0_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_0_6 = Statvalid ? io_Stationary_matrix_0_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_0_7 = Statvalid ? io_Stationary_matrix_0_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_1_0 = Statvalid ? io_Stationary_matrix_1_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_1_1 = Statvalid ? io_Stationary_matrix_1_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_1_2 = Statvalid ? io_Stationary_matrix_1_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_1_3 = Statvalid ? io_Stationary_matrix_1_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_1_4 = Statvalid ? io_Stationary_matrix_1_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_1_5 = Statvalid ? io_Stationary_matrix_1_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_1_6 = Statvalid ? io_Stationary_matrix_1_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_1_7 = Statvalid ? io_Stationary_matrix_1_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_2_0 = Statvalid ? io_Stationary_matrix_2_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_2_1 = Statvalid ? io_Stationary_matrix_2_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_2_2 = Statvalid ? io_Stationary_matrix_2_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_2_3 = Statvalid ? io_Stationary_matrix_2_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_2_4 = Statvalid ? io_Stationary_matrix_2_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_2_5 = Statvalid ? io_Stationary_matrix_2_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_2_6 = Statvalid ? io_Stationary_matrix_2_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_2_7 = Statvalid ? io_Stationary_matrix_2_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_3_0 = Statvalid ? io_Stationary_matrix_3_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_3_1 = Statvalid ? io_Stationary_matrix_3_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_3_2 = Statvalid ? io_Stationary_matrix_3_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_3_3 = Statvalid ? io_Stationary_matrix_3_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_3_4 = Statvalid ? io_Stationary_matrix_3_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_3_5 = Statvalid ? io_Stationary_matrix_3_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_3_6 = Statvalid ? io_Stationary_matrix_3_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_3_7 = Statvalid ? io_Stationary_matrix_3_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_4_0 = Statvalid ? io_Stationary_matrix_4_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_4_1 = Statvalid ? io_Stationary_matrix_4_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_4_2 = Statvalid ? io_Stationary_matrix_4_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_4_3 = Statvalid ? io_Stationary_matrix_4_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_4_4 = Statvalid ? io_Stationary_matrix_4_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_4_5 = Statvalid ? io_Stationary_matrix_4_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_4_6 = Statvalid ? io_Stationary_matrix_4_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_4_7 = Statvalid ? io_Stationary_matrix_4_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_5_0 = Statvalid ? io_Stationary_matrix_5_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_5_1 = Statvalid ? io_Stationary_matrix_5_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_5_2 = Statvalid ? io_Stationary_matrix_5_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_5_3 = Statvalid ? io_Stationary_matrix_5_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_5_4 = Statvalid ? io_Stationary_matrix_5_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_5_5 = Statvalid ? io_Stationary_matrix_5_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_5_6 = Statvalid ? io_Stationary_matrix_5_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_5_7 = Statvalid ? io_Stationary_matrix_5_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_6_0 = Statvalid ? io_Stationary_matrix_6_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_6_1 = Statvalid ? io_Stationary_matrix_6_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_6_2 = Statvalid ? io_Stationary_matrix_6_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_6_3 = Statvalid ? io_Stationary_matrix_6_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_6_4 = Statvalid ? io_Stationary_matrix_6_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_6_5 = Statvalid ? io_Stationary_matrix_6_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_6_6 = Statvalid ? io_Stationary_matrix_6_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_6_7 = Statvalid ? io_Stationary_matrix_6_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_7_0 = Statvalid ? io_Stationary_matrix_7_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_7_1 = Statvalid ? io_Stationary_matrix_7_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_7_2 = Statvalid ? io_Stationary_matrix_7_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_7_3 = Statvalid ? io_Stationary_matrix_7_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_7_4 = Statvalid ? io_Stationary_matrix_7_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_7_5 = Statvalid ? io_Stationary_matrix_7_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_7_6 = Statvalid ? io_Stationary_matrix_7_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_7_7 = Statvalid ? io_Stationary_matrix_7_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_2_io_Streaming_matrix_0 = _GEN_392[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_2_io_Streaming_matrix_1 = _GEN_393[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_2_io_Streaming_matrix_2 = _GEN_394[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_2_io_Streaming_matrix_3 = _GEN_395[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_2_io_Streaming_matrix_4 = _GEN_396[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_2_io_Streaming_matrix_5 = _GEN_397[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_2_io_Streaming_matrix_6 = _GEN_398[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_2_io_Streaming_matrix_7 = _GEN_399[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_2_io_NoDPE = {{30'd0}, _GEN_729}; // @[FlexDPU.scala 77:21]
  assign PathFinder_2_io_DataValid = Statvalid; // @[FlexDPU.scala 98:20 101:25 81:25]
  assign PathFinder_3_clock = clock;
  assign PathFinder_3_reset = reset;
  assign PathFinder_3_io_Stationary_matrix_0_0 = Statvalid ? io_Stationary_matrix_0_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_0_1 = Statvalid ? io_Stationary_matrix_0_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_0_2 = Statvalid ? io_Stationary_matrix_0_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_0_3 = Statvalid ? io_Stationary_matrix_0_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_0_4 = Statvalid ? io_Stationary_matrix_0_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_0_5 = Statvalid ? io_Stationary_matrix_0_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_0_6 = Statvalid ? io_Stationary_matrix_0_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_0_7 = Statvalid ? io_Stationary_matrix_0_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_1_0 = Statvalid ? io_Stationary_matrix_1_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_1_1 = Statvalid ? io_Stationary_matrix_1_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_1_2 = Statvalid ? io_Stationary_matrix_1_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_1_3 = Statvalid ? io_Stationary_matrix_1_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_1_4 = Statvalid ? io_Stationary_matrix_1_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_1_5 = Statvalid ? io_Stationary_matrix_1_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_1_6 = Statvalid ? io_Stationary_matrix_1_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_1_7 = Statvalid ? io_Stationary_matrix_1_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_2_0 = Statvalid ? io_Stationary_matrix_2_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_2_1 = Statvalid ? io_Stationary_matrix_2_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_2_2 = Statvalid ? io_Stationary_matrix_2_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_2_3 = Statvalid ? io_Stationary_matrix_2_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_2_4 = Statvalid ? io_Stationary_matrix_2_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_2_5 = Statvalid ? io_Stationary_matrix_2_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_2_6 = Statvalid ? io_Stationary_matrix_2_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_2_7 = Statvalid ? io_Stationary_matrix_2_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_3_0 = Statvalid ? io_Stationary_matrix_3_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_3_1 = Statvalid ? io_Stationary_matrix_3_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_3_2 = Statvalid ? io_Stationary_matrix_3_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_3_3 = Statvalid ? io_Stationary_matrix_3_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_3_4 = Statvalid ? io_Stationary_matrix_3_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_3_5 = Statvalid ? io_Stationary_matrix_3_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_3_6 = Statvalid ? io_Stationary_matrix_3_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_3_7 = Statvalid ? io_Stationary_matrix_3_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_4_0 = Statvalid ? io_Stationary_matrix_4_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_4_1 = Statvalid ? io_Stationary_matrix_4_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_4_2 = Statvalid ? io_Stationary_matrix_4_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_4_3 = Statvalid ? io_Stationary_matrix_4_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_4_4 = Statvalid ? io_Stationary_matrix_4_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_4_5 = Statvalid ? io_Stationary_matrix_4_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_4_6 = Statvalid ? io_Stationary_matrix_4_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_4_7 = Statvalid ? io_Stationary_matrix_4_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_5_0 = Statvalid ? io_Stationary_matrix_5_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_5_1 = Statvalid ? io_Stationary_matrix_5_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_5_2 = Statvalid ? io_Stationary_matrix_5_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_5_3 = Statvalid ? io_Stationary_matrix_5_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_5_4 = Statvalid ? io_Stationary_matrix_5_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_5_5 = Statvalid ? io_Stationary_matrix_5_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_5_6 = Statvalid ? io_Stationary_matrix_5_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_5_7 = Statvalid ? io_Stationary_matrix_5_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_6_0 = Statvalid ? io_Stationary_matrix_6_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_6_1 = Statvalid ? io_Stationary_matrix_6_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_6_2 = Statvalid ? io_Stationary_matrix_6_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_6_3 = Statvalid ? io_Stationary_matrix_6_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_6_4 = Statvalid ? io_Stationary_matrix_6_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_6_5 = Statvalid ? io_Stationary_matrix_6_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_6_6 = Statvalid ? io_Stationary_matrix_6_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_6_7 = Statvalid ? io_Stationary_matrix_6_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_7_0 = Statvalid ? io_Stationary_matrix_7_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_7_1 = Statvalid ? io_Stationary_matrix_7_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_7_2 = Statvalid ? io_Stationary_matrix_7_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_7_3 = Statvalid ? io_Stationary_matrix_7_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_7_4 = Statvalid ? io_Stationary_matrix_7_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_7_5 = Statvalid ? io_Stationary_matrix_7_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_7_6 = Statvalid ? io_Stationary_matrix_7_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_7_7 = Statvalid ? io_Stationary_matrix_7_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_3_io_Streaming_matrix_0 = _GEN_392[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_3_io_Streaming_matrix_1 = _GEN_393[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_3_io_Streaming_matrix_2 = _GEN_394[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_3_io_Streaming_matrix_3 = _GEN_395[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_3_io_Streaming_matrix_4 = _GEN_396[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_3_io_Streaming_matrix_5 = _GEN_397[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_3_io_Streaming_matrix_6 = _GEN_398[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_3_io_Streaming_matrix_7 = _GEN_399[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_3_io_NoDPE = {{30'd0}, _GEN_802}; // @[FlexDPU.scala 77:21]
  assign PathFinder_3_io_DataValid = Statvalid; // @[FlexDPU.scala 98:20 101:25 81:25]
  assign PathFinder_4_clock = clock;
  assign PathFinder_4_reset = reset;
  assign PathFinder_4_io_Stationary_matrix_0_0 = Statvalid ? io_Stationary_matrix_0_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_0_1 = Statvalid ? io_Stationary_matrix_0_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_0_2 = Statvalid ? io_Stationary_matrix_0_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_0_3 = Statvalid ? io_Stationary_matrix_0_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_0_4 = Statvalid ? io_Stationary_matrix_0_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_0_5 = Statvalid ? io_Stationary_matrix_0_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_0_6 = Statvalid ? io_Stationary_matrix_0_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_0_7 = Statvalid ? io_Stationary_matrix_0_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_1_0 = Statvalid ? io_Stationary_matrix_1_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_1_1 = Statvalid ? io_Stationary_matrix_1_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_1_2 = Statvalid ? io_Stationary_matrix_1_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_1_3 = Statvalid ? io_Stationary_matrix_1_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_1_4 = Statvalid ? io_Stationary_matrix_1_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_1_5 = Statvalid ? io_Stationary_matrix_1_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_1_6 = Statvalid ? io_Stationary_matrix_1_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_1_7 = Statvalid ? io_Stationary_matrix_1_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_2_0 = Statvalid ? io_Stationary_matrix_2_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_2_1 = Statvalid ? io_Stationary_matrix_2_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_2_2 = Statvalid ? io_Stationary_matrix_2_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_2_3 = Statvalid ? io_Stationary_matrix_2_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_2_4 = Statvalid ? io_Stationary_matrix_2_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_2_5 = Statvalid ? io_Stationary_matrix_2_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_2_6 = Statvalid ? io_Stationary_matrix_2_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_2_7 = Statvalid ? io_Stationary_matrix_2_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_3_0 = Statvalid ? io_Stationary_matrix_3_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_3_1 = Statvalid ? io_Stationary_matrix_3_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_3_2 = Statvalid ? io_Stationary_matrix_3_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_3_3 = Statvalid ? io_Stationary_matrix_3_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_3_4 = Statvalid ? io_Stationary_matrix_3_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_3_5 = Statvalid ? io_Stationary_matrix_3_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_3_6 = Statvalid ? io_Stationary_matrix_3_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_3_7 = Statvalid ? io_Stationary_matrix_3_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_4_0 = Statvalid ? io_Stationary_matrix_4_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_4_1 = Statvalid ? io_Stationary_matrix_4_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_4_2 = Statvalid ? io_Stationary_matrix_4_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_4_3 = Statvalid ? io_Stationary_matrix_4_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_4_4 = Statvalid ? io_Stationary_matrix_4_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_4_5 = Statvalid ? io_Stationary_matrix_4_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_4_6 = Statvalid ? io_Stationary_matrix_4_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_4_7 = Statvalid ? io_Stationary_matrix_4_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_5_0 = Statvalid ? io_Stationary_matrix_5_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_5_1 = Statvalid ? io_Stationary_matrix_5_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_5_2 = Statvalid ? io_Stationary_matrix_5_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_5_3 = Statvalid ? io_Stationary_matrix_5_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_5_4 = Statvalid ? io_Stationary_matrix_5_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_5_5 = Statvalid ? io_Stationary_matrix_5_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_5_6 = Statvalid ? io_Stationary_matrix_5_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_5_7 = Statvalid ? io_Stationary_matrix_5_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_6_0 = Statvalid ? io_Stationary_matrix_6_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_6_1 = Statvalid ? io_Stationary_matrix_6_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_6_2 = Statvalid ? io_Stationary_matrix_6_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_6_3 = Statvalid ? io_Stationary_matrix_6_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_6_4 = Statvalid ? io_Stationary_matrix_6_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_6_5 = Statvalid ? io_Stationary_matrix_6_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_6_6 = Statvalid ? io_Stationary_matrix_6_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_6_7 = Statvalid ? io_Stationary_matrix_6_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_7_0 = Statvalid ? io_Stationary_matrix_7_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_7_1 = Statvalid ? io_Stationary_matrix_7_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_7_2 = Statvalid ? io_Stationary_matrix_7_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_7_3 = Statvalid ? io_Stationary_matrix_7_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_7_4 = Statvalid ? io_Stationary_matrix_7_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_7_5 = Statvalid ? io_Stationary_matrix_7_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_7_6 = Statvalid ? io_Stationary_matrix_7_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_7_7 = Statvalid ? io_Stationary_matrix_7_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_4_io_Streaming_matrix_0 = _GEN_392[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_4_io_Streaming_matrix_1 = _GEN_393[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_4_io_Streaming_matrix_2 = _GEN_394[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_4_io_Streaming_matrix_3 = _GEN_395[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_4_io_Streaming_matrix_4 = _GEN_396[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_4_io_Streaming_matrix_5 = _GEN_397[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_4_io_Streaming_matrix_6 = _GEN_398[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_4_io_Streaming_matrix_7 = _GEN_399[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_4_io_NoDPE = {{29'd0}, _GEN_875}; // @[FlexDPU.scala 77:21]
  assign PathFinder_4_io_DataValid = Statvalid; // @[FlexDPU.scala 98:20 101:25 81:25]
  assign PathFinder_5_clock = clock;
  assign PathFinder_5_reset = reset;
  assign PathFinder_5_io_Stationary_matrix_0_0 = Statvalid ? io_Stationary_matrix_0_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_0_1 = Statvalid ? io_Stationary_matrix_0_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_0_2 = Statvalid ? io_Stationary_matrix_0_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_0_3 = Statvalid ? io_Stationary_matrix_0_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_0_4 = Statvalid ? io_Stationary_matrix_0_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_0_5 = Statvalid ? io_Stationary_matrix_0_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_0_6 = Statvalid ? io_Stationary_matrix_0_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_0_7 = Statvalid ? io_Stationary_matrix_0_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_1_0 = Statvalid ? io_Stationary_matrix_1_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_1_1 = Statvalid ? io_Stationary_matrix_1_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_1_2 = Statvalid ? io_Stationary_matrix_1_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_1_3 = Statvalid ? io_Stationary_matrix_1_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_1_4 = Statvalid ? io_Stationary_matrix_1_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_1_5 = Statvalid ? io_Stationary_matrix_1_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_1_6 = Statvalid ? io_Stationary_matrix_1_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_1_7 = Statvalid ? io_Stationary_matrix_1_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_2_0 = Statvalid ? io_Stationary_matrix_2_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_2_1 = Statvalid ? io_Stationary_matrix_2_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_2_2 = Statvalid ? io_Stationary_matrix_2_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_2_3 = Statvalid ? io_Stationary_matrix_2_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_2_4 = Statvalid ? io_Stationary_matrix_2_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_2_5 = Statvalid ? io_Stationary_matrix_2_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_2_6 = Statvalid ? io_Stationary_matrix_2_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_2_7 = Statvalid ? io_Stationary_matrix_2_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_3_0 = Statvalid ? io_Stationary_matrix_3_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_3_1 = Statvalid ? io_Stationary_matrix_3_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_3_2 = Statvalid ? io_Stationary_matrix_3_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_3_3 = Statvalid ? io_Stationary_matrix_3_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_3_4 = Statvalid ? io_Stationary_matrix_3_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_3_5 = Statvalid ? io_Stationary_matrix_3_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_3_6 = Statvalid ? io_Stationary_matrix_3_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_3_7 = Statvalid ? io_Stationary_matrix_3_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_4_0 = Statvalid ? io_Stationary_matrix_4_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_4_1 = Statvalid ? io_Stationary_matrix_4_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_4_2 = Statvalid ? io_Stationary_matrix_4_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_4_3 = Statvalid ? io_Stationary_matrix_4_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_4_4 = Statvalid ? io_Stationary_matrix_4_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_4_5 = Statvalid ? io_Stationary_matrix_4_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_4_6 = Statvalid ? io_Stationary_matrix_4_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_4_7 = Statvalid ? io_Stationary_matrix_4_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_5_0 = Statvalid ? io_Stationary_matrix_5_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_5_1 = Statvalid ? io_Stationary_matrix_5_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_5_2 = Statvalid ? io_Stationary_matrix_5_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_5_3 = Statvalid ? io_Stationary_matrix_5_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_5_4 = Statvalid ? io_Stationary_matrix_5_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_5_5 = Statvalid ? io_Stationary_matrix_5_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_5_6 = Statvalid ? io_Stationary_matrix_5_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_5_7 = Statvalid ? io_Stationary_matrix_5_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_6_0 = Statvalid ? io_Stationary_matrix_6_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_6_1 = Statvalid ? io_Stationary_matrix_6_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_6_2 = Statvalid ? io_Stationary_matrix_6_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_6_3 = Statvalid ? io_Stationary_matrix_6_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_6_4 = Statvalid ? io_Stationary_matrix_6_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_6_5 = Statvalid ? io_Stationary_matrix_6_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_6_6 = Statvalid ? io_Stationary_matrix_6_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_6_7 = Statvalid ? io_Stationary_matrix_6_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_7_0 = Statvalid ? io_Stationary_matrix_7_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_7_1 = Statvalid ? io_Stationary_matrix_7_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_7_2 = Statvalid ? io_Stationary_matrix_7_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_7_3 = Statvalid ? io_Stationary_matrix_7_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_7_4 = Statvalid ? io_Stationary_matrix_7_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_7_5 = Statvalid ? io_Stationary_matrix_7_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_7_6 = Statvalid ? io_Stationary_matrix_7_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_7_7 = Statvalid ? io_Stationary_matrix_7_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_5_io_Streaming_matrix_0 = _GEN_392[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_5_io_Streaming_matrix_1 = _GEN_393[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_5_io_Streaming_matrix_2 = _GEN_394[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_5_io_Streaming_matrix_3 = _GEN_395[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_5_io_Streaming_matrix_4 = _GEN_396[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_5_io_Streaming_matrix_5 = _GEN_397[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_5_io_Streaming_matrix_6 = _GEN_398[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_5_io_Streaming_matrix_7 = _GEN_399[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_5_io_NoDPE = {{29'd0}, _GEN_948}; // @[FlexDPU.scala 77:21]
  assign PathFinder_5_io_DataValid = Statvalid; // @[FlexDPU.scala 98:20 101:25 81:25]
  assign PathFinder_6_clock = clock;
  assign PathFinder_6_reset = reset;
  assign PathFinder_6_io_Stationary_matrix_0_0 = Statvalid ? io_Stationary_matrix_0_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_0_1 = Statvalid ? io_Stationary_matrix_0_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_0_2 = Statvalid ? io_Stationary_matrix_0_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_0_3 = Statvalid ? io_Stationary_matrix_0_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_0_4 = Statvalid ? io_Stationary_matrix_0_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_0_5 = Statvalid ? io_Stationary_matrix_0_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_0_6 = Statvalid ? io_Stationary_matrix_0_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_0_7 = Statvalid ? io_Stationary_matrix_0_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_1_0 = Statvalid ? io_Stationary_matrix_1_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_1_1 = Statvalid ? io_Stationary_matrix_1_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_1_2 = Statvalid ? io_Stationary_matrix_1_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_1_3 = Statvalid ? io_Stationary_matrix_1_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_1_4 = Statvalid ? io_Stationary_matrix_1_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_1_5 = Statvalid ? io_Stationary_matrix_1_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_1_6 = Statvalid ? io_Stationary_matrix_1_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_1_7 = Statvalid ? io_Stationary_matrix_1_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_2_0 = Statvalid ? io_Stationary_matrix_2_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_2_1 = Statvalid ? io_Stationary_matrix_2_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_2_2 = Statvalid ? io_Stationary_matrix_2_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_2_3 = Statvalid ? io_Stationary_matrix_2_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_2_4 = Statvalid ? io_Stationary_matrix_2_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_2_5 = Statvalid ? io_Stationary_matrix_2_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_2_6 = Statvalid ? io_Stationary_matrix_2_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_2_7 = Statvalid ? io_Stationary_matrix_2_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_3_0 = Statvalid ? io_Stationary_matrix_3_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_3_1 = Statvalid ? io_Stationary_matrix_3_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_3_2 = Statvalid ? io_Stationary_matrix_3_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_3_3 = Statvalid ? io_Stationary_matrix_3_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_3_4 = Statvalid ? io_Stationary_matrix_3_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_3_5 = Statvalid ? io_Stationary_matrix_3_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_3_6 = Statvalid ? io_Stationary_matrix_3_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_3_7 = Statvalid ? io_Stationary_matrix_3_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_4_0 = Statvalid ? io_Stationary_matrix_4_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_4_1 = Statvalid ? io_Stationary_matrix_4_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_4_2 = Statvalid ? io_Stationary_matrix_4_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_4_3 = Statvalid ? io_Stationary_matrix_4_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_4_4 = Statvalid ? io_Stationary_matrix_4_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_4_5 = Statvalid ? io_Stationary_matrix_4_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_4_6 = Statvalid ? io_Stationary_matrix_4_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_4_7 = Statvalid ? io_Stationary_matrix_4_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_5_0 = Statvalid ? io_Stationary_matrix_5_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_5_1 = Statvalid ? io_Stationary_matrix_5_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_5_2 = Statvalid ? io_Stationary_matrix_5_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_5_3 = Statvalid ? io_Stationary_matrix_5_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_5_4 = Statvalid ? io_Stationary_matrix_5_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_5_5 = Statvalid ? io_Stationary_matrix_5_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_5_6 = Statvalid ? io_Stationary_matrix_5_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_5_7 = Statvalid ? io_Stationary_matrix_5_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_6_0 = Statvalid ? io_Stationary_matrix_6_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_6_1 = Statvalid ? io_Stationary_matrix_6_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_6_2 = Statvalid ? io_Stationary_matrix_6_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_6_3 = Statvalid ? io_Stationary_matrix_6_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_6_4 = Statvalid ? io_Stationary_matrix_6_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_6_5 = Statvalid ? io_Stationary_matrix_6_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_6_6 = Statvalid ? io_Stationary_matrix_6_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_6_7 = Statvalid ? io_Stationary_matrix_6_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_7_0 = Statvalid ? io_Stationary_matrix_7_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_7_1 = Statvalid ? io_Stationary_matrix_7_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_7_2 = Statvalid ? io_Stationary_matrix_7_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_7_3 = Statvalid ? io_Stationary_matrix_7_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_7_4 = Statvalid ? io_Stationary_matrix_7_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_7_5 = Statvalid ? io_Stationary_matrix_7_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_7_6 = Statvalid ? io_Stationary_matrix_7_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_7_7 = Statvalid ? io_Stationary_matrix_7_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_6_io_Streaming_matrix_0 = _GEN_392[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_6_io_Streaming_matrix_1 = _GEN_393[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_6_io_Streaming_matrix_2 = _GEN_394[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_6_io_Streaming_matrix_3 = _GEN_395[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_6_io_Streaming_matrix_4 = _GEN_396[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_6_io_Streaming_matrix_5 = _GEN_397[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_6_io_Streaming_matrix_6 = _GEN_398[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_6_io_Streaming_matrix_7 = _GEN_399[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_6_io_NoDPE = {{29'd0}, _GEN_1021}; // @[FlexDPU.scala 77:21]
  assign PathFinder_6_io_DataValid = Statvalid; // @[FlexDPU.scala 98:20 101:25 81:25]
  assign PathFinder_7_clock = clock;
  assign PathFinder_7_reset = reset;
  assign PathFinder_7_io_Stationary_matrix_0_0 = Statvalid ? io_Stationary_matrix_0_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_0_1 = Statvalid ? io_Stationary_matrix_0_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_0_2 = Statvalid ? io_Stationary_matrix_0_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_0_3 = Statvalid ? io_Stationary_matrix_0_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_0_4 = Statvalid ? io_Stationary_matrix_0_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_0_5 = Statvalid ? io_Stationary_matrix_0_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_0_6 = Statvalid ? io_Stationary_matrix_0_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_0_7 = Statvalid ? io_Stationary_matrix_0_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_1_0 = Statvalid ? io_Stationary_matrix_1_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_1_1 = Statvalid ? io_Stationary_matrix_1_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_1_2 = Statvalid ? io_Stationary_matrix_1_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_1_3 = Statvalid ? io_Stationary_matrix_1_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_1_4 = Statvalid ? io_Stationary_matrix_1_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_1_5 = Statvalid ? io_Stationary_matrix_1_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_1_6 = Statvalid ? io_Stationary_matrix_1_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_1_7 = Statvalid ? io_Stationary_matrix_1_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_2_0 = Statvalid ? io_Stationary_matrix_2_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_2_1 = Statvalid ? io_Stationary_matrix_2_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_2_2 = Statvalid ? io_Stationary_matrix_2_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_2_3 = Statvalid ? io_Stationary_matrix_2_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_2_4 = Statvalid ? io_Stationary_matrix_2_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_2_5 = Statvalid ? io_Stationary_matrix_2_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_2_6 = Statvalid ? io_Stationary_matrix_2_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_2_7 = Statvalid ? io_Stationary_matrix_2_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_3_0 = Statvalid ? io_Stationary_matrix_3_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_3_1 = Statvalid ? io_Stationary_matrix_3_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_3_2 = Statvalid ? io_Stationary_matrix_3_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_3_3 = Statvalid ? io_Stationary_matrix_3_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_3_4 = Statvalid ? io_Stationary_matrix_3_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_3_5 = Statvalid ? io_Stationary_matrix_3_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_3_6 = Statvalid ? io_Stationary_matrix_3_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_3_7 = Statvalid ? io_Stationary_matrix_3_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_4_0 = Statvalid ? io_Stationary_matrix_4_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_4_1 = Statvalid ? io_Stationary_matrix_4_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_4_2 = Statvalid ? io_Stationary_matrix_4_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_4_3 = Statvalid ? io_Stationary_matrix_4_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_4_4 = Statvalid ? io_Stationary_matrix_4_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_4_5 = Statvalid ? io_Stationary_matrix_4_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_4_6 = Statvalid ? io_Stationary_matrix_4_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_4_7 = Statvalid ? io_Stationary_matrix_4_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_5_0 = Statvalid ? io_Stationary_matrix_5_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_5_1 = Statvalid ? io_Stationary_matrix_5_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_5_2 = Statvalid ? io_Stationary_matrix_5_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_5_3 = Statvalid ? io_Stationary_matrix_5_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_5_4 = Statvalid ? io_Stationary_matrix_5_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_5_5 = Statvalid ? io_Stationary_matrix_5_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_5_6 = Statvalid ? io_Stationary_matrix_5_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_5_7 = Statvalid ? io_Stationary_matrix_5_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_6_0 = Statvalid ? io_Stationary_matrix_6_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_6_1 = Statvalid ? io_Stationary_matrix_6_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_6_2 = Statvalid ? io_Stationary_matrix_6_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_6_3 = Statvalid ? io_Stationary_matrix_6_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_6_4 = Statvalid ? io_Stationary_matrix_6_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_6_5 = Statvalid ? io_Stationary_matrix_6_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_6_6 = Statvalid ? io_Stationary_matrix_6_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_6_7 = Statvalid ? io_Stationary_matrix_6_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_7_0 = Statvalid ? io_Stationary_matrix_7_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_7_1 = Statvalid ? io_Stationary_matrix_7_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_7_2 = Statvalid ? io_Stationary_matrix_7_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_7_3 = Statvalid ? io_Stationary_matrix_7_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_7_4 = Statvalid ? io_Stationary_matrix_7_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_7_5 = Statvalid ? io_Stationary_matrix_7_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_7_6 = Statvalid ? io_Stationary_matrix_7_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_7_7 = Statvalid ? io_Stationary_matrix_7_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_7_io_Streaming_matrix_0 = _GEN_392[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_7_io_Streaming_matrix_1 = _GEN_393[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_7_io_Streaming_matrix_2 = _GEN_394[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_7_io_Streaming_matrix_3 = _GEN_395[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_7_io_Streaming_matrix_4 = _GEN_396[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_7_io_Streaming_matrix_5 = _GEN_397[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_7_io_Streaming_matrix_6 = _GEN_398[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_7_io_Streaming_matrix_7 = _GEN_399[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_7_io_NoDPE = {{29'd0}, _GEN_1094}; // @[FlexDPU.scala 77:21]
  assign PathFinder_7_io_DataValid = Statvalid; // @[FlexDPU.scala 98:20 101:25 81:25]
  assign PathFinder_8_clock = clock;
  assign PathFinder_8_reset = reset;
  assign PathFinder_8_io_Stationary_matrix_0_0 = Statvalid ? io_Stationary_matrix_0_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_0_1 = Statvalid ? io_Stationary_matrix_0_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_0_2 = Statvalid ? io_Stationary_matrix_0_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_0_3 = Statvalid ? io_Stationary_matrix_0_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_0_4 = Statvalid ? io_Stationary_matrix_0_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_0_5 = Statvalid ? io_Stationary_matrix_0_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_0_6 = Statvalid ? io_Stationary_matrix_0_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_0_7 = Statvalid ? io_Stationary_matrix_0_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_1_0 = Statvalid ? io_Stationary_matrix_1_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_1_1 = Statvalid ? io_Stationary_matrix_1_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_1_2 = Statvalid ? io_Stationary_matrix_1_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_1_3 = Statvalid ? io_Stationary_matrix_1_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_1_4 = Statvalid ? io_Stationary_matrix_1_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_1_5 = Statvalid ? io_Stationary_matrix_1_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_1_6 = Statvalid ? io_Stationary_matrix_1_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_1_7 = Statvalid ? io_Stationary_matrix_1_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_2_0 = Statvalid ? io_Stationary_matrix_2_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_2_1 = Statvalid ? io_Stationary_matrix_2_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_2_2 = Statvalid ? io_Stationary_matrix_2_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_2_3 = Statvalid ? io_Stationary_matrix_2_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_2_4 = Statvalid ? io_Stationary_matrix_2_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_2_5 = Statvalid ? io_Stationary_matrix_2_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_2_6 = Statvalid ? io_Stationary_matrix_2_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_2_7 = Statvalid ? io_Stationary_matrix_2_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_3_0 = Statvalid ? io_Stationary_matrix_3_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_3_1 = Statvalid ? io_Stationary_matrix_3_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_3_2 = Statvalid ? io_Stationary_matrix_3_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_3_3 = Statvalid ? io_Stationary_matrix_3_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_3_4 = Statvalid ? io_Stationary_matrix_3_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_3_5 = Statvalid ? io_Stationary_matrix_3_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_3_6 = Statvalid ? io_Stationary_matrix_3_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_3_7 = Statvalid ? io_Stationary_matrix_3_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_4_0 = Statvalid ? io_Stationary_matrix_4_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_4_1 = Statvalid ? io_Stationary_matrix_4_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_4_2 = Statvalid ? io_Stationary_matrix_4_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_4_3 = Statvalid ? io_Stationary_matrix_4_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_4_4 = Statvalid ? io_Stationary_matrix_4_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_4_5 = Statvalid ? io_Stationary_matrix_4_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_4_6 = Statvalid ? io_Stationary_matrix_4_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_4_7 = Statvalid ? io_Stationary_matrix_4_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_5_0 = Statvalid ? io_Stationary_matrix_5_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_5_1 = Statvalid ? io_Stationary_matrix_5_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_5_2 = Statvalid ? io_Stationary_matrix_5_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_5_3 = Statvalid ? io_Stationary_matrix_5_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_5_4 = Statvalid ? io_Stationary_matrix_5_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_5_5 = Statvalid ? io_Stationary_matrix_5_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_5_6 = Statvalid ? io_Stationary_matrix_5_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_5_7 = Statvalid ? io_Stationary_matrix_5_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_6_0 = Statvalid ? io_Stationary_matrix_6_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_6_1 = Statvalid ? io_Stationary_matrix_6_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_6_2 = Statvalid ? io_Stationary_matrix_6_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_6_3 = Statvalid ? io_Stationary_matrix_6_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_6_4 = Statvalid ? io_Stationary_matrix_6_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_6_5 = Statvalid ? io_Stationary_matrix_6_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_6_6 = Statvalid ? io_Stationary_matrix_6_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_6_7 = Statvalid ? io_Stationary_matrix_6_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_7_0 = Statvalid ? io_Stationary_matrix_7_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_7_1 = Statvalid ? io_Stationary_matrix_7_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_7_2 = Statvalid ? io_Stationary_matrix_7_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_7_3 = Statvalid ? io_Stationary_matrix_7_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_7_4 = Statvalid ? io_Stationary_matrix_7_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_7_5 = Statvalid ? io_Stationary_matrix_7_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_7_6 = Statvalid ? io_Stationary_matrix_7_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_7_7 = Statvalid ? io_Stationary_matrix_7_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_8_io_Streaming_matrix_0 = _GEN_392[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_8_io_Streaming_matrix_1 = _GEN_393[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_8_io_Streaming_matrix_2 = _GEN_394[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_8_io_Streaming_matrix_3 = _GEN_395[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_8_io_Streaming_matrix_4 = _GEN_396[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_8_io_Streaming_matrix_5 = _GEN_397[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_8_io_Streaming_matrix_6 = _GEN_398[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_8_io_Streaming_matrix_7 = _GEN_399[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_8_io_NoDPE = {{28'd0}, _GEN_1167}; // @[FlexDPU.scala 77:21]
  assign PathFinder_8_io_DataValid = Statvalid; // @[FlexDPU.scala 98:20 101:25 81:25]
  assign PathFinder_9_clock = clock;
  assign PathFinder_9_reset = reset;
  assign PathFinder_9_io_Stationary_matrix_0_0 = Statvalid ? io_Stationary_matrix_0_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_0_1 = Statvalid ? io_Stationary_matrix_0_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_0_2 = Statvalid ? io_Stationary_matrix_0_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_0_3 = Statvalid ? io_Stationary_matrix_0_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_0_4 = Statvalid ? io_Stationary_matrix_0_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_0_5 = Statvalid ? io_Stationary_matrix_0_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_0_6 = Statvalid ? io_Stationary_matrix_0_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_0_7 = Statvalid ? io_Stationary_matrix_0_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_1_0 = Statvalid ? io_Stationary_matrix_1_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_1_1 = Statvalid ? io_Stationary_matrix_1_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_1_2 = Statvalid ? io_Stationary_matrix_1_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_1_3 = Statvalid ? io_Stationary_matrix_1_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_1_4 = Statvalid ? io_Stationary_matrix_1_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_1_5 = Statvalid ? io_Stationary_matrix_1_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_1_6 = Statvalid ? io_Stationary_matrix_1_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_1_7 = Statvalid ? io_Stationary_matrix_1_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_2_0 = Statvalid ? io_Stationary_matrix_2_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_2_1 = Statvalid ? io_Stationary_matrix_2_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_2_2 = Statvalid ? io_Stationary_matrix_2_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_2_3 = Statvalid ? io_Stationary_matrix_2_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_2_4 = Statvalid ? io_Stationary_matrix_2_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_2_5 = Statvalid ? io_Stationary_matrix_2_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_2_6 = Statvalid ? io_Stationary_matrix_2_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_2_7 = Statvalid ? io_Stationary_matrix_2_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_3_0 = Statvalid ? io_Stationary_matrix_3_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_3_1 = Statvalid ? io_Stationary_matrix_3_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_3_2 = Statvalid ? io_Stationary_matrix_3_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_3_3 = Statvalid ? io_Stationary_matrix_3_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_3_4 = Statvalid ? io_Stationary_matrix_3_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_3_5 = Statvalid ? io_Stationary_matrix_3_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_3_6 = Statvalid ? io_Stationary_matrix_3_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_3_7 = Statvalid ? io_Stationary_matrix_3_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_4_0 = Statvalid ? io_Stationary_matrix_4_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_4_1 = Statvalid ? io_Stationary_matrix_4_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_4_2 = Statvalid ? io_Stationary_matrix_4_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_4_3 = Statvalid ? io_Stationary_matrix_4_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_4_4 = Statvalid ? io_Stationary_matrix_4_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_4_5 = Statvalid ? io_Stationary_matrix_4_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_4_6 = Statvalid ? io_Stationary_matrix_4_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_4_7 = Statvalid ? io_Stationary_matrix_4_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_5_0 = Statvalid ? io_Stationary_matrix_5_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_5_1 = Statvalid ? io_Stationary_matrix_5_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_5_2 = Statvalid ? io_Stationary_matrix_5_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_5_3 = Statvalid ? io_Stationary_matrix_5_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_5_4 = Statvalid ? io_Stationary_matrix_5_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_5_5 = Statvalid ? io_Stationary_matrix_5_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_5_6 = Statvalid ? io_Stationary_matrix_5_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_5_7 = Statvalid ? io_Stationary_matrix_5_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_6_0 = Statvalid ? io_Stationary_matrix_6_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_6_1 = Statvalid ? io_Stationary_matrix_6_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_6_2 = Statvalid ? io_Stationary_matrix_6_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_6_3 = Statvalid ? io_Stationary_matrix_6_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_6_4 = Statvalid ? io_Stationary_matrix_6_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_6_5 = Statvalid ? io_Stationary_matrix_6_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_6_6 = Statvalid ? io_Stationary_matrix_6_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_6_7 = Statvalid ? io_Stationary_matrix_6_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_7_0 = Statvalid ? io_Stationary_matrix_7_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_7_1 = Statvalid ? io_Stationary_matrix_7_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_7_2 = Statvalid ? io_Stationary_matrix_7_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_7_3 = Statvalid ? io_Stationary_matrix_7_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_7_4 = Statvalid ? io_Stationary_matrix_7_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_7_5 = Statvalid ? io_Stationary_matrix_7_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_7_6 = Statvalid ? io_Stationary_matrix_7_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_7_7 = Statvalid ? io_Stationary_matrix_7_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_9_io_Streaming_matrix_0 = _GEN_392[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_9_io_Streaming_matrix_1 = _GEN_393[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_9_io_Streaming_matrix_2 = _GEN_394[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_9_io_Streaming_matrix_3 = _GEN_395[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_9_io_Streaming_matrix_4 = _GEN_396[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_9_io_Streaming_matrix_5 = _GEN_397[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_9_io_Streaming_matrix_6 = _GEN_398[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_9_io_Streaming_matrix_7 = _GEN_399[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_9_io_NoDPE = {{28'd0}, _GEN_1240}; // @[FlexDPU.scala 77:21]
  assign PathFinder_9_io_DataValid = Statvalid; // @[FlexDPU.scala 98:20 101:25 81:25]
  assign PathFinder_10_clock = clock;
  assign PathFinder_10_reset = reset;
  assign PathFinder_10_io_Stationary_matrix_0_0 = Statvalid ? io_Stationary_matrix_0_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_0_1 = Statvalid ? io_Stationary_matrix_0_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_0_2 = Statvalid ? io_Stationary_matrix_0_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_0_3 = Statvalid ? io_Stationary_matrix_0_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_0_4 = Statvalid ? io_Stationary_matrix_0_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_0_5 = Statvalid ? io_Stationary_matrix_0_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_0_6 = Statvalid ? io_Stationary_matrix_0_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_0_7 = Statvalid ? io_Stationary_matrix_0_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_1_0 = Statvalid ? io_Stationary_matrix_1_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_1_1 = Statvalid ? io_Stationary_matrix_1_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_1_2 = Statvalid ? io_Stationary_matrix_1_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_1_3 = Statvalid ? io_Stationary_matrix_1_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_1_4 = Statvalid ? io_Stationary_matrix_1_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_1_5 = Statvalid ? io_Stationary_matrix_1_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_1_6 = Statvalid ? io_Stationary_matrix_1_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_1_7 = Statvalid ? io_Stationary_matrix_1_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_2_0 = Statvalid ? io_Stationary_matrix_2_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_2_1 = Statvalid ? io_Stationary_matrix_2_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_2_2 = Statvalid ? io_Stationary_matrix_2_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_2_3 = Statvalid ? io_Stationary_matrix_2_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_2_4 = Statvalid ? io_Stationary_matrix_2_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_2_5 = Statvalid ? io_Stationary_matrix_2_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_2_6 = Statvalid ? io_Stationary_matrix_2_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_2_7 = Statvalid ? io_Stationary_matrix_2_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_3_0 = Statvalid ? io_Stationary_matrix_3_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_3_1 = Statvalid ? io_Stationary_matrix_3_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_3_2 = Statvalid ? io_Stationary_matrix_3_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_3_3 = Statvalid ? io_Stationary_matrix_3_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_3_4 = Statvalid ? io_Stationary_matrix_3_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_3_5 = Statvalid ? io_Stationary_matrix_3_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_3_6 = Statvalid ? io_Stationary_matrix_3_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_3_7 = Statvalid ? io_Stationary_matrix_3_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_4_0 = Statvalid ? io_Stationary_matrix_4_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_4_1 = Statvalid ? io_Stationary_matrix_4_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_4_2 = Statvalid ? io_Stationary_matrix_4_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_4_3 = Statvalid ? io_Stationary_matrix_4_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_4_4 = Statvalid ? io_Stationary_matrix_4_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_4_5 = Statvalid ? io_Stationary_matrix_4_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_4_6 = Statvalid ? io_Stationary_matrix_4_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_4_7 = Statvalid ? io_Stationary_matrix_4_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_5_0 = Statvalid ? io_Stationary_matrix_5_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_5_1 = Statvalid ? io_Stationary_matrix_5_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_5_2 = Statvalid ? io_Stationary_matrix_5_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_5_3 = Statvalid ? io_Stationary_matrix_5_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_5_4 = Statvalid ? io_Stationary_matrix_5_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_5_5 = Statvalid ? io_Stationary_matrix_5_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_5_6 = Statvalid ? io_Stationary_matrix_5_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_5_7 = Statvalid ? io_Stationary_matrix_5_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_6_0 = Statvalid ? io_Stationary_matrix_6_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_6_1 = Statvalid ? io_Stationary_matrix_6_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_6_2 = Statvalid ? io_Stationary_matrix_6_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_6_3 = Statvalid ? io_Stationary_matrix_6_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_6_4 = Statvalid ? io_Stationary_matrix_6_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_6_5 = Statvalid ? io_Stationary_matrix_6_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_6_6 = Statvalid ? io_Stationary_matrix_6_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_6_7 = Statvalid ? io_Stationary_matrix_6_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_7_0 = Statvalid ? io_Stationary_matrix_7_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_7_1 = Statvalid ? io_Stationary_matrix_7_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_7_2 = Statvalid ? io_Stationary_matrix_7_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_7_3 = Statvalid ? io_Stationary_matrix_7_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_7_4 = Statvalid ? io_Stationary_matrix_7_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_7_5 = Statvalid ? io_Stationary_matrix_7_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_7_6 = Statvalid ? io_Stationary_matrix_7_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_7_7 = Statvalid ? io_Stationary_matrix_7_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_10_io_Streaming_matrix_0 = _GEN_392[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_10_io_Streaming_matrix_1 = _GEN_393[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_10_io_Streaming_matrix_2 = _GEN_394[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_10_io_Streaming_matrix_3 = _GEN_395[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_10_io_Streaming_matrix_4 = _GEN_396[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_10_io_Streaming_matrix_5 = _GEN_397[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_10_io_Streaming_matrix_6 = _GEN_398[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_10_io_Streaming_matrix_7 = _GEN_399[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_10_io_NoDPE = {{28'd0}, _GEN_1313}; // @[FlexDPU.scala 77:21]
  assign PathFinder_10_io_DataValid = Statvalid; // @[FlexDPU.scala 98:20 101:25 81:25]
  assign PathFinder_11_clock = clock;
  assign PathFinder_11_reset = reset;
  assign PathFinder_11_io_Stationary_matrix_0_0 = Statvalid ? io_Stationary_matrix_0_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_0_1 = Statvalid ? io_Stationary_matrix_0_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_0_2 = Statvalid ? io_Stationary_matrix_0_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_0_3 = Statvalid ? io_Stationary_matrix_0_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_0_4 = Statvalid ? io_Stationary_matrix_0_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_0_5 = Statvalid ? io_Stationary_matrix_0_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_0_6 = Statvalid ? io_Stationary_matrix_0_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_0_7 = Statvalid ? io_Stationary_matrix_0_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_1_0 = Statvalid ? io_Stationary_matrix_1_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_1_1 = Statvalid ? io_Stationary_matrix_1_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_1_2 = Statvalid ? io_Stationary_matrix_1_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_1_3 = Statvalid ? io_Stationary_matrix_1_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_1_4 = Statvalid ? io_Stationary_matrix_1_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_1_5 = Statvalid ? io_Stationary_matrix_1_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_1_6 = Statvalid ? io_Stationary_matrix_1_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_1_7 = Statvalid ? io_Stationary_matrix_1_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_2_0 = Statvalid ? io_Stationary_matrix_2_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_2_1 = Statvalid ? io_Stationary_matrix_2_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_2_2 = Statvalid ? io_Stationary_matrix_2_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_2_3 = Statvalid ? io_Stationary_matrix_2_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_2_4 = Statvalid ? io_Stationary_matrix_2_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_2_5 = Statvalid ? io_Stationary_matrix_2_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_2_6 = Statvalid ? io_Stationary_matrix_2_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_2_7 = Statvalid ? io_Stationary_matrix_2_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_3_0 = Statvalid ? io_Stationary_matrix_3_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_3_1 = Statvalid ? io_Stationary_matrix_3_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_3_2 = Statvalid ? io_Stationary_matrix_3_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_3_3 = Statvalid ? io_Stationary_matrix_3_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_3_4 = Statvalid ? io_Stationary_matrix_3_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_3_5 = Statvalid ? io_Stationary_matrix_3_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_3_6 = Statvalid ? io_Stationary_matrix_3_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_3_7 = Statvalid ? io_Stationary_matrix_3_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_4_0 = Statvalid ? io_Stationary_matrix_4_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_4_1 = Statvalid ? io_Stationary_matrix_4_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_4_2 = Statvalid ? io_Stationary_matrix_4_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_4_3 = Statvalid ? io_Stationary_matrix_4_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_4_4 = Statvalid ? io_Stationary_matrix_4_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_4_5 = Statvalid ? io_Stationary_matrix_4_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_4_6 = Statvalid ? io_Stationary_matrix_4_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_4_7 = Statvalid ? io_Stationary_matrix_4_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_5_0 = Statvalid ? io_Stationary_matrix_5_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_5_1 = Statvalid ? io_Stationary_matrix_5_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_5_2 = Statvalid ? io_Stationary_matrix_5_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_5_3 = Statvalid ? io_Stationary_matrix_5_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_5_4 = Statvalid ? io_Stationary_matrix_5_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_5_5 = Statvalid ? io_Stationary_matrix_5_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_5_6 = Statvalid ? io_Stationary_matrix_5_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_5_7 = Statvalid ? io_Stationary_matrix_5_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_6_0 = Statvalid ? io_Stationary_matrix_6_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_6_1 = Statvalid ? io_Stationary_matrix_6_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_6_2 = Statvalid ? io_Stationary_matrix_6_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_6_3 = Statvalid ? io_Stationary_matrix_6_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_6_4 = Statvalid ? io_Stationary_matrix_6_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_6_5 = Statvalid ? io_Stationary_matrix_6_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_6_6 = Statvalid ? io_Stationary_matrix_6_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_6_7 = Statvalid ? io_Stationary_matrix_6_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_7_0 = Statvalid ? io_Stationary_matrix_7_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_7_1 = Statvalid ? io_Stationary_matrix_7_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_7_2 = Statvalid ? io_Stationary_matrix_7_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_7_3 = Statvalid ? io_Stationary_matrix_7_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_7_4 = Statvalid ? io_Stationary_matrix_7_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_7_5 = Statvalid ? io_Stationary_matrix_7_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_7_6 = Statvalid ? io_Stationary_matrix_7_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_7_7 = Statvalid ? io_Stationary_matrix_7_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_11_io_Streaming_matrix_0 = _GEN_392[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_11_io_Streaming_matrix_1 = _GEN_393[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_11_io_Streaming_matrix_2 = _GEN_394[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_11_io_Streaming_matrix_3 = _GEN_395[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_11_io_Streaming_matrix_4 = _GEN_396[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_11_io_Streaming_matrix_5 = _GEN_397[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_11_io_Streaming_matrix_6 = _GEN_398[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_11_io_Streaming_matrix_7 = _GEN_399[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_11_io_NoDPE = {{28'd0}, _GEN_1386}; // @[FlexDPU.scala 77:21]
  assign PathFinder_11_io_DataValid = Statvalid; // @[FlexDPU.scala 98:20 101:25 81:25]
  assign PathFinder_12_clock = clock;
  assign PathFinder_12_reset = reset;
  assign PathFinder_12_io_Stationary_matrix_0_0 = Statvalid ? io_Stationary_matrix_0_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_0_1 = Statvalid ? io_Stationary_matrix_0_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_0_2 = Statvalid ? io_Stationary_matrix_0_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_0_3 = Statvalid ? io_Stationary_matrix_0_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_0_4 = Statvalid ? io_Stationary_matrix_0_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_0_5 = Statvalid ? io_Stationary_matrix_0_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_0_6 = Statvalid ? io_Stationary_matrix_0_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_0_7 = Statvalid ? io_Stationary_matrix_0_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_1_0 = Statvalid ? io_Stationary_matrix_1_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_1_1 = Statvalid ? io_Stationary_matrix_1_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_1_2 = Statvalid ? io_Stationary_matrix_1_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_1_3 = Statvalid ? io_Stationary_matrix_1_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_1_4 = Statvalid ? io_Stationary_matrix_1_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_1_5 = Statvalid ? io_Stationary_matrix_1_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_1_6 = Statvalid ? io_Stationary_matrix_1_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_1_7 = Statvalid ? io_Stationary_matrix_1_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_2_0 = Statvalid ? io_Stationary_matrix_2_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_2_1 = Statvalid ? io_Stationary_matrix_2_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_2_2 = Statvalid ? io_Stationary_matrix_2_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_2_3 = Statvalid ? io_Stationary_matrix_2_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_2_4 = Statvalid ? io_Stationary_matrix_2_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_2_5 = Statvalid ? io_Stationary_matrix_2_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_2_6 = Statvalid ? io_Stationary_matrix_2_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_2_7 = Statvalid ? io_Stationary_matrix_2_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_3_0 = Statvalid ? io_Stationary_matrix_3_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_3_1 = Statvalid ? io_Stationary_matrix_3_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_3_2 = Statvalid ? io_Stationary_matrix_3_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_3_3 = Statvalid ? io_Stationary_matrix_3_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_3_4 = Statvalid ? io_Stationary_matrix_3_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_3_5 = Statvalid ? io_Stationary_matrix_3_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_3_6 = Statvalid ? io_Stationary_matrix_3_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_3_7 = Statvalid ? io_Stationary_matrix_3_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_4_0 = Statvalid ? io_Stationary_matrix_4_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_4_1 = Statvalid ? io_Stationary_matrix_4_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_4_2 = Statvalid ? io_Stationary_matrix_4_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_4_3 = Statvalid ? io_Stationary_matrix_4_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_4_4 = Statvalid ? io_Stationary_matrix_4_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_4_5 = Statvalid ? io_Stationary_matrix_4_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_4_6 = Statvalid ? io_Stationary_matrix_4_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_4_7 = Statvalid ? io_Stationary_matrix_4_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_5_0 = Statvalid ? io_Stationary_matrix_5_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_5_1 = Statvalid ? io_Stationary_matrix_5_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_5_2 = Statvalid ? io_Stationary_matrix_5_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_5_3 = Statvalid ? io_Stationary_matrix_5_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_5_4 = Statvalid ? io_Stationary_matrix_5_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_5_5 = Statvalid ? io_Stationary_matrix_5_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_5_6 = Statvalid ? io_Stationary_matrix_5_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_5_7 = Statvalid ? io_Stationary_matrix_5_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_6_0 = Statvalid ? io_Stationary_matrix_6_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_6_1 = Statvalid ? io_Stationary_matrix_6_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_6_2 = Statvalid ? io_Stationary_matrix_6_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_6_3 = Statvalid ? io_Stationary_matrix_6_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_6_4 = Statvalid ? io_Stationary_matrix_6_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_6_5 = Statvalid ? io_Stationary_matrix_6_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_6_6 = Statvalid ? io_Stationary_matrix_6_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_6_7 = Statvalid ? io_Stationary_matrix_6_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_7_0 = Statvalid ? io_Stationary_matrix_7_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_7_1 = Statvalid ? io_Stationary_matrix_7_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_7_2 = Statvalid ? io_Stationary_matrix_7_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_7_3 = Statvalid ? io_Stationary_matrix_7_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_7_4 = Statvalid ? io_Stationary_matrix_7_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_7_5 = Statvalid ? io_Stationary_matrix_7_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_7_6 = Statvalid ? io_Stationary_matrix_7_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_7_7 = Statvalid ? io_Stationary_matrix_7_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_12_io_Streaming_matrix_0 = _GEN_392[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_12_io_Streaming_matrix_1 = _GEN_393[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_12_io_Streaming_matrix_2 = _GEN_394[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_12_io_Streaming_matrix_3 = _GEN_395[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_12_io_Streaming_matrix_4 = _GEN_396[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_12_io_Streaming_matrix_5 = _GEN_397[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_12_io_Streaming_matrix_6 = _GEN_398[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_12_io_Streaming_matrix_7 = _GEN_399[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_12_io_NoDPE = {{28'd0}, _GEN_1459}; // @[FlexDPU.scala 77:21]
  assign PathFinder_12_io_DataValid = Statvalid; // @[FlexDPU.scala 98:20 101:25 81:25]
  assign PathFinder_13_clock = clock;
  assign PathFinder_13_reset = reset;
  assign PathFinder_13_io_Stationary_matrix_0_0 = Statvalid ? io_Stationary_matrix_0_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_0_1 = Statvalid ? io_Stationary_matrix_0_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_0_2 = Statvalid ? io_Stationary_matrix_0_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_0_3 = Statvalid ? io_Stationary_matrix_0_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_0_4 = Statvalid ? io_Stationary_matrix_0_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_0_5 = Statvalid ? io_Stationary_matrix_0_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_0_6 = Statvalid ? io_Stationary_matrix_0_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_0_7 = Statvalid ? io_Stationary_matrix_0_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_1_0 = Statvalid ? io_Stationary_matrix_1_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_1_1 = Statvalid ? io_Stationary_matrix_1_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_1_2 = Statvalid ? io_Stationary_matrix_1_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_1_3 = Statvalid ? io_Stationary_matrix_1_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_1_4 = Statvalid ? io_Stationary_matrix_1_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_1_5 = Statvalid ? io_Stationary_matrix_1_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_1_6 = Statvalid ? io_Stationary_matrix_1_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_1_7 = Statvalid ? io_Stationary_matrix_1_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_2_0 = Statvalid ? io_Stationary_matrix_2_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_2_1 = Statvalid ? io_Stationary_matrix_2_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_2_2 = Statvalid ? io_Stationary_matrix_2_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_2_3 = Statvalid ? io_Stationary_matrix_2_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_2_4 = Statvalid ? io_Stationary_matrix_2_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_2_5 = Statvalid ? io_Stationary_matrix_2_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_2_6 = Statvalid ? io_Stationary_matrix_2_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_2_7 = Statvalid ? io_Stationary_matrix_2_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_3_0 = Statvalid ? io_Stationary_matrix_3_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_3_1 = Statvalid ? io_Stationary_matrix_3_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_3_2 = Statvalid ? io_Stationary_matrix_3_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_3_3 = Statvalid ? io_Stationary_matrix_3_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_3_4 = Statvalid ? io_Stationary_matrix_3_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_3_5 = Statvalid ? io_Stationary_matrix_3_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_3_6 = Statvalid ? io_Stationary_matrix_3_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_3_7 = Statvalid ? io_Stationary_matrix_3_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_4_0 = Statvalid ? io_Stationary_matrix_4_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_4_1 = Statvalid ? io_Stationary_matrix_4_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_4_2 = Statvalid ? io_Stationary_matrix_4_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_4_3 = Statvalid ? io_Stationary_matrix_4_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_4_4 = Statvalid ? io_Stationary_matrix_4_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_4_5 = Statvalid ? io_Stationary_matrix_4_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_4_6 = Statvalid ? io_Stationary_matrix_4_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_4_7 = Statvalid ? io_Stationary_matrix_4_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_5_0 = Statvalid ? io_Stationary_matrix_5_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_5_1 = Statvalid ? io_Stationary_matrix_5_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_5_2 = Statvalid ? io_Stationary_matrix_5_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_5_3 = Statvalid ? io_Stationary_matrix_5_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_5_4 = Statvalid ? io_Stationary_matrix_5_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_5_5 = Statvalid ? io_Stationary_matrix_5_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_5_6 = Statvalid ? io_Stationary_matrix_5_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_5_7 = Statvalid ? io_Stationary_matrix_5_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_6_0 = Statvalid ? io_Stationary_matrix_6_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_6_1 = Statvalid ? io_Stationary_matrix_6_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_6_2 = Statvalid ? io_Stationary_matrix_6_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_6_3 = Statvalid ? io_Stationary_matrix_6_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_6_4 = Statvalid ? io_Stationary_matrix_6_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_6_5 = Statvalid ? io_Stationary_matrix_6_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_6_6 = Statvalid ? io_Stationary_matrix_6_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_6_7 = Statvalid ? io_Stationary_matrix_6_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_7_0 = Statvalid ? io_Stationary_matrix_7_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_7_1 = Statvalid ? io_Stationary_matrix_7_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_7_2 = Statvalid ? io_Stationary_matrix_7_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_7_3 = Statvalid ? io_Stationary_matrix_7_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_7_4 = Statvalid ? io_Stationary_matrix_7_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_7_5 = Statvalid ? io_Stationary_matrix_7_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_7_6 = Statvalid ? io_Stationary_matrix_7_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_7_7 = Statvalid ? io_Stationary_matrix_7_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_13_io_Streaming_matrix_0 = _GEN_392[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_13_io_Streaming_matrix_1 = _GEN_393[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_13_io_Streaming_matrix_2 = _GEN_394[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_13_io_Streaming_matrix_3 = _GEN_395[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_13_io_Streaming_matrix_4 = _GEN_396[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_13_io_Streaming_matrix_5 = _GEN_397[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_13_io_Streaming_matrix_6 = _GEN_398[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_13_io_Streaming_matrix_7 = _GEN_399[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_13_io_NoDPE = {{28'd0}, _GEN_1532}; // @[FlexDPU.scala 77:21]
  assign PathFinder_13_io_DataValid = Statvalid; // @[FlexDPU.scala 98:20 101:25 81:25]
  assign PathFinder_14_clock = clock;
  assign PathFinder_14_reset = reset;
  assign PathFinder_14_io_Stationary_matrix_0_0 = Statvalid ? io_Stationary_matrix_0_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_0_1 = Statvalid ? io_Stationary_matrix_0_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_0_2 = Statvalid ? io_Stationary_matrix_0_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_0_3 = Statvalid ? io_Stationary_matrix_0_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_0_4 = Statvalid ? io_Stationary_matrix_0_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_0_5 = Statvalid ? io_Stationary_matrix_0_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_0_6 = Statvalid ? io_Stationary_matrix_0_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_0_7 = Statvalid ? io_Stationary_matrix_0_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_1_0 = Statvalid ? io_Stationary_matrix_1_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_1_1 = Statvalid ? io_Stationary_matrix_1_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_1_2 = Statvalid ? io_Stationary_matrix_1_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_1_3 = Statvalid ? io_Stationary_matrix_1_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_1_4 = Statvalid ? io_Stationary_matrix_1_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_1_5 = Statvalid ? io_Stationary_matrix_1_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_1_6 = Statvalid ? io_Stationary_matrix_1_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_1_7 = Statvalid ? io_Stationary_matrix_1_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_2_0 = Statvalid ? io_Stationary_matrix_2_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_2_1 = Statvalid ? io_Stationary_matrix_2_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_2_2 = Statvalid ? io_Stationary_matrix_2_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_2_3 = Statvalid ? io_Stationary_matrix_2_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_2_4 = Statvalid ? io_Stationary_matrix_2_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_2_5 = Statvalid ? io_Stationary_matrix_2_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_2_6 = Statvalid ? io_Stationary_matrix_2_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_2_7 = Statvalid ? io_Stationary_matrix_2_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_3_0 = Statvalid ? io_Stationary_matrix_3_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_3_1 = Statvalid ? io_Stationary_matrix_3_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_3_2 = Statvalid ? io_Stationary_matrix_3_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_3_3 = Statvalid ? io_Stationary_matrix_3_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_3_4 = Statvalid ? io_Stationary_matrix_3_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_3_5 = Statvalid ? io_Stationary_matrix_3_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_3_6 = Statvalid ? io_Stationary_matrix_3_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_3_7 = Statvalid ? io_Stationary_matrix_3_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_4_0 = Statvalid ? io_Stationary_matrix_4_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_4_1 = Statvalid ? io_Stationary_matrix_4_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_4_2 = Statvalid ? io_Stationary_matrix_4_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_4_3 = Statvalid ? io_Stationary_matrix_4_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_4_4 = Statvalid ? io_Stationary_matrix_4_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_4_5 = Statvalid ? io_Stationary_matrix_4_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_4_6 = Statvalid ? io_Stationary_matrix_4_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_4_7 = Statvalid ? io_Stationary_matrix_4_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_5_0 = Statvalid ? io_Stationary_matrix_5_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_5_1 = Statvalid ? io_Stationary_matrix_5_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_5_2 = Statvalid ? io_Stationary_matrix_5_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_5_3 = Statvalid ? io_Stationary_matrix_5_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_5_4 = Statvalid ? io_Stationary_matrix_5_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_5_5 = Statvalid ? io_Stationary_matrix_5_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_5_6 = Statvalid ? io_Stationary_matrix_5_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_5_7 = Statvalid ? io_Stationary_matrix_5_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_6_0 = Statvalid ? io_Stationary_matrix_6_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_6_1 = Statvalid ? io_Stationary_matrix_6_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_6_2 = Statvalid ? io_Stationary_matrix_6_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_6_3 = Statvalid ? io_Stationary_matrix_6_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_6_4 = Statvalid ? io_Stationary_matrix_6_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_6_5 = Statvalid ? io_Stationary_matrix_6_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_6_6 = Statvalid ? io_Stationary_matrix_6_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_6_7 = Statvalid ? io_Stationary_matrix_6_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_7_0 = Statvalid ? io_Stationary_matrix_7_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_7_1 = Statvalid ? io_Stationary_matrix_7_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_7_2 = Statvalid ? io_Stationary_matrix_7_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_7_3 = Statvalid ? io_Stationary_matrix_7_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_7_4 = Statvalid ? io_Stationary_matrix_7_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_7_5 = Statvalid ? io_Stationary_matrix_7_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_7_6 = Statvalid ? io_Stationary_matrix_7_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_7_7 = Statvalid ? io_Stationary_matrix_7_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_14_io_Streaming_matrix_0 = _GEN_392[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_14_io_Streaming_matrix_1 = _GEN_393[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_14_io_Streaming_matrix_2 = _GEN_394[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_14_io_Streaming_matrix_3 = _GEN_395[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_14_io_Streaming_matrix_4 = _GEN_396[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_14_io_Streaming_matrix_5 = _GEN_397[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_14_io_Streaming_matrix_6 = _GEN_398[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_14_io_Streaming_matrix_7 = _GEN_399[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_14_io_NoDPE = {{28'd0}, _GEN_1605}; // @[FlexDPU.scala 77:21]
  assign PathFinder_14_io_DataValid = Statvalid; // @[FlexDPU.scala 98:20 101:25 81:25]
  assign PathFinder_15_clock = clock;
  assign PathFinder_15_reset = reset;
  assign PathFinder_15_io_Stationary_matrix_0_0 = Statvalid ? io_Stationary_matrix_0_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_0_1 = Statvalid ? io_Stationary_matrix_0_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_0_2 = Statvalid ? io_Stationary_matrix_0_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_0_3 = Statvalid ? io_Stationary_matrix_0_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_0_4 = Statvalid ? io_Stationary_matrix_0_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_0_5 = Statvalid ? io_Stationary_matrix_0_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_0_6 = Statvalid ? io_Stationary_matrix_0_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_0_7 = Statvalid ? io_Stationary_matrix_0_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_1_0 = Statvalid ? io_Stationary_matrix_1_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_1_1 = Statvalid ? io_Stationary_matrix_1_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_1_2 = Statvalid ? io_Stationary_matrix_1_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_1_3 = Statvalid ? io_Stationary_matrix_1_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_1_4 = Statvalid ? io_Stationary_matrix_1_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_1_5 = Statvalid ? io_Stationary_matrix_1_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_1_6 = Statvalid ? io_Stationary_matrix_1_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_1_7 = Statvalid ? io_Stationary_matrix_1_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_2_0 = Statvalid ? io_Stationary_matrix_2_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_2_1 = Statvalid ? io_Stationary_matrix_2_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_2_2 = Statvalid ? io_Stationary_matrix_2_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_2_3 = Statvalid ? io_Stationary_matrix_2_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_2_4 = Statvalid ? io_Stationary_matrix_2_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_2_5 = Statvalid ? io_Stationary_matrix_2_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_2_6 = Statvalid ? io_Stationary_matrix_2_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_2_7 = Statvalid ? io_Stationary_matrix_2_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_3_0 = Statvalid ? io_Stationary_matrix_3_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_3_1 = Statvalid ? io_Stationary_matrix_3_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_3_2 = Statvalid ? io_Stationary_matrix_3_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_3_3 = Statvalid ? io_Stationary_matrix_3_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_3_4 = Statvalid ? io_Stationary_matrix_3_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_3_5 = Statvalid ? io_Stationary_matrix_3_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_3_6 = Statvalid ? io_Stationary_matrix_3_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_3_7 = Statvalid ? io_Stationary_matrix_3_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_4_0 = Statvalid ? io_Stationary_matrix_4_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_4_1 = Statvalid ? io_Stationary_matrix_4_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_4_2 = Statvalid ? io_Stationary_matrix_4_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_4_3 = Statvalid ? io_Stationary_matrix_4_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_4_4 = Statvalid ? io_Stationary_matrix_4_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_4_5 = Statvalid ? io_Stationary_matrix_4_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_4_6 = Statvalid ? io_Stationary_matrix_4_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_4_7 = Statvalid ? io_Stationary_matrix_4_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_5_0 = Statvalid ? io_Stationary_matrix_5_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_5_1 = Statvalid ? io_Stationary_matrix_5_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_5_2 = Statvalid ? io_Stationary_matrix_5_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_5_3 = Statvalid ? io_Stationary_matrix_5_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_5_4 = Statvalid ? io_Stationary_matrix_5_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_5_5 = Statvalid ? io_Stationary_matrix_5_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_5_6 = Statvalid ? io_Stationary_matrix_5_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_5_7 = Statvalid ? io_Stationary_matrix_5_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_6_0 = Statvalid ? io_Stationary_matrix_6_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_6_1 = Statvalid ? io_Stationary_matrix_6_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_6_2 = Statvalid ? io_Stationary_matrix_6_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_6_3 = Statvalid ? io_Stationary_matrix_6_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_6_4 = Statvalid ? io_Stationary_matrix_6_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_6_5 = Statvalid ? io_Stationary_matrix_6_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_6_6 = Statvalid ? io_Stationary_matrix_6_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_6_7 = Statvalid ? io_Stationary_matrix_6_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_7_0 = Statvalid ? io_Stationary_matrix_7_0 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_7_1 = Statvalid ? io_Stationary_matrix_7_1 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_7_2 = Statvalid ? io_Stationary_matrix_7_2 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_7_3 = Statvalid ? io_Stationary_matrix_7_3 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_7_4 = Statvalid ? io_Stationary_matrix_7_4 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_7_5 = Statvalid ? io_Stationary_matrix_7_5 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_7_6 = Statvalid ? io_Stationary_matrix_7_6 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_7_7 = Statvalid ? io_Stationary_matrix_7_7 : 16'h0; // @[FlexDPU.scala 98:20 102:33 82:33]
  assign PathFinder_15_io_Streaming_matrix_0 = _GEN_392[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_15_io_Streaming_matrix_1 = _GEN_393[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_15_io_Streaming_matrix_2 = _GEN_394[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_15_io_Streaming_matrix_3 = _GEN_395[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_15_io_Streaming_matrix_4 = _GEN_396[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_15_io_Streaming_matrix_5 = _GEN_397[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_15_io_Streaming_matrix_6 = _GEN_398[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_15_io_Streaming_matrix_7 = _GEN_399[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_15_io_NoDPE = {{28'd0}, _GEN_1678}; // @[FlexDPU.scala 77:21]
  assign PathFinder_15_io_DataValid = Statvalid; // @[FlexDPU.scala 98:20 101:25 81:25]
  assign flexdpecom4_clock = clock;
  assign flexdpecom4_reset = reset;
  assign flexdpecom4_io_i_data_valid = 1'h1; // @[FlexDPU.scala 110:27 114:34]
  assign flexdpecom4_io_i_data_bus_0 = PathFinder_io_Source_0; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_io_i_data_bus_1 = PathFinder_io_Source_1; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_io_i_data_bus_2 = PathFinder_io_Source_2; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_io_i_data_bus_3 = PathFinder_io_Source_3; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_io_i_data_bus2_0 = PathFinder_io_destination_0; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_io_i_data_bus2_1 = PathFinder_io_destination_1; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_io_i_data_bus2_2 = PathFinder_io_destination_2; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_io_i_data_bus2_3 = PathFinder_io_destination_3; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_io_i_mux_bus_0 = PathFinder_io_i_mux_bus_0; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_io_i_mux_bus_1 = PathFinder_io_i_mux_bus_1; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_io_i_mux_bus_2 = PathFinder_io_i_mux_bus_2; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_io_i_mux_bus_3 = PathFinder_io_i_mux_bus_3; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_1_clock = clock;
  assign flexdpecom4_1_reset = reset;
  assign flexdpecom4_1_io_i_data_valid = 1'h1; // @[FlexDPU.scala 110:27 114:34]
  assign flexdpecom4_1_io_i_data_bus_0 = PathFinder_1_io_Source_0; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_1_io_i_data_bus_1 = PathFinder_1_io_Source_1; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_1_io_i_data_bus_2 = PathFinder_1_io_Source_2; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_1_io_i_data_bus_3 = PathFinder_1_io_Source_3; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_1_io_i_data_bus2_0 = PathFinder_1_io_destination_0; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_1_io_i_data_bus2_1 = PathFinder_1_io_destination_1; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_1_io_i_data_bus2_2 = PathFinder_1_io_destination_2; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_1_io_i_data_bus2_3 = PathFinder_1_io_destination_3; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_1_io_i_mux_bus_0 = PathFinder_1_io_i_mux_bus_0; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_1_io_i_mux_bus_1 = PathFinder_1_io_i_mux_bus_1; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_1_io_i_mux_bus_2 = PathFinder_1_io_i_mux_bus_2; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_1_io_i_mux_bus_3 = PathFinder_1_io_i_mux_bus_3; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_2_clock = clock;
  assign flexdpecom4_2_reset = reset;
  assign flexdpecom4_2_io_i_data_valid = 1'h1; // @[FlexDPU.scala 110:27 114:34]
  assign flexdpecom4_2_io_i_data_bus_0 = PathFinder_2_io_Source_0; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_2_io_i_data_bus_1 = PathFinder_2_io_Source_1; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_2_io_i_data_bus_2 = PathFinder_2_io_Source_2; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_2_io_i_data_bus_3 = PathFinder_2_io_Source_3; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_2_io_i_data_bus2_0 = PathFinder_2_io_destination_0; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_2_io_i_data_bus2_1 = PathFinder_2_io_destination_1; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_2_io_i_data_bus2_2 = PathFinder_2_io_destination_2; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_2_io_i_data_bus2_3 = PathFinder_2_io_destination_3; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_2_io_i_mux_bus_0 = PathFinder_2_io_i_mux_bus_0; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_2_io_i_mux_bus_1 = PathFinder_2_io_i_mux_bus_1; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_2_io_i_mux_bus_2 = PathFinder_2_io_i_mux_bus_2; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_2_io_i_mux_bus_3 = PathFinder_2_io_i_mux_bus_3; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_3_clock = clock;
  assign flexdpecom4_3_reset = reset;
  assign flexdpecom4_3_io_i_data_valid = 1'h1; // @[FlexDPU.scala 110:27 114:34]
  assign flexdpecom4_3_io_i_data_bus_0 = PathFinder_3_io_Source_0; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_3_io_i_data_bus_1 = PathFinder_3_io_Source_1; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_3_io_i_data_bus_2 = PathFinder_3_io_Source_2; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_3_io_i_data_bus_3 = PathFinder_3_io_Source_3; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_3_io_i_data_bus2_0 = PathFinder_3_io_destination_0; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_3_io_i_data_bus2_1 = PathFinder_3_io_destination_1; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_3_io_i_data_bus2_2 = PathFinder_3_io_destination_2; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_3_io_i_data_bus2_3 = PathFinder_3_io_destination_3; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_3_io_i_mux_bus_0 = PathFinder_3_io_i_mux_bus_0; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_3_io_i_mux_bus_1 = PathFinder_3_io_i_mux_bus_1; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_3_io_i_mux_bus_2 = PathFinder_3_io_i_mux_bus_2; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_3_io_i_mux_bus_3 = PathFinder_3_io_i_mux_bus_3; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_4_clock = clock;
  assign flexdpecom4_4_reset = reset;
  assign flexdpecom4_4_io_i_data_valid = 1'h1; // @[FlexDPU.scala 110:27 114:34]
  assign flexdpecom4_4_io_i_data_bus_0 = PathFinder_4_io_Source_0; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_4_io_i_data_bus_1 = PathFinder_4_io_Source_1; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_4_io_i_data_bus_2 = PathFinder_4_io_Source_2; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_4_io_i_data_bus_3 = PathFinder_4_io_Source_3; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_4_io_i_data_bus2_0 = PathFinder_4_io_destination_0; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_4_io_i_data_bus2_1 = PathFinder_4_io_destination_1; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_4_io_i_data_bus2_2 = PathFinder_4_io_destination_2; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_4_io_i_data_bus2_3 = PathFinder_4_io_destination_3; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_4_io_i_mux_bus_0 = PathFinder_4_io_i_mux_bus_0; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_4_io_i_mux_bus_1 = PathFinder_4_io_i_mux_bus_1; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_4_io_i_mux_bus_2 = PathFinder_4_io_i_mux_bus_2; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_4_io_i_mux_bus_3 = PathFinder_4_io_i_mux_bus_3; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_5_clock = clock;
  assign flexdpecom4_5_reset = reset;
  assign flexdpecom4_5_io_i_data_valid = 1'h1; // @[FlexDPU.scala 110:27 114:34]
  assign flexdpecom4_5_io_i_data_bus_0 = PathFinder_5_io_Source_0; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_5_io_i_data_bus_1 = PathFinder_5_io_Source_1; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_5_io_i_data_bus_2 = PathFinder_5_io_Source_2; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_5_io_i_data_bus_3 = PathFinder_5_io_Source_3; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_5_io_i_data_bus2_0 = PathFinder_5_io_destination_0; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_5_io_i_data_bus2_1 = PathFinder_5_io_destination_1; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_5_io_i_data_bus2_2 = PathFinder_5_io_destination_2; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_5_io_i_data_bus2_3 = PathFinder_5_io_destination_3; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_5_io_i_mux_bus_0 = PathFinder_5_io_i_mux_bus_0; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_5_io_i_mux_bus_1 = PathFinder_5_io_i_mux_bus_1; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_5_io_i_mux_bus_2 = PathFinder_5_io_i_mux_bus_2; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_5_io_i_mux_bus_3 = PathFinder_5_io_i_mux_bus_3; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_6_clock = clock;
  assign flexdpecom4_6_reset = reset;
  assign flexdpecom4_6_io_i_data_valid = 1'h1; // @[FlexDPU.scala 110:27 114:34]
  assign flexdpecom4_6_io_i_data_bus_0 = PathFinder_6_io_Source_0; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_6_io_i_data_bus_1 = PathFinder_6_io_Source_1; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_6_io_i_data_bus_2 = PathFinder_6_io_Source_2; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_6_io_i_data_bus_3 = PathFinder_6_io_Source_3; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_6_io_i_data_bus2_0 = PathFinder_6_io_destination_0; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_6_io_i_data_bus2_1 = PathFinder_6_io_destination_1; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_6_io_i_data_bus2_2 = PathFinder_6_io_destination_2; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_6_io_i_data_bus2_3 = PathFinder_6_io_destination_3; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_6_io_i_mux_bus_0 = PathFinder_6_io_i_mux_bus_0; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_6_io_i_mux_bus_1 = PathFinder_6_io_i_mux_bus_1; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_6_io_i_mux_bus_2 = PathFinder_6_io_i_mux_bus_2; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_6_io_i_mux_bus_3 = PathFinder_6_io_i_mux_bus_3; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_7_clock = clock;
  assign flexdpecom4_7_reset = reset;
  assign flexdpecom4_7_io_i_data_valid = 1'h1; // @[FlexDPU.scala 110:27 114:34]
  assign flexdpecom4_7_io_i_data_bus_0 = PathFinder_7_io_Source_0; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_7_io_i_data_bus_1 = PathFinder_7_io_Source_1; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_7_io_i_data_bus_2 = PathFinder_7_io_Source_2; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_7_io_i_data_bus_3 = PathFinder_7_io_Source_3; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_7_io_i_data_bus2_0 = PathFinder_7_io_destination_0; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_7_io_i_data_bus2_1 = PathFinder_7_io_destination_1; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_7_io_i_data_bus2_2 = PathFinder_7_io_destination_2; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_7_io_i_data_bus2_3 = PathFinder_7_io_destination_3; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_7_io_i_mux_bus_0 = PathFinder_7_io_i_mux_bus_0; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_7_io_i_mux_bus_1 = PathFinder_7_io_i_mux_bus_1; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_7_io_i_mux_bus_2 = PathFinder_7_io_i_mux_bus_2; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_7_io_i_mux_bus_3 = PathFinder_7_io_i_mux_bus_3; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_8_clock = clock;
  assign flexdpecom4_8_reset = reset;
  assign flexdpecom4_8_io_i_data_valid = 1'h1; // @[FlexDPU.scala 110:27 114:34]
  assign flexdpecom4_8_io_i_data_bus_0 = PathFinder_8_io_Source_0; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_8_io_i_data_bus_1 = PathFinder_8_io_Source_1; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_8_io_i_data_bus_2 = PathFinder_8_io_Source_2; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_8_io_i_data_bus_3 = PathFinder_8_io_Source_3; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_8_io_i_data_bus2_0 = PathFinder_8_io_destination_0; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_8_io_i_data_bus2_1 = PathFinder_8_io_destination_1; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_8_io_i_data_bus2_2 = PathFinder_8_io_destination_2; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_8_io_i_data_bus2_3 = PathFinder_8_io_destination_3; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_8_io_i_mux_bus_0 = PathFinder_8_io_i_mux_bus_0; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_8_io_i_mux_bus_1 = PathFinder_8_io_i_mux_bus_1; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_8_io_i_mux_bus_2 = PathFinder_8_io_i_mux_bus_2; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_8_io_i_mux_bus_3 = PathFinder_8_io_i_mux_bus_3; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_9_clock = clock;
  assign flexdpecom4_9_reset = reset;
  assign flexdpecom4_9_io_i_data_valid = 1'h1; // @[FlexDPU.scala 110:27 114:34]
  assign flexdpecom4_9_io_i_data_bus_0 = PathFinder_9_io_Source_0; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_9_io_i_data_bus_1 = PathFinder_9_io_Source_1; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_9_io_i_data_bus_2 = PathFinder_9_io_Source_2; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_9_io_i_data_bus_3 = PathFinder_9_io_Source_3; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_9_io_i_data_bus2_0 = PathFinder_9_io_destination_0; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_9_io_i_data_bus2_1 = PathFinder_9_io_destination_1; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_9_io_i_data_bus2_2 = PathFinder_9_io_destination_2; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_9_io_i_data_bus2_3 = PathFinder_9_io_destination_3; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_9_io_i_mux_bus_0 = PathFinder_9_io_i_mux_bus_0; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_9_io_i_mux_bus_1 = PathFinder_9_io_i_mux_bus_1; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_9_io_i_mux_bus_2 = PathFinder_9_io_i_mux_bus_2; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_9_io_i_mux_bus_3 = PathFinder_9_io_i_mux_bus_3; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_10_clock = clock;
  assign flexdpecom4_10_reset = reset;
  assign flexdpecom4_10_io_i_data_valid = 1'h1; // @[FlexDPU.scala 110:27 114:34]
  assign flexdpecom4_10_io_i_data_bus_0 = PathFinder_10_io_Source_0; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_10_io_i_data_bus_1 = PathFinder_10_io_Source_1; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_10_io_i_data_bus_2 = PathFinder_10_io_Source_2; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_10_io_i_data_bus_3 = PathFinder_10_io_Source_3; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_10_io_i_data_bus2_0 = PathFinder_10_io_destination_0; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_10_io_i_data_bus2_1 = PathFinder_10_io_destination_1; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_10_io_i_data_bus2_2 = PathFinder_10_io_destination_2; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_10_io_i_data_bus2_3 = PathFinder_10_io_destination_3; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_10_io_i_mux_bus_0 = PathFinder_10_io_i_mux_bus_0; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_10_io_i_mux_bus_1 = PathFinder_10_io_i_mux_bus_1; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_10_io_i_mux_bus_2 = PathFinder_10_io_i_mux_bus_2; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_10_io_i_mux_bus_3 = PathFinder_10_io_i_mux_bus_3; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_11_clock = clock;
  assign flexdpecom4_11_reset = reset;
  assign flexdpecom4_11_io_i_data_valid = 1'h1; // @[FlexDPU.scala 110:27 114:34]
  assign flexdpecom4_11_io_i_data_bus_0 = PathFinder_11_io_Source_0; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_11_io_i_data_bus_1 = PathFinder_11_io_Source_1; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_11_io_i_data_bus_2 = PathFinder_11_io_Source_2; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_11_io_i_data_bus_3 = PathFinder_11_io_Source_3; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_11_io_i_data_bus2_0 = PathFinder_11_io_destination_0; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_11_io_i_data_bus2_1 = PathFinder_11_io_destination_1; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_11_io_i_data_bus2_2 = PathFinder_11_io_destination_2; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_11_io_i_data_bus2_3 = PathFinder_11_io_destination_3; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_11_io_i_mux_bus_0 = PathFinder_11_io_i_mux_bus_0; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_11_io_i_mux_bus_1 = PathFinder_11_io_i_mux_bus_1; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_11_io_i_mux_bus_2 = PathFinder_11_io_i_mux_bus_2; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_11_io_i_mux_bus_3 = PathFinder_11_io_i_mux_bus_3; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_12_clock = clock;
  assign flexdpecom4_12_reset = reset;
  assign flexdpecom4_12_io_i_data_valid = 1'h1; // @[FlexDPU.scala 110:27 114:34]
  assign flexdpecom4_12_io_i_data_bus_0 = PathFinder_12_io_Source_0; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_12_io_i_data_bus_1 = PathFinder_12_io_Source_1; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_12_io_i_data_bus_2 = PathFinder_12_io_Source_2; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_12_io_i_data_bus_3 = PathFinder_12_io_Source_3; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_12_io_i_data_bus2_0 = PathFinder_12_io_destination_0; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_12_io_i_data_bus2_1 = PathFinder_12_io_destination_1; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_12_io_i_data_bus2_2 = PathFinder_12_io_destination_2; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_12_io_i_data_bus2_3 = PathFinder_12_io_destination_3; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_12_io_i_mux_bus_0 = PathFinder_12_io_i_mux_bus_0; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_12_io_i_mux_bus_1 = PathFinder_12_io_i_mux_bus_1; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_12_io_i_mux_bus_2 = PathFinder_12_io_i_mux_bus_2; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_12_io_i_mux_bus_3 = PathFinder_12_io_i_mux_bus_3; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_13_clock = clock;
  assign flexdpecom4_13_reset = reset;
  assign flexdpecom4_13_io_i_data_valid = 1'h1; // @[FlexDPU.scala 110:27 114:34]
  assign flexdpecom4_13_io_i_data_bus_0 = PathFinder_13_io_Source_0; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_13_io_i_data_bus_1 = PathFinder_13_io_Source_1; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_13_io_i_data_bus_2 = PathFinder_13_io_Source_2; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_13_io_i_data_bus_3 = PathFinder_13_io_Source_3; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_13_io_i_data_bus2_0 = PathFinder_13_io_destination_0; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_13_io_i_data_bus2_1 = PathFinder_13_io_destination_1; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_13_io_i_data_bus2_2 = PathFinder_13_io_destination_2; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_13_io_i_data_bus2_3 = PathFinder_13_io_destination_3; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_13_io_i_mux_bus_0 = PathFinder_13_io_i_mux_bus_0; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_13_io_i_mux_bus_1 = PathFinder_13_io_i_mux_bus_1; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_13_io_i_mux_bus_2 = PathFinder_13_io_i_mux_bus_2; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_13_io_i_mux_bus_3 = PathFinder_13_io_i_mux_bus_3; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_14_clock = clock;
  assign flexdpecom4_14_reset = reset;
  assign flexdpecom4_14_io_i_data_valid = 1'h1; // @[FlexDPU.scala 110:27 114:34]
  assign flexdpecom4_14_io_i_data_bus_0 = PathFinder_14_io_Source_0; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_14_io_i_data_bus_1 = PathFinder_14_io_Source_1; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_14_io_i_data_bus_2 = PathFinder_14_io_Source_2; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_14_io_i_data_bus_3 = PathFinder_14_io_Source_3; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_14_io_i_data_bus2_0 = PathFinder_14_io_destination_0; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_14_io_i_data_bus2_1 = PathFinder_14_io_destination_1; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_14_io_i_data_bus2_2 = PathFinder_14_io_destination_2; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_14_io_i_data_bus2_3 = PathFinder_14_io_destination_3; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_14_io_i_mux_bus_0 = PathFinder_14_io_i_mux_bus_0; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_14_io_i_mux_bus_1 = PathFinder_14_io_i_mux_bus_1; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_14_io_i_mux_bus_2 = PathFinder_14_io_i_mux_bus_2; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_14_io_i_mux_bus_3 = PathFinder_14_io_i_mux_bus_3; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_15_clock = clock;
  assign flexdpecom4_15_reset = reset;
  assign flexdpecom4_15_io_i_data_valid = 1'h1; // @[FlexDPU.scala 110:27 114:34]
  assign flexdpecom4_15_io_i_data_bus_0 = PathFinder_15_io_Source_0; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_15_io_i_data_bus_1 = PathFinder_15_io_Source_1; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_15_io_i_data_bus_2 = PathFinder_15_io_Source_2; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_15_io_i_data_bus_3 = PathFinder_15_io_Source_3; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_15_io_i_data_bus2_0 = PathFinder_15_io_destination_0; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_15_io_i_data_bus2_1 = PathFinder_15_io_destination_1; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_15_io_i_data_bus2_2 = PathFinder_15_io_destination_2; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_15_io_i_data_bus2_3 = PathFinder_15_io_destination_3; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_15_io_i_mux_bus_0 = PathFinder_15_io_i_mux_bus_0; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_15_io_i_mux_bus_1 = PathFinder_15_io_i_mux_bus_1; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_15_io_i_mux_bus_2 = PathFinder_15_io_i_mux_bus_2; // @[FlexDPU.scala 77:{21,21}]
  assign flexdpecom4_15_io_i_mux_bus_3 = PathFinder_15_io_i_mux_bus_3; // @[FlexDPU.scala 77:{21,21}]
  always @(posedge clock) begin
    if (2'h0 < remainingDistribution) begin // @[FlexDPU.scala 25:29]
      used_FlexDPE_0 <= _used_FlexDPE_0_T_2;
    end else begin
      used_FlexDPE_0 <= equalDistribution;
    end
    if (2'h1 < remainingDistribution) begin // @[FlexDPU.scala 25:29]
      used_FlexDPE_1 <= _used_FlexDPE_0_T_2;
    end else begin
      used_FlexDPE_1 <= equalDistribution;
    end
    if (reset) begin // @[FlexDPU.scala 33:24]
      iloop <= 32'h0; // @[FlexDPU.scala 33:24]
    end else if (iloop < 32'h7 & _Statvalid_T_1) begin // @[FlexDPU.scala 43:77]
      iloop <= _iloop_T_1; // @[FlexDPU.scala 44:15]
    end
    if (reset) begin // @[FlexDPU.scala 34:24]
      jloop <= 32'h0; // @[FlexDPU.scala 34:24]
    end else if (iloop <= 32'h7 & jloop < 32'h7) begin // @[FlexDPU.scala 47:76]
      jloop <= _jloop_T_1; // @[FlexDPU.scala 48:15]
    end else if (!(_Statvalid_T_2)) begin // @[FlexDPU.scala 49:83]
      jloop <= 32'h0; // @[FlexDPU.scala 52:15]
    end
    if (reset) begin // @[FlexDPU.scala 35:28]
      Statvalid <= 1'h0; // @[FlexDPU.scala 35:28]
    end else begin
      Statvalid <= iloop == 32'h7 & jloop == 32'h7; // @[FlexDPU.scala 37:15]
    end
    if (reset) begin // @[FlexDPU.scala 61:33]
      PF1_Stream_Col_0 <= 32'h0; // @[FlexDPU.scala 61:33]
    end else if (Statvalid) begin // @[FlexDPU.scala 98:20]
      PF1_Stream_Col_0 <= {{16'd0}, _GEN_269}; // @[FlexDPU.scala 164:31]
    end
    if (reset) begin // @[FlexDPU.scala 61:33]
      PF1_Stream_Col_1 <= 32'h0; // @[FlexDPU.scala 61:33]
    end else if (Statvalid) begin // @[FlexDPU.scala 98:20]
      PF1_Stream_Col_1 <= {{16'd0}, _GEN_277}; // @[FlexDPU.scala 164:31]
    end
    if (reset) begin // @[FlexDPU.scala 61:33]
      PF1_Stream_Col_2 <= 32'h0; // @[FlexDPU.scala 61:33]
    end else if (Statvalid) begin // @[FlexDPU.scala 98:20]
      PF1_Stream_Col_2 <= {{16'd0}, _GEN_285}; // @[FlexDPU.scala 164:31]
    end
    if (reset) begin // @[FlexDPU.scala 61:33]
      PF1_Stream_Col_3 <= 32'h0; // @[FlexDPU.scala 61:33]
    end else if (Statvalid) begin // @[FlexDPU.scala 98:20]
      PF1_Stream_Col_3 <= {{16'd0}, _GEN_293}; // @[FlexDPU.scala 164:31]
    end
    if (reset) begin // @[FlexDPU.scala 61:33]
      PF1_Stream_Col_4 <= 32'h0; // @[FlexDPU.scala 61:33]
    end else if (Statvalid) begin // @[FlexDPU.scala 98:20]
      PF1_Stream_Col_4 <= {{16'd0}, _GEN_301}; // @[FlexDPU.scala 164:31]
    end
    if (reset) begin // @[FlexDPU.scala 61:33]
      PF1_Stream_Col_5 <= 32'h0; // @[FlexDPU.scala 61:33]
    end else if (Statvalid) begin // @[FlexDPU.scala 98:20]
      PF1_Stream_Col_5 <= {{16'd0}, _GEN_309}; // @[FlexDPU.scala 164:31]
    end
    if (reset) begin // @[FlexDPU.scala 61:33]
      PF1_Stream_Col_6 <= 32'h0; // @[FlexDPU.scala 61:33]
    end else if (Statvalid) begin // @[FlexDPU.scala 98:20]
      PF1_Stream_Col_6 <= {{16'd0}, _GEN_317}; // @[FlexDPU.scala 164:31]
    end
    if (reset) begin // @[FlexDPU.scala 61:33]
      PF1_Stream_Col_7 <= 32'h0; // @[FlexDPU.scala 61:33]
    end else if (Statvalid) begin // @[FlexDPU.scala 98:20]
      PF1_Stream_Col_7 <= {{16'd0}, _GEN_325}; // @[FlexDPU.scala 164:31]
    end
    if (reset) begin // @[FlexDPU.scala 62:30]
      ModuleIndex <= 32'h0; // @[FlexDPU.scala 62:30]
    end else if (Statvalid) begin // @[FlexDPU.scala 98:20]
      if (!(ModuleIndex == 32'h7 & PF_0_PF_Valid)) begin // @[FlexDPU.scala 157:71]
        if (PF_0_PF_Valid) begin // @[FlexDPU.scala 152:29]
          ModuleIndex <= _ModuleIndex_T_1; // @[FlexDPU.scala 154:25]
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  used_FlexDPE_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  used_FlexDPE_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  iloop = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  jloop = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  Statvalid = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  PF1_Stream_Col_0 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  PF1_Stream_Col_1 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  PF1_Stream_Col_2 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  PF1_Stream_Col_3 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  PF1_Stream_Col_4 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  PF1_Stream_Col_5 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  PF1_Stream_Col_6 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  PF1_Stream_Col_7 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  ModuleIndex = _RAND_13[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
