/* verilator lint_off WIDTH */
module Bitmap(
  input         clock,
  input         reset,
  input  [15:0] io_mat1_0_0,
  input  [15:0] io_mat1_0_1,
  input  [15:0] io_mat1_0_2,
  input  [15:0] io_mat1_0_3,
  input  [15:0] io_mat1_0_4,
  input  [15:0] io_mat1_0_5,
  input  [15:0] io_mat1_0_6,
  input  [15:0] io_mat1_0_7,
  input  [15:0] io_mat1_1_0,
  input  [15:0] io_mat1_1_1,
  input  [15:0] io_mat1_1_2,
  input  [15:0] io_mat1_1_3,
  input  [15:0] io_mat1_1_4,
  input  [15:0] io_mat1_1_5,
  input  [15:0] io_mat1_1_6,
  input  [15:0] io_mat1_1_7,
  input  [15:0] io_mat1_2_0,
  input  [15:0] io_mat1_2_1,
  input  [15:0] io_mat1_2_2,
  input  [15:0] io_mat1_2_3,
  input  [15:0] io_mat1_2_4,
  input  [15:0] io_mat1_2_5,
  input  [15:0] io_mat1_2_6,
  input  [15:0] io_mat1_2_7,
  input  [15:0] io_mat1_3_0,
  input  [15:0] io_mat1_3_1,
  input  [15:0] io_mat1_3_2,
  input  [15:0] io_mat1_3_3,
  input  [15:0] io_mat1_3_4,
  input  [15:0] io_mat1_3_5,
  input  [15:0] io_mat1_3_6,
  input  [15:0] io_mat1_3_7,
  input  [15:0] io_mat1_4_0,
  input  [15:0] io_mat1_4_1,
  input  [15:0] io_mat1_4_2,
  input  [15:0] io_mat1_4_3,
  input  [15:0] io_mat1_4_4,
  input  [15:0] io_mat1_4_5,
  input  [15:0] io_mat1_4_6,
  input  [15:0] io_mat1_4_7,
  input  [15:0] io_mat1_5_0,
  input  [15:0] io_mat1_5_1,
  input  [15:0] io_mat1_5_2,
  input  [15:0] io_mat1_5_3,
  input  [15:0] io_mat1_5_4,
  input  [15:0] io_mat1_5_5,
  input  [15:0] io_mat1_5_6,
  input  [15:0] io_mat1_5_7,
  input  [15:0] io_mat1_6_0,
  input  [15:0] io_mat1_6_1,
  input  [15:0] io_mat1_6_2,
  input  [15:0] io_mat1_6_3,
  input  [15:0] io_mat1_6_4,
  input  [15:0] io_mat1_6_5,
  input  [15:0] io_mat1_6_6,
  input  [15:0] io_mat1_6_7,
  input  [15:0] io_mat1_7_0,
  input  [15:0] io_mat1_7_1,
  input  [15:0] io_mat1_7_2,
  input  [15:0] io_mat1_7_3,
  input  [15:0] io_mat1_7_4,
  input  [15:0] io_mat1_7_5,
  input  [15:0] io_mat1_7_6,
  input  [15:0] io_mat1_7_7,
  output [15:0] io_bitmap1_0_0,
  output [15:0] io_bitmap1_0_1,
  output [15:0] io_bitmap1_0_2,
  output [15:0] io_bitmap1_0_3,
  output [15:0] io_bitmap1_0_4,
  output [15:0] io_bitmap1_0_5,
  output [15:0] io_bitmap1_0_6,
  output [15:0] io_bitmap1_0_7,
  output [15:0] io_bitmap1_1_0,
  output [15:0] io_bitmap1_1_1,
  output [15:0] io_bitmap1_1_2,
  output [15:0] io_bitmap1_1_3,
  output [15:0] io_bitmap1_1_4,
  output [15:0] io_bitmap1_1_5,
  output [15:0] io_bitmap1_1_6,
  output [15:0] io_bitmap1_1_7,
  output [15:0] io_bitmap1_2_0,
  output [15:0] io_bitmap1_2_1,
  output [15:0] io_bitmap1_2_2,
  output [15:0] io_bitmap1_2_3,
  output [15:0] io_bitmap1_2_4,
  output [15:0] io_bitmap1_2_5,
  output [15:0] io_bitmap1_2_6,
  output [15:0] io_bitmap1_2_7,
  output [15:0] io_bitmap1_3_0,
  output [15:0] io_bitmap1_3_1,
  output [15:0] io_bitmap1_3_2,
  output [15:0] io_bitmap1_3_3,
  output [15:0] io_bitmap1_3_4,
  output [15:0] io_bitmap1_3_5,
  output [15:0] io_bitmap1_3_6,
  output [15:0] io_bitmap1_3_7,
  output [15:0] io_bitmap1_4_0,
  output [15:0] io_bitmap1_4_1,
  output [15:0] io_bitmap1_4_2,
  output [15:0] io_bitmap1_4_3,
  output [15:0] io_bitmap1_4_4,
  output [15:0] io_bitmap1_4_5,
  output [15:0] io_bitmap1_4_6,
  output [15:0] io_bitmap1_4_7,
  output [15:0] io_bitmap1_5_0,
  output [15:0] io_bitmap1_5_1,
  output [15:0] io_bitmap1_5_2,
  output [15:0] io_bitmap1_5_3,
  output [15:0] io_bitmap1_5_4,
  output [15:0] io_bitmap1_5_5,
  output [15:0] io_bitmap1_5_6,
  output [15:0] io_bitmap1_5_7,
  output [15:0] io_bitmap1_6_0,
  output [15:0] io_bitmap1_6_1,
  output [15:0] io_bitmap1_6_2,
  output [15:0] io_bitmap1_6_3,
  output [15:0] io_bitmap1_6_4,
  output [15:0] io_bitmap1_6_5,
  output [15:0] io_bitmap1_6_6,
  output [15:0] io_bitmap1_6_7,
  output [15:0] io_bitmap1_7_0,
  output [15:0] io_bitmap1_7_1,
  output [15:0] io_bitmap1_7_2,
  output [15:0] io_bitmap1_7_3,
  output [15:0] io_bitmap1_7_4,
  output [15:0] io_bitmap1_7_5,
  output [15:0] io_bitmap1_7_6,
  output [15:0] io_bitmap1_7_7
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
`endif // RANDOMIZE_REG_INIT
  reg [15:0] matReg1_0_0; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_0_1; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_0_2; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_0_3; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_0_4; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_0_5; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_0_6; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_0_7; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_1_0; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_1_1; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_1_2; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_1_3; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_1_4; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_1_5; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_1_6; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_1_7; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_2_0; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_2_1; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_2_2; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_2_3; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_2_4; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_2_5; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_2_6; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_2_7; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_3_0; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_3_1; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_3_2; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_3_3; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_3_4; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_3_5; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_3_6; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_3_7; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_4_0; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_4_1; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_4_2; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_4_3; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_4_4; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_4_5; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_4_6; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_4_7; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_5_0; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_5_1; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_5_2; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_5_3; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_5_4; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_5_5; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_5_6; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_5_7; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_6_0; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_6_1; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_6_2; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_6_3; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_6_4; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_6_5; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_6_6; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_6_7; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_7_0; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_7_1; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_7_2; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_7_3; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_7_4; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_7_5; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_7_6; // @[Bitmap.scala 14:26]
  reg [15:0] matReg1_7_7; // @[Bitmap.scala 14:26]
  reg [2:0] i; // @[Bitmap.scala 19:20]
  reg [2:0] j; // @[Bitmap.scala 20:20]
  wire  _GEN_642 = 3'h0 == i; // @[Bitmap.scala 23:{41,41}]
  wire  _GEN_643 = 3'h1 == j; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_1 = 3'h0 == i & 3'h1 == j ? io_mat1_0_1 : io_mat1_0_0; // @[Bitmap.scala 23:{41,41}]
  wire  _GEN_645 = 3'h2 == j; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_2 = 3'h0 == i & 3'h2 == j ? io_mat1_0_2 : _GEN_1; // @[Bitmap.scala 23:{41,41}]
  wire  _GEN_647 = 3'h3 == j; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_3 = 3'h0 == i & 3'h3 == j ? io_mat1_0_3 : _GEN_2; // @[Bitmap.scala 23:{41,41}]
  wire  _GEN_649 = 3'h4 == j; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_4 = 3'h0 == i & 3'h4 == j ? io_mat1_0_4 : _GEN_3; // @[Bitmap.scala 23:{41,41}]
  wire  _GEN_651 = 3'h5 == j; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_5 = 3'h0 == i & 3'h5 == j ? io_mat1_0_5 : _GEN_4; // @[Bitmap.scala 23:{41,41}]
  wire  _GEN_653 = 3'h6 == j; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_6 = 3'h0 == i & 3'h6 == j ? io_mat1_0_6 : _GEN_5; // @[Bitmap.scala 23:{41,41}]
  wire  _GEN_655 = 3'h7 == j; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_7 = 3'h0 == i & 3'h7 == j ? io_mat1_0_7 : _GEN_6; // @[Bitmap.scala 23:{41,41}]
  wire  _GEN_656 = 3'h1 == i; // @[Bitmap.scala 23:{41,41}]
  wire  _GEN_657 = 3'h0 == j; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_8 = 3'h1 == i & 3'h0 == j ? io_mat1_1_0 : _GEN_7; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_9 = 3'h1 == i & 3'h1 == j ? io_mat1_1_1 : _GEN_8; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_10 = 3'h1 == i & 3'h2 == j ? io_mat1_1_2 : _GEN_9; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_11 = 3'h1 == i & 3'h3 == j ? io_mat1_1_3 : _GEN_10; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_12 = 3'h1 == i & 3'h4 == j ? io_mat1_1_4 : _GEN_11; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_13 = 3'h1 == i & 3'h5 == j ? io_mat1_1_5 : _GEN_12; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_14 = 3'h1 == i & 3'h6 == j ? io_mat1_1_6 : _GEN_13; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_15 = 3'h1 == i & 3'h7 == j ? io_mat1_1_7 : _GEN_14; // @[Bitmap.scala 23:{41,41}]
  wire  _GEN_672 = 3'h2 == i; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_16 = 3'h2 == i & 3'h0 == j ? io_mat1_2_0 : _GEN_15; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_17 = 3'h2 == i & 3'h1 == j ? io_mat1_2_1 : _GEN_16; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_18 = 3'h2 == i & 3'h2 == j ? io_mat1_2_2 : _GEN_17; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_19 = 3'h2 == i & 3'h3 == j ? io_mat1_2_3 : _GEN_18; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_20 = 3'h2 == i & 3'h4 == j ? io_mat1_2_4 : _GEN_19; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_21 = 3'h2 == i & 3'h5 == j ? io_mat1_2_5 : _GEN_20; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_22 = 3'h2 == i & 3'h6 == j ? io_mat1_2_6 : _GEN_21; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_23 = 3'h2 == i & 3'h7 == j ? io_mat1_2_7 : _GEN_22; // @[Bitmap.scala 23:{41,41}]
  wire  _GEN_688 = 3'h3 == i; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_24 = 3'h3 == i & 3'h0 == j ? io_mat1_3_0 : _GEN_23; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_25 = 3'h3 == i & 3'h1 == j ? io_mat1_3_1 : _GEN_24; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_26 = 3'h3 == i & 3'h2 == j ? io_mat1_3_2 : _GEN_25; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_27 = 3'h3 == i & 3'h3 == j ? io_mat1_3_3 : _GEN_26; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_28 = 3'h3 == i & 3'h4 == j ? io_mat1_3_4 : _GEN_27; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_29 = 3'h3 == i & 3'h5 == j ? io_mat1_3_5 : _GEN_28; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_30 = 3'h3 == i & 3'h6 == j ? io_mat1_3_6 : _GEN_29; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_31 = 3'h3 == i & 3'h7 == j ? io_mat1_3_7 : _GEN_30; // @[Bitmap.scala 23:{41,41}]
  wire  _GEN_704 = 3'h4 == i; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_32 = 3'h4 == i & 3'h0 == j ? io_mat1_4_0 : _GEN_31; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_33 = 3'h4 == i & 3'h1 == j ? io_mat1_4_1 : _GEN_32; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_34 = 3'h4 == i & 3'h2 == j ? io_mat1_4_2 : _GEN_33; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_35 = 3'h4 == i & 3'h3 == j ? io_mat1_4_3 : _GEN_34; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_36 = 3'h4 == i & 3'h4 == j ? io_mat1_4_4 : _GEN_35; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_37 = 3'h4 == i & 3'h5 == j ? io_mat1_4_5 : _GEN_36; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_38 = 3'h4 == i & 3'h6 == j ? io_mat1_4_6 : _GEN_37; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_39 = 3'h4 == i & 3'h7 == j ? io_mat1_4_7 : _GEN_38; // @[Bitmap.scala 23:{41,41}]
  wire  _GEN_720 = 3'h5 == i; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_40 = 3'h5 == i & 3'h0 == j ? io_mat1_5_0 : _GEN_39; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_41 = 3'h5 == i & 3'h1 == j ? io_mat1_5_1 : _GEN_40; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_42 = 3'h5 == i & 3'h2 == j ? io_mat1_5_2 : _GEN_41; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_43 = 3'h5 == i & 3'h3 == j ? io_mat1_5_3 : _GEN_42; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_44 = 3'h5 == i & 3'h4 == j ? io_mat1_5_4 : _GEN_43; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_45 = 3'h5 == i & 3'h5 == j ? io_mat1_5_5 : _GEN_44; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_46 = 3'h5 == i & 3'h6 == j ? io_mat1_5_6 : _GEN_45; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_47 = 3'h5 == i & 3'h7 == j ? io_mat1_5_7 : _GEN_46; // @[Bitmap.scala 23:{41,41}]
  wire  _GEN_736 = 3'h6 == i; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_48 = 3'h6 == i & 3'h0 == j ? io_mat1_6_0 : _GEN_47; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_49 = 3'h6 == i & 3'h1 == j ? io_mat1_6_1 : _GEN_48; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_50 = 3'h6 == i & 3'h2 == j ? io_mat1_6_2 : _GEN_49; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_51 = 3'h6 == i & 3'h3 == j ? io_mat1_6_3 : _GEN_50; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_52 = 3'h6 == i & 3'h4 == j ? io_mat1_6_4 : _GEN_51; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_53 = 3'h6 == i & 3'h5 == j ? io_mat1_6_5 : _GEN_52; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_54 = 3'h6 == i & 3'h6 == j ? io_mat1_6_6 : _GEN_53; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_55 = 3'h6 == i & 3'h7 == j ? io_mat1_6_7 : _GEN_54; // @[Bitmap.scala 23:{41,41}]
  wire  _GEN_752 = 3'h7 == i; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_56 = 3'h7 == i & 3'h0 == j ? io_mat1_7_0 : _GEN_55; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_57 = 3'h7 == i & 3'h1 == j ? io_mat1_7_1 : _GEN_56; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_58 = 3'h7 == i & 3'h2 == j ? io_mat1_7_2 : _GEN_57; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_59 = 3'h7 == i & 3'h3 == j ? io_mat1_7_3 : _GEN_58; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_60 = 3'h7 == i & 3'h4 == j ? io_mat1_7_4 : _GEN_59; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_61 = 3'h7 == i & 3'h5 == j ? io_mat1_7_5 : _GEN_60; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_62 = 3'h7 == i & 3'h6 == j ? io_mat1_7_6 : _GEN_61; // @[Bitmap.scala 23:{41,41}]
  wire [15:0] _GEN_63 = 3'h7 == i & 3'h7 == j ? io_mat1_7_7 : _GEN_62; // @[Bitmap.scala 23:{41,41}]
  wire [2:0] _j_T_1 = j + 3'h1; // @[Bitmap.scala 33:17]
  wire [2:0] _i_T_1 = i + 3'h1; // @[Bitmap.scala 36:12]
  assign io_bitmap1_0_0 = matReg1_0_0; // @[Bitmap.scala 16:16]
  assign io_bitmap1_0_1 = matReg1_0_1; // @[Bitmap.scala 16:16]
  assign io_bitmap1_0_2 = matReg1_0_2; // @[Bitmap.scala 16:16]
  assign io_bitmap1_0_3 = matReg1_0_3; // @[Bitmap.scala 16:16]
  assign io_bitmap1_0_4 = matReg1_0_4; // @[Bitmap.scala 16:16]
  assign io_bitmap1_0_5 = matReg1_0_5; // @[Bitmap.scala 16:16]
  assign io_bitmap1_0_6 = matReg1_0_6; // @[Bitmap.scala 16:16]
  assign io_bitmap1_0_7 = matReg1_0_7; // @[Bitmap.scala 16:16]
  assign io_bitmap1_1_0 = matReg1_1_0; // @[Bitmap.scala 16:16]
  assign io_bitmap1_1_1 = matReg1_1_1; // @[Bitmap.scala 16:16]
  assign io_bitmap1_1_2 = matReg1_1_2; // @[Bitmap.scala 16:16]
  assign io_bitmap1_1_3 = matReg1_1_3; // @[Bitmap.scala 16:16]
  assign io_bitmap1_1_4 = matReg1_1_4; // @[Bitmap.scala 16:16]
  assign io_bitmap1_1_5 = matReg1_1_5; // @[Bitmap.scala 16:16]
  assign io_bitmap1_1_6 = matReg1_1_6; // @[Bitmap.scala 16:16]
  assign io_bitmap1_1_7 = matReg1_1_7; // @[Bitmap.scala 16:16]
  assign io_bitmap1_2_0 = matReg1_2_0; // @[Bitmap.scala 16:16]
  assign io_bitmap1_2_1 = matReg1_2_1; // @[Bitmap.scala 16:16]
  assign io_bitmap1_2_2 = matReg1_2_2; // @[Bitmap.scala 16:16]
  assign io_bitmap1_2_3 = matReg1_2_3; // @[Bitmap.scala 16:16]
  assign io_bitmap1_2_4 = matReg1_2_4; // @[Bitmap.scala 16:16]
  assign io_bitmap1_2_5 = matReg1_2_5; // @[Bitmap.scala 16:16]
  assign io_bitmap1_2_6 = matReg1_2_6; // @[Bitmap.scala 16:16]
  assign io_bitmap1_2_7 = matReg1_2_7; // @[Bitmap.scala 16:16]
  assign io_bitmap1_3_0 = matReg1_3_0; // @[Bitmap.scala 16:16]
  assign io_bitmap1_3_1 = matReg1_3_1; // @[Bitmap.scala 16:16]
  assign io_bitmap1_3_2 = matReg1_3_2; // @[Bitmap.scala 16:16]
  assign io_bitmap1_3_3 = matReg1_3_3; // @[Bitmap.scala 16:16]
  assign io_bitmap1_3_4 = matReg1_3_4; // @[Bitmap.scala 16:16]
  assign io_bitmap1_3_5 = matReg1_3_5; // @[Bitmap.scala 16:16]
  assign io_bitmap1_3_6 = matReg1_3_6; // @[Bitmap.scala 16:16]
  assign io_bitmap1_3_7 = matReg1_3_7; // @[Bitmap.scala 16:16]
  assign io_bitmap1_4_0 = matReg1_4_0; // @[Bitmap.scala 16:16]
  assign io_bitmap1_4_1 = matReg1_4_1; // @[Bitmap.scala 16:16]
  assign io_bitmap1_4_2 = matReg1_4_2; // @[Bitmap.scala 16:16]
  assign io_bitmap1_4_3 = matReg1_4_3; // @[Bitmap.scala 16:16]
  assign io_bitmap1_4_4 = matReg1_4_4; // @[Bitmap.scala 16:16]
  assign io_bitmap1_4_5 = matReg1_4_5; // @[Bitmap.scala 16:16]
  assign io_bitmap1_4_6 = matReg1_4_6; // @[Bitmap.scala 16:16]
  assign io_bitmap1_4_7 = matReg1_4_7; // @[Bitmap.scala 16:16]
  assign io_bitmap1_5_0 = matReg1_5_0; // @[Bitmap.scala 16:16]
  assign io_bitmap1_5_1 = matReg1_5_1; // @[Bitmap.scala 16:16]
  assign io_bitmap1_5_2 = matReg1_5_2; // @[Bitmap.scala 16:16]
  assign io_bitmap1_5_3 = matReg1_5_3; // @[Bitmap.scala 16:16]
  assign io_bitmap1_5_4 = matReg1_5_4; // @[Bitmap.scala 16:16]
  assign io_bitmap1_5_5 = matReg1_5_5; // @[Bitmap.scala 16:16]
  assign io_bitmap1_5_6 = matReg1_5_6; // @[Bitmap.scala 16:16]
  assign io_bitmap1_5_7 = matReg1_5_7; // @[Bitmap.scala 16:16]
  assign io_bitmap1_6_0 = matReg1_6_0; // @[Bitmap.scala 16:16]
  assign io_bitmap1_6_1 = matReg1_6_1; // @[Bitmap.scala 16:16]
  assign io_bitmap1_6_2 = matReg1_6_2; // @[Bitmap.scala 16:16]
  assign io_bitmap1_6_3 = matReg1_6_3; // @[Bitmap.scala 16:16]
  assign io_bitmap1_6_4 = matReg1_6_4; // @[Bitmap.scala 16:16]
  assign io_bitmap1_6_5 = matReg1_6_5; // @[Bitmap.scala 16:16]
  assign io_bitmap1_6_6 = matReg1_6_6; // @[Bitmap.scala 16:16]
  assign io_bitmap1_6_7 = matReg1_6_7; // @[Bitmap.scala 16:16]
  assign io_bitmap1_7_0 = matReg1_7_0; // @[Bitmap.scala 16:16]
  assign io_bitmap1_7_1 = matReg1_7_1; // @[Bitmap.scala 16:16]
  assign io_bitmap1_7_2 = matReg1_7_2; // @[Bitmap.scala 16:16]
  assign io_bitmap1_7_3 = matReg1_7_3; // @[Bitmap.scala 16:16]
  assign io_bitmap1_7_4 = matReg1_7_4; // @[Bitmap.scala 16:16]
  assign io_bitmap1_7_5 = matReg1_7_5; // @[Bitmap.scala 16:16]
  assign io_bitmap1_7_6 = matReg1_7_6; // @[Bitmap.scala 16:16]
  assign io_bitmap1_7_7 = matReg1_7_7; // @[Bitmap.scala 16:16]
  always @(posedge clock) begin
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_0_0 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_642 & _GEN_657) begin // @[Bitmap.scala 24:31]
        matReg1_0_0 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_642 & _GEN_657) begin // @[Bitmap.scala 26:31]
      matReg1_0_0 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_0_1 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_642 & _GEN_643) begin // @[Bitmap.scala 24:31]
        matReg1_0_1 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_642 & _GEN_643) begin // @[Bitmap.scala 26:31]
      matReg1_0_1 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_0_2 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_642 & _GEN_645) begin // @[Bitmap.scala 24:31]
        matReg1_0_2 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_642 & _GEN_645) begin // @[Bitmap.scala 26:31]
      matReg1_0_2 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_0_3 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_642 & _GEN_647) begin // @[Bitmap.scala 24:31]
        matReg1_0_3 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_642 & _GEN_647) begin // @[Bitmap.scala 26:31]
      matReg1_0_3 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_0_4 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_642 & _GEN_649) begin // @[Bitmap.scala 24:31]
        matReg1_0_4 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_642 & _GEN_649) begin // @[Bitmap.scala 26:31]
      matReg1_0_4 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_0_5 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_642 & _GEN_651) begin // @[Bitmap.scala 24:31]
        matReg1_0_5 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_642 & _GEN_651) begin // @[Bitmap.scala 26:31]
      matReg1_0_5 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_0_6 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_642 & _GEN_653) begin // @[Bitmap.scala 24:31]
        matReg1_0_6 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_642 & _GEN_653) begin // @[Bitmap.scala 26:31]
      matReg1_0_6 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_0_7 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_642 & _GEN_655) begin // @[Bitmap.scala 24:31]
        matReg1_0_7 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_642 & _GEN_655) begin // @[Bitmap.scala 26:31]
      matReg1_0_7 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_1_0 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_656 & _GEN_657) begin // @[Bitmap.scala 24:31]
        matReg1_1_0 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_656 & _GEN_657) begin // @[Bitmap.scala 26:31]
      matReg1_1_0 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_1_1 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_656 & _GEN_643) begin // @[Bitmap.scala 24:31]
        matReg1_1_1 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_656 & _GEN_643) begin // @[Bitmap.scala 26:31]
      matReg1_1_1 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_1_2 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_656 & _GEN_645) begin // @[Bitmap.scala 24:31]
        matReg1_1_2 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_656 & _GEN_645) begin // @[Bitmap.scala 26:31]
      matReg1_1_2 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_1_3 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_656 & _GEN_647) begin // @[Bitmap.scala 24:31]
        matReg1_1_3 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_656 & _GEN_647) begin // @[Bitmap.scala 26:31]
      matReg1_1_3 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_1_4 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_656 & _GEN_649) begin // @[Bitmap.scala 24:31]
        matReg1_1_4 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_656 & _GEN_649) begin // @[Bitmap.scala 26:31]
      matReg1_1_4 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_1_5 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_656 & _GEN_651) begin // @[Bitmap.scala 24:31]
        matReg1_1_5 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_656 & _GEN_651) begin // @[Bitmap.scala 26:31]
      matReg1_1_5 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_1_6 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_656 & _GEN_653) begin // @[Bitmap.scala 24:31]
        matReg1_1_6 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_656 & _GEN_653) begin // @[Bitmap.scala 26:31]
      matReg1_1_6 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_1_7 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_656 & _GEN_655) begin // @[Bitmap.scala 24:31]
        matReg1_1_7 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_656 & _GEN_655) begin // @[Bitmap.scala 26:31]
      matReg1_1_7 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_2_0 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_672 & _GEN_657) begin // @[Bitmap.scala 24:31]
        matReg1_2_0 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_672 & _GEN_657) begin // @[Bitmap.scala 26:31]
      matReg1_2_0 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_2_1 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_672 & _GEN_643) begin // @[Bitmap.scala 24:31]
        matReg1_2_1 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_672 & _GEN_643) begin // @[Bitmap.scala 26:31]
      matReg1_2_1 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_2_2 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_672 & _GEN_645) begin // @[Bitmap.scala 24:31]
        matReg1_2_2 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_672 & _GEN_645) begin // @[Bitmap.scala 26:31]
      matReg1_2_2 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_2_3 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_672 & _GEN_647) begin // @[Bitmap.scala 24:31]
        matReg1_2_3 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_672 & _GEN_647) begin // @[Bitmap.scala 26:31]
      matReg1_2_3 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_2_4 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_672 & _GEN_649) begin // @[Bitmap.scala 24:31]
        matReg1_2_4 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_672 & _GEN_649) begin // @[Bitmap.scala 26:31]
      matReg1_2_4 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_2_5 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_672 & _GEN_651) begin // @[Bitmap.scala 24:31]
        matReg1_2_5 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_672 & _GEN_651) begin // @[Bitmap.scala 26:31]
      matReg1_2_5 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_2_6 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_672 & _GEN_653) begin // @[Bitmap.scala 24:31]
        matReg1_2_6 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_672 & _GEN_653) begin // @[Bitmap.scala 26:31]
      matReg1_2_6 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_2_7 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_672 & _GEN_655) begin // @[Bitmap.scala 24:31]
        matReg1_2_7 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_672 & _GEN_655) begin // @[Bitmap.scala 26:31]
      matReg1_2_7 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_3_0 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_688 & _GEN_657) begin // @[Bitmap.scala 24:31]
        matReg1_3_0 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_688 & _GEN_657) begin // @[Bitmap.scala 26:31]
      matReg1_3_0 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_3_1 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_688 & _GEN_643) begin // @[Bitmap.scala 24:31]
        matReg1_3_1 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_688 & _GEN_643) begin // @[Bitmap.scala 26:31]
      matReg1_3_1 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_3_2 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_688 & _GEN_645) begin // @[Bitmap.scala 24:31]
        matReg1_3_2 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_688 & _GEN_645) begin // @[Bitmap.scala 26:31]
      matReg1_3_2 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_3_3 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_688 & _GEN_647) begin // @[Bitmap.scala 24:31]
        matReg1_3_3 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_688 & _GEN_647) begin // @[Bitmap.scala 26:31]
      matReg1_3_3 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_3_4 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_688 & _GEN_649) begin // @[Bitmap.scala 24:31]
        matReg1_3_4 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_688 & _GEN_649) begin // @[Bitmap.scala 26:31]
      matReg1_3_4 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_3_5 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_688 & _GEN_651) begin // @[Bitmap.scala 24:31]
        matReg1_3_5 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_688 & _GEN_651) begin // @[Bitmap.scala 26:31]
      matReg1_3_5 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_3_6 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_688 & _GEN_653) begin // @[Bitmap.scala 24:31]
        matReg1_3_6 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_688 & _GEN_653) begin // @[Bitmap.scala 26:31]
      matReg1_3_6 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_3_7 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_688 & _GEN_655) begin // @[Bitmap.scala 24:31]
        matReg1_3_7 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_688 & _GEN_655) begin // @[Bitmap.scala 26:31]
      matReg1_3_7 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_4_0 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_704 & _GEN_657) begin // @[Bitmap.scala 24:31]
        matReg1_4_0 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_704 & _GEN_657) begin // @[Bitmap.scala 26:31]
      matReg1_4_0 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_4_1 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_704 & _GEN_643) begin // @[Bitmap.scala 24:31]
        matReg1_4_1 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_704 & _GEN_643) begin // @[Bitmap.scala 26:31]
      matReg1_4_1 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_4_2 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_704 & _GEN_645) begin // @[Bitmap.scala 24:31]
        matReg1_4_2 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_704 & _GEN_645) begin // @[Bitmap.scala 26:31]
      matReg1_4_2 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_4_3 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_704 & _GEN_647) begin // @[Bitmap.scala 24:31]
        matReg1_4_3 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_704 & _GEN_647) begin // @[Bitmap.scala 26:31]
      matReg1_4_3 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_4_4 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_704 & _GEN_649) begin // @[Bitmap.scala 24:31]
        matReg1_4_4 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_704 & _GEN_649) begin // @[Bitmap.scala 26:31]
      matReg1_4_4 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_4_5 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_704 & _GEN_651) begin // @[Bitmap.scala 24:31]
        matReg1_4_5 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_704 & _GEN_651) begin // @[Bitmap.scala 26:31]
      matReg1_4_5 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_4_6 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_704 & _GEN_653) begin // @[Bitmap.scala 24:31]
        matReg1_4_6 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_704 & _GEN_653) begin // @[Bitmap.scala 26:31]
      matReg1_4_6 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_4_7 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_704 & _GEN_655) begin // @[Bitmap.scala 24:31]
        matReg1_4_7 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_704 & _GEN_655) begin // @[Bitmap.scala 26:31]
      matReg1_4_7 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_5_0 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_720 & _GEN_657) begin // @[Bitmap.scala 24:31]
        matReg1_5_0 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_720 & _GEN_657) begin // @[Bitmap.scala 26:31]
      matReg1_5_0 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_5_1 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_720 & _GEN_643) begin // @[Bitmap.scala 24:31]
        matReg1_5_1 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_720 & _GEN_643) begin // @[Bitmap.scala 26:31]
      matReg1_5_1 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_5_2 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_720 & _GEN_645) begin // @[Bitmap.scala 24:31]
        matReg1_5_2 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_720 & _GEN_645) begin // @[Bitmap.scala 26:31]
      matReg1_5_2 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_5_3 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_720 & _GEN_647) begin // @[Bitmap.scala 24:31]
        matReg1_5_3 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_720 & _GEN_647) begin // @[Bitmap.scala 26:31]
      matReg1_5_3 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_5_4 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_720 & _GEN_649) begin // @[Bitmap.scala 24:31]
        matReg1_5_4 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_720 & _GEN_649) begin // @[Bitmap.scala 26:31]
      matReg1_5_4 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_5_5 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_720 & _GEN_651) begin // @[Bitmap.scala 24:31]
        matReg1_5_5 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_720 & _GEN_651) begin // @[Bitmap.scala 26:31]
      matReg1_5_5 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_5_6 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_720 & _GEN_653) begin // @[Bitmap.scala 24:31]
        matReg1_5_6 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_720 & _GEN_653) begin // @[Bitmap.scala 26:31]
      matReg1_5_6 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_5_7 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_720 & _GEN_655) begin // @[Bitmap.scala 24:31]
        matReg1_5_7 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_720 & _GEN_655) begin // @[Bitmap.scala 26:31]
      matReg1_5_7 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_6_0 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_736 & _GEN_657) begin // @[Bitmap.scala 24:31]
        matReg1_6_0 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_736 & _GEN_657) begin // @[Bitmap.scala 26:31]
      matReg1_6_0 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_6_1 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_736 & _GEN_643) begin // @[Bitmap.scala 24:31]
        matReg1_6_1 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_736 & _GEN_643) begin // @[Bitmap.scala 26:31]
      matReg1_6_1 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_6_2 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_736 & _GEN_645) begin // @[Bitmap.scala 24:31]
        matReg1_6_2 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_736 & _GEN_645) begin // @[Bitmap.scala 26:31]
      matReg1_6_2 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_6_3 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_736 & _GEN_647) begin // @[Bitmap.scala 24:31]
        matReg1_6_3 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_736 & _GEN_647) begin // @[Bitmap.scala 26:31]
      matReg1_6_3 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_6_4 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_736 & _GEN_649) begin // @[Bitmap.scala 24:31]
        matReg1_6_4 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_736 & _GEN_649) begin // @[Bitmap.scala 26:31]
      matReg1_6_4 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_6_5 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_736 & _GEN_651) begin // @[Bitmap.scala 24:31]
        matReg1_6_5 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_736 & _GEN_651) begin // @[Bitmap.scala 26:31]
      matReg1_6_5 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_6_6 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_736 & _GEN_653) begin // @[Bitmap.scala 24:31]
        matReg1_6_6 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_736 & _GEN_653) begin // @[Bitmap.scala 26:31]
      matReg1_6_6 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_6_7 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_736 & _GEN_655) begin // @[Bitmap.scala 24:31]
        matReg1_6_7 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_736 & _GEN_655) begin // @[Bitmap.scala 26:31]
      matReg1_6_7 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_7_0 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_752 & _GEN_657) begin // @[Bitmap.scala 24:31]
        matReg1_7_0 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_752 & _GEN_657) begin // @[Bitmap.scala 26:31]
      matReg1_7_0 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_7_1 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_752 & _GEN_643) begin // @[Bitmap.scala 24:31]
        matReg1_7_1 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_752 & _GEN_643) begin // @[Bitmap.scala 26:31]
      matReg1_7_1 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_7_2 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_752 & _GEN_645) begin // @[Bitmap.scala 24:31]
        matReg1_7_2 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_752 & _GEN_645) begin // @[Bitmap.scala 26:31]
      matReg1_7_2 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_7_3 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_752 & _GEN_647) begin // @[Bitmap.scala 24:31]
        matReg1_7_3 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_752 & _GEN_647) begin // @[Bitmap.scala 26:31]
      matReg1_7_3 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_7_4 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_752 & _GEN_649) begin // @[Bitmap.scala 24:31]
        matReg1_7_4 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_752 & _GEN_649) begin // @[Bitmap.scala 26:31]
      matReg1_7_4 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_7_5 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_752 & _GEN_651) begin // @[Bitmap.scala 24:31]
        matReg1_7_5 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_752 & _GEN_651) begin // @[Bitmap.scala 26:31]
      matReg1_7_5 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_7_6 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_752 & _GEN_653) begin // @[Bitmap.scala 24:31]
        matReg1_7_6 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_752 & _GEN_653) begin // @[Bitmap.scala 26:31]
      matReg1_7_6 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 14:26]
      matReg1_7_7 <= 16'h0; // @[Bitmap.scala 14:26]
    end else if (_GEN_63 != 16'h0) begin // @[Bitmap.scala 23:49]
      if (_GEN_752 & _GEN_655) begin // @[Bitmap.scala 24:31]
        matReg1_7_7 <= 16'h1; // @[Bitmap.scala 24:31]
      end
    end else if (_GEN_752 & _GEN_655) begin // @[Bitmap.scala 26:31]
      matReg1_7_7 <= 16'h0; // @[Bitmap.scala 26:31]
    end
    if (reset) begin // @[Bitmap.scala 19:20]
      i <= 3'h0; // @[Bitmap.scala 19:20]
    end else if (j == 3'h7) begin // @[Bitmap.scala 35:36]
      i <= _i_T_1; // @[Bitmap.scala 36:7]
    end
    if (reset) begin // @[Bitmap.scala 20:20]
      j <= 3'h0; // @[Bitmap.scala 20:20]
    end else begin
      j <= _j_T_1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  matReg1_0_0 = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  matReg1_0_1 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  matReg1_0_2 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  matReg1_0_3 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  matReg1_0_4 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  matReg1_0_5 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  matReg1_0_6 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  matReg1_0_7 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  matReg1_1_0 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  matReg1_1_1 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  matReg1_1_2 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  matReg1_1_3 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  matReg1_1_4 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  matReg1_1_5 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  matReg1_1_6 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  matReg1_1_7 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  matReg1_2_0 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  matReg1_2_1 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  matReg1_2_2 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  matReg1_2_3 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  matReg1_2_4 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  matReg1_2_5 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  matReg1_2_6 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  matReg1_2_7 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  matReg1_3_0 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  matReg1_3_1 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  matReg1_3_2 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  matReg1_3_3 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  matReg1_3_4 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  matReg1_3_5 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  matReg1_3_6 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  matReg1_3_7 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  matReg1_4_0 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  matReg1_4_1 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  matReg1_4_2 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  matReg1_4_3 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  matReg1_4_4 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  matReg1_4_5 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  matReg1_4_6 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  matReg1_4_7 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  matReg1_5_0 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  matReg1_5_1 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  matReg1_5_2 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  matReg1_5_3 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  matReg1_5_4 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  matReg1_5_5 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  matReg1_5_6 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  matReg1_5_7 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  matReg1_6_0 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  matReg1_6_1 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  matReg1_6_2 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  matReg1_6_3 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  matReg1_6_4 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  matReg1_6_5 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  matReg1_6_6 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  matReg1_6_7 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  matReg1_7_0 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  matReg1_7_1 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  matReg1_7_2 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  matReg1_7_3 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  matReg1_7_4 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  matReg1_7_5 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  matReg1_7_6 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  matReg1_7_7 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  i = _RAND_64[2:0];
  _RAND_65 = {1{`RANDOM}};
  j = _RAND_65[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Regor(
  input         clock,
  input         reset,
  input  [15:0] io_mat1_0_0,
  input  [15:0] io_mat1_0_1,
  input  [15:0] io_mat1_0_2,
  input  [15:0] io_mat1_0_3,
  input  [15:0] io_mat1_0_4,
  input  [15:0] io_mat1_0_5,
  input  [15:0] io_mat1_0_6,
  input  [15:0] io_mat1_0_7,
  input  [15:0] io_mat1_1_0,
  input  [15:0] io_mat1_1_1,
  input  [15:0] io_mat1_1_2,
  input  [15:0] io_mat1_1_3,
  input  [15:0] io_mat1_1_4,
  input  [15:0] io_mat1_1_5,
  input  [15:0] io_mat1_1_6,
  input  [15:0] io_mat1_1_7,
  input  [15:0] io_mat1_2_0,
  input  [15:0] io_mat1_2_1,
  input  [15:0] io_mat1_2_2,
  input  [15:0] io_mat1_2_3,
  input  [15:0] io_mat1_2_4,
  input  [15:0] io_mat1_2_5,
  input  [15:0] io_mat1_2_6,
  input  [15:0] io_mat1_2_7,
  input  [15:0] io_mat1_3_0,
  input  [15:0] io_mat1_3_1,
  input  [15:0] io_mat1_3_2,
  input  [15:0] io_mat1_3_3,
  input  [15:0] io_mat1_3_4,
  input  [15:0] io_mat1_3_5,
  input  [15:0] io_mat1_3_6,
  input  [15:0] io_mat1_3_7,
  input  [15:0] io_mat1_4_0,
  input  [15:0] io_mat1_4_1,
  input  [15:0] io_mat1_4_2,
  input  [15:0] io_mat1_4_3,
  input  [15:0] io_mat1_4_4,
  input  [15:0] io_mat1_4_5,
  input  [15:0] io_mat1_4_6,
  input  [15:0] io_mat1_4_7,
  input  [15:0] io_mat1_5_0,
  input  [15:0] io_mat1_5_1,
  input  [15:0] io_mat1_5_2,
  input  [15:0] io_mat1_5_3,
  input  [15:0] io_mat1_5_4,
  input  [15:0] io_mat1_5_5,
  input  [15:0] io_mat1_5_6,
  input  [15:0] io_mat1_5_7,
  input  [15:0] io_mat1_6_0,
  input  [15:0] io_mat1_6_1,
  input  [15:0] io_mat1_6_2,
  input  [15:0] io_mat1_6_3,
  input  [15:0] io_mat1_6_4,
  input  [15:0] io_mat1_6_5,
  input  [15:0] io_mat1_6_6,
  input  [15:0] io_mat1_6_7,
  input  [15:0] io_mat1_7_0,
  input  [15:0] io_mat1_7_1,
  input  [15:0] io_mat1_7_2,
  input  [15:0] io_mat1_7_3,
  input  [15:0] io_mat1_7_4,
  input  [15:0] io_mat1_7_5,
  input  [15:0] io_mat1_7_6,
  input  [15:0] io_mat1_7_7,
  input  [15:0] io_mat2_0_0,
  input  [15:0] io_mat2_0_1,
  input  [15:0] io_mat2_0_2,
  input  [15:0] io_mat2_0_3,
  input  [15:0] io_mat2_0_4,
  input  [15:0] io_mat2_0_5,
  input  [15:0] io_mat2_0_6,
  input  [15:0] io_mat2_0_7,
  input  [15:0] io_mat2_1_0,
  input  [15:0] io_mat2_1_1,
  input  [15:0] io_mat2_1_2,
  input  [15:0] io_mat2_1_3,
  input  [15:0] io_mat2_1_4,
  input  [15:0] io_mat2_1_5,
  input  [15:0] io_mat2_1_6,
  input  [15:0] io_mat2_1_7,
  input  [15:0] io_mat2_2_0,
  input  [15:0] io_mat2_2_1,
  input  [15:0] io_mat2_2_2,
  input  [15:0] io_mat2_2_3,
  input  [15:0] io_mat2_2_4,
  input  [15:0] io_mat2_2_5,
  input  [15:0] io_mat2_2_6,
  input  [15:0] io_mat2_2_7,
  input  [15:0] io_mat2_3_0,
  input  [15:0] io_mat2_3_1,
  input  [15:0] io_mat2_3_2,
  input  [15:0] io_mat2_3_3,
  input  [15:0] io_mat2_3_4,
  input  [15:0] io_mat2_3_5,
  input  [15:0] io_mat2_3_6,
  input  [15:0] io_mat2_3_7,
  input  [15:0] io_mat2_4_0,
  input  [15:0] io_mat2_4_1,
  input  [15:0] io_mat2_4_2,
  input  [15:0] io_mat2_4_3,
  input  [15:0] io_mat2_4_4,
  input  [15:0] io_mat2_4_5,
  input  [15:0] io_mat2_4_6,
  input  [15:0] io_mat2_4_7,
  input  [15:0] io_mat2_5_0,
  input  [15:0] io_mat2_5_1,
  input  [15:0] io_mat2_5_2,
  input  [15:0] io_mat2_5_3,
  input  [15:0] io_mat2_5_4,
  input  [15:0] io_mat2_5_5,
  input  [15:0] io_mat2_5_6,
  input  [15:0] io_mat2_5_7,
  input  [15:0] io_mat2_6_0,
  input  [15:0] io_mat2_6_1,
  input  [15:0] io_mat2_6_2,
  input  [15:0] io_mat2_6_3,
  input  [15:0] io_mat2_6_4,
  input  [15:0] io_mat2_6_5,
  input  [15:0] io_mat2_6_6,
  input  [15:0] io_mat2_6_7,
  input  [15:0] io_mat2_7_0,
  input  [15:0] io_mat2_7_1,
  input  [15:0] io_mat2_7_2,
  input  [15:0] io_mat2_7_3,
  input  [15:0] io_mat2_7_4,
  input  [15:0] io_mat2_7_5,
  input  [15:0] io_mat2_7_6,
  input  [15:0] io_mat2_7_7,
  output [15:0] io_compressedBitmap_0_0,
  output [15:0] io_compressedBitmap_0_1,
  output [15:0] io_compressedBitmap_0_2,
  output [15:0] io_compressedBitmap_0_3,
  output [15:0] io_compressedBitmap_0_4,
  output [15:0] io_compressedBitmap_0_5,
  output [15:0] io_compressedBitmap_0_6,
  output [15:0] io_compressedBitmap_0_7,
  output [15:0] io_compressedBitmap_1_0,
  output [15:0] io_compressedBitmap_1_1,
  output [15:0] io_compressedBitmap_1_2,
  output [15:0] io_compressedBitmap_1_3,
  output [15:0] io_compressedBitmap_1_4,
  output [15:0] io_compressedBitmap_1_5,
  output [15:0] io_compressedBitmap_1_6,
  output [15:0] io_compressedBitmap_1_7,
  output [15:0] io_compressedBitmap_2_0,
  output [15:0] io_compressedBitmap_2_1,
  output [15:0] io_compressedBitmap_2_2,
  output [15:0] io_compressedBitmap_2_3,
  output [15:0] io_compressedBitmap_2_4,
  output [15:0] io_compressedBitmap_2_5,
  output [15:0] io_compressedBitmap_2_6,
  output [15:0] io_compressedBitmap_2_7,
  output [15:0] io_compressedBitmap_3_0,
  output [15:0] io_compressedBitmap_3_1,
  output [15:0] io_compressedBitmap_3_2,
  output [15:0] io_compressedBitmap_3_3,
  output [15:0] io_compressedBitmap_3_4,
  output [15:0] io_compressedBitmap_3_5,
  output [15:0] io_compressedBitmap_3_6,
  output [15:0] io_compressedBitmap_3_7,
  output [15:0] io_compressedBitmap_4_0,
  output [15:0] io_compressedBitmap_4_1,
  output [15:0] io_compressedBitmap_4_2,
  output [15:0] io_compressedBitmap_4_3,
  output [15:0] io_compressedBitmap_4_4,
  output [15:0] io_compressedBitmap_4_5,
  output [15:0] io_compressedBitmap_4_6,
  output [15:0] io_compressedBitmap_4_7,
  output [15:0] io_compressedBitmap_5_0,
  output [15:0] io_compressedBitmap_5_1,
  output [15:0] io_compressedBitmap_5_2,
  output [15:0] io_compressedBitmap_5_3,
  output [15:0] io_compressedBitmap_5_4,
  output [15:0] io_compressedBitmap_5_5,
  output [15:0] io_compressedBitmap_5_6,
  output [15:0] io_compressedBitmap_5_7,
  output [15:0] io_compressedBitmap_6_0,
  output [15:0] io_compressedBitmap_6_1,
  output [15:0] io_compressedBitmap_6_2,
  output [15:0] io_compressedBitmap_6_3,
  output [15:0] io_compressedBitmap_6_4,
  output [15:0] io_compressedBitmap_6_5,
  output [15:0] io_compressedBitmap_6_6,
  output [15:0] io_compressedBitmap_6_7,
  output [15:0] io_compressedBitmap_7_0,
  output [15:0] io_compressedBitmap_7_1,
  output [15:0] io_compressedBitmap_7_2,
  output [15:0] io_compressedBitmap_7_3,
  output [15:0] io_compressedBitmap_7_4,
  output [15:0] io_compressedBitmap_7_5,
  output [15:0] io_compressedBitmap_7_6,
  output [15:0] io_compressedBitmap_7_7
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
`endif // RANDOMIZE_REG_INIT
  wire  bitmap_clock; // @[MatrixPRE-Processor.scala 17:24]
  wire  bitmap_reset; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_0_0; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_0_1; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_0_2; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_0_3; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_0_4; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_0_5; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_0_6; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_0_7; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_1_0; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_1_1; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_1_2; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_1_3; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_1_4; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_1_5; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_1_6; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_1_7; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_2_0; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_2_1; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_2_2; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_2_3; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_2_4; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_2_5; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_2_6; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_2_7; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_3_0; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_3_1; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_3_2; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_3_3; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_3_4; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_3_5; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_3_6; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_3_7; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_4_0; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_4_1; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_4_2; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_4_3; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_4_4; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_4_5; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_4_6; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_4_7; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_5_0; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_5_1; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_5_2; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_5_3; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_5_4; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_5_5; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_5_6; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_5_7; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_6_0; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_6_1; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_6_2; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_6_3; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_6_4; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_6_5; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_6_6; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_6_7; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_7_0; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_7_1; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_7_2; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_7_3; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_7_4; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_7_5; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_7_6; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_mat1_7_7; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_0_0; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_0_1; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_0_2; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_0_3; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_0_4; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_0_5; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_0_6; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_0_7; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_1_0; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_1_1; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_1_2; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_1_3; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_1_4; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_1_5; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_1_6; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_1_7; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_2_0; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_2_1; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_2_2; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_2_3; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_2_4; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_2_5; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_2_6; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_2_7; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_3_0; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_3_1; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_3_2; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_3_3; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_3_4; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_3_5; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_3_6; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_3_7; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_4_0; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_4_1; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_4_2; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_4_3; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_4_4; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_4_5; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_4_6; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_4_7; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_5_0; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_5_1; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_5_2; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_5_3; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_5_4; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_5_5; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_5_6; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_5_7; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_6_0; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_6_1; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_6_2; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_6_3; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_6_4; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_6_5; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_6_6; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_6_7; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_7_0; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_7_1; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_7_2; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_7_3; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_7_4; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_7_5; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_7_6; // @[MatrixPRE-Processor.scala 17:24]
  wire [15:0] bitmap_io_bitmap1_7_7; // @[MatrixPRE-Processor.scala 17:24]
  reg [15:0] matReg1_0_0; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_0_1; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_0_2; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_0_3; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_0_4; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_0_5; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_0_6; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_0_7; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_1_0; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_1_1; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_1_2; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_1_3; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_1_4; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_1_5; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_1_6; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_1_7; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_2_0; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_2_1; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_2_2; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_2_3; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_2_4; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_2_5; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_2_6; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_2_7; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_3_0; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_3_1; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_3_2; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_3_3; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_3_4; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_3_5; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_3_6; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_3_7; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_4_0; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_4_1; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_4_2; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_4_3; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_4_4; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_4_5; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_4_6; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_4_7; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_5_0; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_5_1; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_5_2; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_5_3; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_5_4; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_5_5; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_5_6; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_5_7; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_6_0; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_6_1; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_6_2; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_6_3; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_6_4; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_6_5; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_6_6; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_6_7; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_7_0; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_7_1; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_7_2; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_7_3; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_7_4; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_7_5; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_7_6; // @[MatrixPRE-Processor.scala 14:26]
  reg [15:0] matReg1_7_7; // @[MatrixPRE-Processor.scala 14:26]
  reg  reg_0; // @[MatrixPRE-Processor.scala 21:22]
  reg  reg_1; // @[MatrixPRE-Processor.scala 21:22]
  reg  reg_2; // @[MatrixPRE-Processor.scala 21:22]
  reg  reg_3; // @[MatrixPRE-Processor.scala 21:22]
  reg  reg_4; // @[MatrixPRE-Processor.scala 21:22]
  reg  reg_5; // @[MatrixPRE-Processor.scala 21:22]
  reg  reg_6; // @[MatrixPRE-Processor.scala 21:22]
  reg  reg_7; // @[MatrixPRE-Processor.scala 21:22]
  reg [2:0] i; // @[MatrixPRE-Processor.scala 28:20]
  reg [2:0] j; // @[MatrixPRE-Processor.scala 29:20]
  wire  _GEN_1 = 3'h1 == j ? reg_1 : reg_0; // @[MatrixPRE-Processor.scala 35:{23,23}]
  wire  _GEN_2 = 3'h2 == j ? reg_2 : _GEN_1; // @[MatrixPRE-Processor.scala 35:{23,23}]
  wire  _GEN_3 = 3'h3 == j ? reg_3 : _GEN_2; // @[MatrixPRE-Processor.scala 35:{23,23}]
  wire  _GEN_4 = 3'h4 == j ? reg_4 : _GEN_3; // @[MatrixPRE-Processor.scala 35:{23,23}]
  wire  _GEN_5 = 3'h5 == j ? reg_5 : _GEN_4; // @[MatrixPRE-Processor.scala 35:{23,23}]
  wire  _GEN_6 = 3'h6 == j ? reg_6 : _GEN_5; // @[MatrixPRE-Processor.scala 35:{23,23}]
  wire  _GEN_7 = 3'h7 == j ? reg_7 : _GEN_6; // @[MatrixPRE-Processor.scala 35:{23,23}]
  wire [15:0] _GEN_8 = bitmap_io_bitmap1_0_0; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire  _GEN_394 = 3'h0 == i; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire  _GEN_395 = 3'h1 == j; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_9 = 3'h0 == i & 3'h1 == j ? bitmap_io_bitmap1_0_1 : _GEN_8; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire  _GEN_397 = 3'h2 == j; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_10 = 3'h0 == i & 3'h2 == j ? bitmap_io_bitmap1_0_2 : _GEN_9; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire  _GEN_399 = 3'h3 == j; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_11 = 3'h0 == i & 3'h3 == j ? bitmap_io_bitmap1_0_3 : _GEN_10; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire  _GEN_401 = 3'h4 == j; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_12 = 3'h0 == i & 3'h4 == j ? bitmap_io_bitmap1_0_4 : _GEN_11; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire  _GEN_403 = 3'h5 == j; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_13 = 3'h0 == i & 3'h5 == j ? bitmap_io_bitmap1_0_5 : _GEN_12; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire  _GEN_405 = 3'h6 == j; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_14 = 3'h0 == i & 3'h6 == j ? bitmap_io_bitmap1_0_6 : _GEN_13; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire  _GEN_407 = 3'h7 == j; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_15 = 3'h0 == i & 3'h7 == j ? bitmap_io_bitmap1_0_7 : _GEN_14; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire  _GEN_408 = 3'h1 == i; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire  _GEN_409 = 3'h0 == j; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_16 = 3'h1 == i & 3'h0 == j ? bitmap_io_bitmap1_1_0 : _GEN_15; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_17 = 3'h1 == i & 3'h1 == j ? bitmap_io_bitmap1_1_1 : _GEN_16; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_18 = 3'h1 == i & 3'h2 == j ? bitmap_io_bitmap1_1_2 : _GEN_17; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_19 = 3'h1 == i & 3'h3 == j ? bitmap_io_bitmap1_1_3 : _GEN_18; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_20 = 3'h1 == i & 3'h4 == j ? bitmap_io_bitmap1_1_4 : _GEN_19; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_21 = 3'h1 == i & 3'h5 == j ? bitmap_io_bitmap1_1_5 : _GEN_20; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_22 = 3'h1 == i & 3'h6 == j ? bitmap_io_bitmap1_1_6 : _GEN_21; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_23 = 3'h1 == i & 3'h7 == j ? bitmap_io_bitmap1_1_7 : _GEN_22; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire  _GEN_424 = 3'h2 == i; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_24 = 3'h2 == i & 3'h0 == j ? bitmap_io_bitmap1_2_0 : _GEN_23; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_25 = 3'h2 == i & 3'h1 == j ? bitmap_io_bitmap1_2_1 : _GEN_24; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_26 = 3'h2 == i & 3'h2 == j ? bitmap_io_bitmap1_2_2 : _GEN_25; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_27 = 3'h2 == i & 3'h3 == j ? bitmap_io_bitmap1_2_3 : _GEN_26; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_28 = 3'h2 == i & 3'h4 == j ? bitmap_io_bitmap1_2_4 : _GEN_27; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_29 = 3'h2 == i & 3'h5 == j ? bitmap_io_bitmap1_2_5 : _GEN_28; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_30 = 3'h2 == i & 3'h6 == j ? bitmap_io_bitmap1_2_6 : _GEN_29; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_31 = 3'h2 == i & 3'h7 == j ? bitmap_io_bitmap1_2_7 : _GEN_30; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire  _GEN_440 = 3'h3 == i; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_32 = 3'h3 == i & 3'h0 == j ? bitmap_io_bitmap1_3_0 : _GEN_31; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_33 = 3'h3 == i & 3'h1 == j ? bitmap_io_bitmap1_3_1 : _GEN_32; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_34 = 3'h3 == i & 3'h2 == j ? bitmap_io_bitmap1_3_2 : _GEN_33; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_35 = 3'h3 == i & 3'h3 == j ? bitmap_io_bitmap1_3_3 : _GEN_34; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_36 = 3'h3 == i & 3'h4 == j ? bitmap_io_bitmap1_3_4 : _GEN_35; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_37 = 3'h3 == i & 3'h5 == j ? bitmap_io_bitmap1_3_5 : _GEN_36; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_38 = 3'h3 == i & 3'h6 == j ? bitmap_io_bitmap1_3_6 : _GEN_37; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_39 = 3'h3 == i & 3'h7 == j ? bitmap_io_bitmap1_3_7 : _GEN_38; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire  _GEN_456 = 3'h4 == i; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_40 = 3'h4 == i & 3'h0 == j ? bitmap_io_bitmap1_4_0 : _GEN_39; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_41 = 3'h4 == i & 3'h1 == j ? bitmap_io_bitmap1_4_1 : _GEN_40; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_42 = 3'h4 == i & 3'h2 == j ? bitmap_io_bitmap1_4_2 : _GEN_41; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_43 = 3'h4 == i & 3'h3 == j ? bitmap_io_bitmap1_4_3 : _GEN_42; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_44 = 3'h4 == i & 3'h4 == j ? bitmap_io_bitmap1_4_4 : _GEN_43; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_45 = 3'h4 == i & 3'h5 == j ? bitmap_io_bitmap1_4_5 : _GEN_44; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_46 = 3'h4 == i & 3'h6 == j ? bitmap_io_bitmap1_4_6 : _GEN_45; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_47 = 3'h4 == i & 3'h7 == j ? bitmap_io_bitmap1_4_7 : _GEN_46; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire  _GEN_472 = 3'h5 == i; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_48 = 3'h5 == i & 3'h0 == j ? bitmap_io_bitmap1_5_0 : _GEN_47; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_49 = 3'h5 == i & 3'h1 == j ? bitmap_io_bitmap1_5_1 : _GEN_48; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_50 = 3'h5 == i & 3'h2 == j ? bitmap_io_bitmap1_5_2 : _GEN_49; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_51 = 3'h5 == i & 3'h3 == j ? bitmap_io_bitmap1_5_3 : _GEN_50; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_52 = 3'h5 == i & 3'h4 == j ? bitmap_io_bitmap1_5_4 : _GEN_51; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_53 = 3'h5 == i & 3'h5 == j ? bitmap_io_bitmap1_5_5 : _GEN_52; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_54 = 3'h5 == i & 3'h6 == j ? bitmap_io_bitmap1_5_6 : _GEN_53; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_55 = 3'h5 == i & 3'h7 == j ? bitmap_io_bitmap1_5_7 : _GEN_54; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire  _GEN_488 = 3'h6 == i; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_56 = 3'h6 == i & 3'h0 == j ? bitmap_io_bitmap1_6_0 : _GEN_55; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_57 = 3'h6 == i & 3'h1 == j ? bitmap_io_bitmap1_6_1 : _GEN_56; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_58 = 3'h6 == i & 3'h2 == j ? bitmap_io_bitmap1_6_2 : _GEN_57; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_59 = 3'h6 == i & 3'h3 == j ? bitmap_io_bitmap1_6_3 : _GEN_58; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_60 = 3'h6 == i & 3'h4 == j ? bitmap_io_bitmap1_6_4 : _GEN_59; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_61 = 3'h6 == i & 3'h5 == j ? bitmap_io_bitmap1_6_5 : _GEN_60; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_62 = 3'h6 == i & 3'h6 == j ? bitmap_io_bitmap1_6_6 : _GEN_61; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_63 = 3'h6 == i & 3'h7 == j ? bitmap_io_bitmap1_6_7 : _GEN_62; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire  _GEN_504 = 3'h7 == i; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_64 = 3'h7 == i & 3'h0 == j ? bitmap_io_bitmap1_7_0 : _GEN_63; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_65 = 3'h7 == i & 3'h1 == j ? bitmap_io_bitmap1_7_1 : _GEN_64; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_66 = 3'h7 == i & 3'h2 == j ? bitmap_io_bitmap1_7_2 : _GEN_65; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_67 = 3'h7 == i & 3'h3 == j ? bitmap_io_bitmap1_7_3 : _GEN_66; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_68 = 3'h7 == i & 3'h4 == j ? bitmap_io_bitmap1_7_4 : _GEN_67; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_69 = 3'h7 == i & 3'h5 == j ? bitmap_io_bitmap1_7_5 : _GEN_68; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_70 = 3'h7 == i & 3'h6 == j ? bitmap_io_bitmap1_7_6 : _GEN_69; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_71 = 3'h7 == i & 3'h7 == j ? bitmap_io_bitmap1_7_7 : _GEN_70; // @[MatrixPRE-Processor.scala 35:{60,60}]
  wire [15:0] _GEN_201 = _GEN_394 & _GEN_395 ? io_mat1_0_1 : io_mat1_0_0; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_202 = _GEN_394 & _GEN_397 ? io_mat1_0_2 : _GEN_201; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_203 = _GEN_394 & _GEN_399 ? io_mat1_0_3 : _GEN_202; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_204 = _GEN_394 & _GEN_401 ? io_mat1_0_4 : _GEN_203; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_205 = _GEN_394 & _GEN_403 ? io_mat1_0_5 : _GEN_204; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_206 = _GEN_394 & _GEN_405 ? io_mat1_0_6 : _GEN_205; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_207 = _GEN_394 & _GEN_407 ? io_mat1_0_7 : _GEN_206; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_208 = _GEN_408 & _GEN_409 ? io_mat1_1_0 : _GEN_207; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_209 = _GEN_408 & _GEN_395 ? io_mat1_1_1 : _GEN_208; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_210 = _GEN_408 & _GEN_397 ? io_mat1_1_2 : _GEN_209; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_211 = _GEN_408 & _GEN_399 ? io_mat1_1_3 : _GEN_210; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_212 = _GEN_408 & _GEN_401 ? io_mat1_1_4 : _GEN_211; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_213 = _GEN_408 & _GEN_403 ? io_mat1_1_5 : _GEN_212; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_214 = _GEN_408 & _GEN_405 ? io_mat1_1_6 : _GEN_213; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_215 = _GEN_408 & _GEN_407 ? io_mat1_1_7 : _GEN_214; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_216 = _GEN_424 & _GEN_409 ? io_mat1_2_0 : _GEN_215; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_217 = _GEN_424 & _GEN_395 ? io_mat1_2_1 : _GEN_216; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_218 = _GEN_424 & _GEN_397 ? io_mat1_2_2 : _GEN_217; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_219 = _GEN_424 & _GEN_399 ? io_mat1_2_3 : _GEN_218; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_220 = _GEN_424 & _GEN_401 ? io_mat1_2_4 : _GEN_219; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_221 = _GEN_424 & _GEN_403 ? io_mat1_2_5 : _GEN_220; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_222 = _GEN_424 & _GEN_405 ? io_mat1_2_6 : _GEN_221; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_223 = _GEN_424 & _GEN_407 ? io_mat1_2_7 : _GEN_222; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_224 = _GEN_440 & _GEN_409 ? io_mat1_3_0 : _GEN_223; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_225 = _GEN_440 & _GEN_395 ? io_mat1_3_1 : _GEN_224; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_226 = _GEN_440 & _GEN_397 ? io_mat1_3_2 : _GEN_225; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_227 = _GEN_440 & _GEN_399 ? io_mat1_3_3 : _GEN_226; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_228 = _GEN_440 & _GEN_401 ? io_mat1_3_4 : _GEN_227; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_229 = _GEN_440 & _GEN_403 ? io_mat1_3_5 : _GEN_228; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_230 = _GEN_440 & _GEN_405 ? io_mat1_3_6 : _GEN_229; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_231 = _GEN_440 & _GEN_407 ? io_mat1_3_7 : _GEN_230; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_232 = _GEN_456 & _GEN_409 ? io_mat1_4_0 : _GEN_231; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_233 = _GEN_456 & _GEN_395 ? io_mat1_4_1 : _GEN_232; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_234 = _GEN_456 & _GEN_397 ? io_mat1_4_2 : _GEN_233; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_235 = _GEN_456 & _GEN_399 ? io_mat1_4_3 : _GEN_234; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_236 = _GEN_456 & _GEN_401 ? io_mat1_4_4 : _GEN_235; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_237 = _GEN_456 & _GEN_403 ? io_mat1_4_5 : _GEN_236; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_238 = _GEN_456 & _GEN_405 ? io_mat1_4_6 : _GEN_237; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_239 = _GEN_456 & _GEN_407 ? io_mat1_4_7 : _GEN_238; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_240 = _GEN_472 & _GEN_409 ? io_mat1_5_0 : _GEN_239; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_241 = _GEN_472 & _GEN_395 ? io_mat1_5_1 : _GEN_240; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_242 = _GEN_472 & _GEN_397 ? io_mat1_5_2 : _GEN_241; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_243 = _GEN_472 & _GEN_399 ? io_mat1_5_3 : _GEN_242; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_244 = _GEN_472 & _GEN_401 ? io_mat1_5_4 : _GEN_243; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_245 = _GEN_472 & _GEN_403 ? io_mat1_5_5 : _GEN_244; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_246 = _GEN_472 & _GEN_405 ? io_mat1_5_6 : _GEN_245; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_247 = _GEN_472 & _GEN_407 ? io_mat1_5_7 : _GEN_246; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_248 = _GEN_488 & _GEN_409 ? io_mat1_6_0 : _GEN_247; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_249 = _GEN_488 & _GEN_395 ? io_mat1_6_1 : _GEN_248; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_250 = _GEN_488 & _GEN_397 ? io_mat1_6_2 : _GEN_249; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_251 = _GEN_488 & _GEN_399 ? io_mat1_6_3 : _GEN_250; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_252 = _GEN_488 & _GEN_401 ? io_mat1_6_4 : _GEN_251; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_253 = _GEN_488 & _GEN_403 ? io_mat1_6_5 : _GEN_252; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_254 = _GEN_488 & _GEN_405 ? io_mat1_6_6 : _GEN_253; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_255 = _GEN_488 & _GEN_407 ? io_mat1_6_7 : _GEN_254; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_256 = _GEN_504 & _GEN_409 ? io_mat1_7_0 : _GEN_255; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_257 = _GEN_504 & _GEN_395 ? io_mat1_7_1 : _GEN_256; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_258 = _GEN_504 & _GEN_397 ? io_mat1_7_2 : _GEN_257; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_259 = _GEN_504 & _GEN_399 ? io_mat1_7_3 : _GEN_258; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_260 = _GEN_504 & _GEN_401 ? io_mat1_7_4 : _GEN_259; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_261 = _GEN_504 & _GEN_403 ? io_mat1_7_5 : _GEN_260; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [15:0] _GEN_262 = _GEN_504 & _GEN_405 ? io_mat1_7_6 : _GEN_261; // @[MatrixPRE-Processor.scala 38:{27,27}]
  wire [2:0] _i_T_1 = i + 3'h1; // @[MatrixPRE-Processor.scala 40:16]
  wire [2:0] _j_T_1 = j + 3'h1; // @[MatrixPRE-Processor.scala 43:16]
  Bitmap bitmap ( // @[MatrixPRE-Processor.scala 17:24]
    .clock(bitmap_clock),
    .reset(bitmap_reset),
    .io_mat1_0_0(bitmap_io_mat1_0_0),
    .io_mat1_0_1(bitmap_io_mat1_0_1),
    .io_mat1_0_2(bitmap_io_mat1_0_2),
    .io_mat1_0_3(bitmap_io_mat1_0_3),
    .io_mat1_0_4(bitmap_io_mat1_0_4),
    .io_mat1_0_5(bitmap_io_mat1_0_5),
    .io_mat1_0_6(bitmap_io_mat1_0_6),
    .io_mat1_0_7(bitmap_io_mat1_0_7),
    .io_mat1_1_0(bitmap_io_mat1_1_0),
    .io_mat1_1_1(bitmap_io_mat1_1_1),
    .io_mat1_1_2(bitmap_io_mat1_1_2),
    .io_mat1_1_3(bitmap_io_mat1_1_3),
    .io_mat1_1_4(bitmap_io_mat1_1_4),
    .io_mat1_1_5(bitmap_io_mat1_1_5),
    .io_mat1_1_6(bitmap_io_mat1_1_6),
    .io_mat1_1_7(bitmap_io_mat1_1_7),
    .io_mat1_2_0(bitmap_io_mat1_2_0),
    .io_mat1_2_1(bitmap_io_mat1_2_1),
    .io_mat1_2_2(bitmap_io_mat1_2_2),
    .io_mat1_2_3(bitmap_io_mat1_2_3),
    .io_mat1_2_4(bitmap_io_mat1_2_4),
    .io_mat1_2_5(bitmap_io_mat1_2_5),
    .io_mat1_2_6(bitmap_io_mat1_2_6),
    .io_mat1_2_7(bitmap_io_mat1_2_7),
    .io_mat1_3_0(bitmap_io_mat1_3_0),
    .io_mat1_3_1(bitmap_io_mat1_3_1),
    .io_mat1_3_2(bitmap_io_mat1_3_2),
    .io_mat1_3_3(bitmap_io_mat1_3_3),
    .io_mat1_3_4(bitmap_io_mat1_3_4),
    .io_mat1_3_5(bitmap_io_mat1_3_5),
    .io_mat1_3_6(bitmap_io_mat1_3_6),
    .io_mat1_3_7(bitmap_io_mat1_3_7),
    .io_mat1_4_0(bitmap_io_mat1_4_0),
    .io_mat1_4_1(bitmap_io_mat1_4_1),
    .io_mat1_4_2(bitmap_io_mat1_4_2),
    .io_mat1_4_3(bitmap_io_mat1_4_3),
    .io_mat1_4_4(bitmap_io_mat1_4_4),
    .io_mat1_4_5(bitmap_io_mat1_4_5),
    .io_mat1_4_6(bitmap_io_mat1_4_6),
    .io_mat1_4_7(bitmap_io_mat1_4_7),
    .io_mat1_5_0(bitmap_io_mat1_5_0),
    .io_mat1_5_1(bitmap_io_mat1_5_1),
    .io_mat1_5_2(bitmap_io_mat1_5_2),
    .io_mat1_5_3(bitmap_io_mat1_5_3),
    .io_mat1_5_4(bitmap_io_mat1_5_4),
    .io_mat1_5_5(bitmap_io_mat1_5_5),
    .io_mat1_5_6(bitmap_io_mat1_5_6),
    .io_mat1_5_7(bitmap_io_mat1_5_7),
    .io_mat1_6_0(bitmap_io_mat1_6_0),
    .io_mat1_6_1(bitmap_io_mat1_6_1),
    .io_mat1_6_2(bitmap_io_mat1_6_2),
    .io_mat1_6_3(bitmap_io_mat1_6_3),
    .io_mat1_6_4(bitmap_io_mat1_6_4),
    .io_mat1_6_5(bitmap_io_mat1_6_5),
    .io_mat1_6_6(bitmap_io_mat1_6_6),
    .io_mat1_6_7(bitmap_io_mat1_6_7),
    .io_mat1_7_0(bitmap_io_mat1_7_0),
    .io_mat1_7_1(bitmap_io_mat1_7_1),
    .io_mat1_7_2(bitmap_io_mat1_7_2),
    .io_mat1_7_3(bitmap_io_mat1_7_3),
    .io_mat1_7_4(bitmap_io_mat1_7_4),
    .io_mat1_7_5(bitmap_io_mat1_7_5),
    .io_mat1_7_6(bitmap_io_mat1_7_6),
    .io_mat1_7_7(bitmap_io_mat1_7_7),
    .io_bitmap1_0_0(bitmap_io_bitmap1_0_0),
    .io_bitmap1_0_1(bitmap_io_bitmap1_0_1),
    .io_bitmap1_0_2(bitmap_io_bitmap1_0_2),
    .io_bitmap1_0_3(bitmap_io_bitmap1_0_3),
    .io_bitmap1_0_4(bitmap_io_bitmap1_0_4),
    .io_bitmap1_0_5(bitmap_io_bitmap1_0_5),
    .io_bitmap1_0_6(bitmap_io_bitmap1_0_6),
    .io_bitmap1_0_7(bitmap_io_bitmap1_0_7),
    .io_bitmap1_1_0(bitmap_io_bitmap1_1_0),
    .io_bitmap1_1_1(bitmap_io_bitmap1_1_1),
    .io_bitmap1_1_2(bitmap_io_bitmap1_1_2),
    .io_bitmap1_1_3(bitmap_io_bitmap1_1_3),
    .io_bitmap1_1_4(bitmap_io_bitmap1_1_4),
    .io_bitmap1_1_5(bitmap_io_bitmap1_1_5),
    .io_bitmap1_1_6(bitmap_io_bitmap1_1_6),
    .io_bitmap1_1_7(bitmap_io_bitmap1_1_7),
    .io_bitmap1_2_0(bitmap_io_bitmap1_2_0),
    .io_bitmap1_2_1(bitmap_io_bitmap1_2_1),
    .io_bitmap1_2_2(bitmap_io_bitmap1_2_2),
    .io_bitmap1_2_3(bitmap_io_bitmap1_2_3),
    .io_bitmap1_2_4(bitmap_io_bitmap1_2_4),
    .io_bitmap1_2_5(bitmap_io_bitmap1_2_5),
    .io_bitmap1_2_6(bitmap_io_bitmap1_2_6),
    .io_bitmap1_2_7(bitmap_io_bitmap1_2_7),
    .io_bitmap1_3_0(bitmap_io_bitmap1_3_0),
    .io_bitmap1_3_1(bitmap_io_bitmap1_3_1),
    .io_bitmap1_3_2(bitmap_io_bitmap1_3_2),
    .io_bitmap1_3_3(bitmap_io_bitmap1_3_3),
    .io_bitmap1_3_4(bitmap_io_bitmap1_3_4),
    .io_bitmap1_3_5(bitmap_io_bitmap1_3_5),
    .io_bitmap1_3_6(bitmap_io_bitmap1_3_6),
    .io_bitmap1_3_7(bitmap_io_bitmap1_3_7),
    .io_bitmap1_4_0(bitmap_io_bitmap1_4_0),
    .io_bitmap1_4_1(bitmap_io_bitmap1_4_1),
    .io_bitmap1_4_2(bitmap_io_bitmap1_4_2),
    .io_bitmap1_4_3(bitmap_io_bitmap1_4_3),
    .io_bitmap1_4_4(bitmap_io_bitmap1_4_4),
    .io_bitmap1_4_5(bitmap_io_bitmap1_4_5),
    .io_bitmap1_4_6(bitmap_io_bitmap1_4_6),
    .io_bitmap1_4_7(bitmap_io_bitmap1_4_7),
    .io_bitmap1_5_0(bitmap_io_bitmap1_5_0),
    .io_bitmap1_5_1(bitmap_io_bitmap1_5_1),
    .io_bitmap1_5_2(bitmap_io_bitmap1_5_2),
    .io_bitmap1_5_3(bitmap_io_bitmap1_5_3),
    .io_bitmap1_5_4(bitmap_io_bitmap1_5_4),
    .io_bitmap1_5_5(bitmap_io_bitmap1_5_5),
    .io_bitmap1_5_6(bitmap_io_bitmap1_5_6),
    .io_bitmap1_5_7(bitmap_io_bitmap1_5_7),
    .io_bitmap1_6_0(bitmap_io_bitmap1_6_0),
    .io_bitmap1_6_1(bitmap_io_bitmap1_6_1),
    .io_bitmap1_6_2(bitmap_io_bitmap1_6_2),
    .io_bitmap1_6_3(bitmap_io_bitmap1_6_3),
    .io_bitmap1_6_4(bitmap_io_bitmap1_6_4),
    .io_bitmap1_6_5(bitmap_io_bitmap1_6_5),
    .io_bitmap1_6_6(bitmap_io_bitmap1_6_6),
    .io_bitmap1_6_7(bitmap_io_bitmap1_6_7),
    .io_bitmap1_7_0(bitmap_io_bitmap1_7_0),
    .io_bitmap1_7_1(bitmap_io_bitmap1_7_1),
    .io_bitmap1_7_2(bitmap_io_bitmap1_7_2),
    .io_bitmap1_7_3(bitmap_io_bitmap1_7_3),
    .io_bitmap1_7_4(bitmap_io_bitmap1_7_4),
    .io_bitmap1_7_5(bitmap_io_bitmap1_7_5),
    .io_bitmap1_7_6(bitmap_io_bitmap1_7_6),
    .io_bitmap1_7_7(bitmap_io_bitmap1_7_7)
  );
  assign io_compressedBitmap_0_0 = matReg1_0_0; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_0_1 = matReg1_0_1; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_0_2 = matReg1_0_2; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_0_3 = matReg1_0_3; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_0_4 = matReg1_0_4; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_0_5 = matReg1_0_5; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_0_6 = matReg1_0_6; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_0_7 = matReg1_0_7; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_1_0 = matReg1_1_0; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_1_1 = matReg1_1_1; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_1_2 = matReg1_1_2; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_1_3 = matReg1_1_3; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_1_4 = matReg1_1_4; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_1_5 = matReg1_1_5; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_1_6 = matReg1_1_6; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_1_7 = matReg1_1_7; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_2_0 = matReg1_2_0; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_2_1 = matReg1_2_1; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_2_2 = matReg1_2_2; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_2_3 = matReg1_2_3; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_2_4 = matReg1_2_4; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_2_5 = matReg1_2_5; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_2_6 = matReg1_2_6; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_2_7 = matReg1_2_7; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_3_0 = matReg1_3_0; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_3_1 = matReg1_3_1; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_3_2 = matReg1_3_2; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_3_3 = matReg1_3_3; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_3_4 = matReg1_3_4; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_3_5 = matReg1_3_5; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_3_6 = matReg1_3_6; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_3_7 = matReg1_3_7; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_4_0 = matReg1_4_0; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_4_1 = matReg1_4_1; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_4_2 = matReg1_4_2; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_4_3 = matReg1_4_3; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_4_4 = matReg1_4_4; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_4_5 = matReg1_4_5; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_4_6 = matReg1_4_6; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_4_7 = matReg1_4_7; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_5_0 = matReg1_5_0; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_5_1 = matReg1_5_1; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_5_2 = matReg1_5_2; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_5_3 = matReg1_5_3; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_5_4 = matReg1_5_4; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_5_5 = matReg1_5_5; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_5_6 = matReg1_5_6; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_5_7 = matReg1_5_7; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_6_0 = matReg1_6_0; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_6_1 = matReg1_6_1; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_6_2 = matReg1_6_2; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_6_3 = matReg1_6_3; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_6_4 = matReg1_6_4; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_6_5 = matReg1_6_5; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_6_6 = matReg1_6_6; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_6_7 = matReg1_6_7; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_7_0 = matReg1_7_0; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_7_1 = matReg1_7_1; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_7_2 = matReg1_7_2; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_7_3 = matReg1_7_3; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_7_4 = matReg1_7_4; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_7_5 = matReg1_7_5; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_7_6 = matReg1_7_6; // @[MatrixPRE-Processor.scala 15:25]
  assign io_compressedBitmap_7_7 = matReg1_7_7; // @[MatrixPRE-Processor.scala 15:25]
  assign bitmap_clock = clock;
  assign bitmap_reset = reset;
  assign bitmap_io_mat1_0_0 = io_mat1_0_0; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_0_1 = io_mat1_0_1; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_0_2 = io_mat1_0_2; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_0_3 = io_mat1_0_3; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_0_4 = io_mat1_0_4; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_0_5 = io_mat1_0_5; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_0_6 = io_mat1_0_6; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_0_7 = io_mat1_0_7; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_1_0 = io_mat1_1_0; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_1_1 = io_mat1_1_1; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_1_2 = io_mat1_1_2; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_1_3 = io_mat1_1_3; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_1_4 = io_mat1_1_4; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_1_5 = io_mat1_1_5; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_1_6 = io_mat1_1_6; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_1_7 = io_mat1_1_7; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_2_0 = io_mat1_2_0; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_2_1 = io_mat1_2_1; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_2_2 = io_mat1_2_2; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_2_3 = io_mat1_2_3; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_2_4 = io_mat1_2_4; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_2_5 = io_mat1_2_5; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_2_6 = io_mat1_2_6; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_2_7 = io_mat1_2_7; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_3_0 = io_mat1_3_0; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_3_1 = io_mat1_3_1; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_3_2 = io_mat1_3_2; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_3_3 = io_mat1_3_3; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_3_4 = io_mat1_3_4; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_3_5 = io_mat1_3_5; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_3_6 = io_mat1_3_6; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_3_7 = io_mat1_3_7; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_4_0 = io_mat1_4_0; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_4_1 = io_mat1_4_1; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_4_2 = io_mat1_4_2; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_4_3 = io_mat1_4_3; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_4_4 = io_mat1_4_4; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_4_5 = io_mat1_4_5; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_4_6 = io_mat1_4_6; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_4_7 = io_mat1_4_7; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_5_0 = io_mat1_5_0; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_5_1 = io_mat1_5_1; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_5_2 = io_mat1_5_2; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_5_3 = io_mat1_5_3; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_5_4 = io_mat1_5_4; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_5_5 = io_mat1_5_5; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_5_6 = io_mat1_5_6; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_5_7 = io_mat1_5_7; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_6_0 = io_mat1_6_0; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_6_1 = io_mat1_6_1; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_6_2 = io_mat1_6_2; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_6_3 = io_mat1_6_3; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_6_4 = io_mat1_6_4; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_6_5 = io_mat1_6_5; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_6_6 = io_mat1_6_6; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_6_7 = io_mat1_6_7; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_7_0 = io_mat1_7_0; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_7_1 = io_mat1_7_1; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_7_2 = io_mat1_7_2; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_7_3 = io_mat1_7_3; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_7_4 = io_mat1_7_4; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_7_5 = io_mat1_7_5; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_7_6 = io_mat1_7_6; // @[MatrixPRE-Processor.scala 18:20]
  assign bitmap_io_mat1_7_7 = io_mat1_7_7; // @[MatrixPRE-Processor.scala 18:20]
  always @(posedge clock) begin
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_0_0 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_394 & _GEN_409) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_0_0 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_394 & _GEN_409) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_0_0 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_0_0 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_0_1 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_394 & _GEN_395) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_0_1 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_394 & _GEN_395) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_0_1 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_0_1 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_0_2 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_394 & _GEN_397) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_0_2 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_394 & _GEN_397) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_0_2 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_0_2 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_0_3 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_394 & _GEN_399) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_0_3 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_394 & _GEN_399) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_0_3 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_0_3 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_0_4 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_394 & _GEN_401) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_0_4 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_394 & _GEN_401) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_0_4 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_0_4 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_0_5 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_394 & _GEN_403) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_0_5 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_394 & _GEN_403) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_0_5 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_0_5 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_0_6 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_394 & _GEN_405) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_0_6 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_394 & _GEN_405) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_0_6 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_0_6 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_0_7 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_394 & _GEN_407) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_0_7 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_394 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_0_7 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_0_7 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_1_0 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_408 & _GEN_409) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_1_0 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_408 & _GEN_409) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_1_0 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_1_0 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_1_1 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_408 & _GEN_395) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_1_1 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_408 & _GEN_395) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_1_1 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_1_1 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_1_2 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_408 & _GEN_397) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_1_2 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_408 & _GEN_397) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_1_2 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_1_2 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_1_3 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_408 & _GEN_399) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_1_3 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_408 & _GEN_399) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_1_3 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_1_3 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_1_4 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_408 & _GEN_401) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_1_4 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_408 & _GEN_401) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_1_4 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_1_4 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_1_5 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_408 & _GEN_403) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_1_5 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_408 & _GEN_403) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_1_5 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_1_5 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_1_6 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_408 & _GEN_405) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_1_6 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_408 & _GEN_405) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_1_6 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_1_6 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_1_7 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_408 & _GEN_407) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_1_7 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_408 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_1_7 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_1_7 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_2_0 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_424 & _GEN_409) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_2_0 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_424 & _GEN_409) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_2_0 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_2_0 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_2_1 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_424 & _GEN_395) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_2_1 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_424 & _GEN_395) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_2_1 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_2_1 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_2_2 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_424 & _GEN_397) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_2_2 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_424 & _GEN_397) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_2_2 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_2_2 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_2_3 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_424 & _GEN_399) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_2_3 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_424 & _GEN_399) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_2_3 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_2_3 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_2_4 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_424 & _GEN_401) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_2_4 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_424 & _GEN_401) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_2_4 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_2_4 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_2_5 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_424 & _GEN_403) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_2_5 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_424 & _GEN_403) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_2_5 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_2_5 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_2_6 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_424 & _GEN_405) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_2_6 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_424 & _GEN_405) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_2_6 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_2_6 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_2_7 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_424 & _GEN_407) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_2_7 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_424 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_2_7 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_2_7 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_3_0 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_440 & _GEN_409) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_3_0 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_440 & _GEN_409) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_3_0 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_3_0 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_3_1 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_440 & _GEN_395) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_3_1 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_440 & _GEN_395) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_3_1 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_3_1 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_3_2 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_440 & _GEN_397) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_3_2 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_440 & _GEN_397) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_3_2 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_3_2 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_3_3 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_440 & _GEN_399) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_3_3 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_440 & _GEN_399) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_3_3 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_3_3 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_3_4 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_440 & _GEN_401) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_3_4 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_440 & _GEN_401) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_3_4 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_3_4 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_3_5 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_440 & _GEN_403) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_3_5 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_440 & _GEN_403) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_3_5 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_3_5 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_3_6 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_440 & _GEN_405) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_3_6 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_440 & _GEN_405) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_3_6 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_3_6 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_3_7 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_440 & _GEN_407) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_3_7 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_440 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_3_7 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_3_7 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_4_0 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_456 & _GEN_409) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_4_0 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_456 & _GEN_409) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_4_0 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_4_0 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_4_1 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_456 & _GEN_395) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_4_1 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_456 & _GEN_395) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_4_1 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_4_1 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_4_2 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_456 & _GEN_397) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_4_2 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_456 & _GEN_397) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_4_2 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_4_2 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_4_3 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_456 & _GEN_399) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_4_3 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_456 & _GEN_399) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_4_3 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_4_3 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_4_4 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_456 & _GEN_401) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_4_4 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_456 & _GEN_401) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_4_4 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_4_4 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_4_5 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_456 & _GEN_403) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_4_5 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_456 & _GEN_403) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_4_5 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_4_5 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_4_6 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_456 & _GEN_405) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_4_6 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_456 & _GEN_405) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_4_6 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_4_6 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_4_7 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_456 & _GEN_407) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_4_7 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_456 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_4_7 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_4_7 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_5_0 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_472 & _GEN_409) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_5_0 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_472 & _GEN_409) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_5_0 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_5_0 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_5_1 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_472 & _GEN_395) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_5_1 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_472 & _GEN_395) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_5_1 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_5_1 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_5_2 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_472 & _GEN_397) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_5_2 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_472 & _GEN_397) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_5_2 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_5_2 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_5_3 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_472 & _GEN_399) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_5_3 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_472 & _GEN_399) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_5_3 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_5_3 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_5_4 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_472 & _GEN_401) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_5_4 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_472 & _GEN_401) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_5_4 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_5_4 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_5_5 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_472 & _GEN_403) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_5_5 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_472 & _GEN_403) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_5_5 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_5_5 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_5_6 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_472 & _GEN_405) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_5_6 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_472 & _GEN_405) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_5_6 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_5_6 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_5_7 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_472 & _GEN_407) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_5_7 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_472 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_5_7 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_5_7 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_6_0 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_488 & _GEN_409) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_6_0 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_488 & _GEN_409) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_6_0 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_6_0 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_6_1 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_488 & _GEN_395) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_6_1 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_488 & _GEN_395) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_6_1 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_6_1 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_6_2 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_488 & _GEN_397) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_6_2 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_488 & _GEN_397) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_6_2 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_6_2 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_6_3 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_488 & _GEN_399) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_6_3 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_488 & _GEN_399) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_6_3 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_6_3 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_6_4 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_488 & _GEN_401) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_6_4 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_488 & _GEN_401) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_6_4 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_6_4 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_6_5 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_488 & _GEN_403) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_6_5 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_488 & _GEN_403) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_6_5 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_6_5 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_6_6 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_488 & _GEN_405) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_6_6 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_488 & _GEN_405) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_6_6 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_6_6 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_6_7 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_488 & _GEN_407) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_6_7 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_488 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_6_7 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_6_7 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_7_0 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_504 & _GEN_409) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_7_0 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_504 & _GEN_409) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_7_0 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_7_0 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_7_1 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_504 & _GEN_395) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_7_1 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_504 & _GEN_395) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_7_1 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_7_1 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_7_2 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_504 & _GEN_397) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_7_2 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_504 & _GEN_397) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_7_2 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_7_2 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_7_3 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_504 & _GEN_399) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_7_3 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_504 & _GEN_399) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_7_3 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_7_3 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_7_4 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_504 & _GEN_401) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_7_4 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_504 & _GEN_401) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_7_4 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_7_4 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_7_5 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_504 & _GEN_403) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_7_5 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_504 & _GEN_403) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_7_5 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_7_5 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_7_6 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_504 & _GEN_405) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_7_6 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_504 & _GEN_405) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_7_6 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_7_6 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 14:26]
      matReg1_7_7 <= 16'h0; // @[MatrixPRE-Processor.scala 14:26]
    end else if (~_GEN_7 & _GEN_71 == 16'h1) begin // @[MatrixPRE-Processor.scala 35:69]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 36:27]
        matReg1_7_7 <= 16'h0; // @[MatrixPRE-Processor.scala 36:27]
      end
    end else if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
      if (_GEN_504 & _GEN_407) begin // @[MatrixPRE-Processor.scala 38:27]
        matReg1_7_7 <= io_mat1_7_7; // @[MatrixPRE-Processor.scala 38:27]
      end else begin
        matReg1_7_7 <= _GEN_262;
      end
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 21:22]
      reg_0 <= 1'h0; // @[MatrixPRE-Processor.scala 21:22]
    end else begin
      reg_0 <= io_mat2_0_0 != 16'h0 | io_mat2_0_1 != 16'h0 | io_mat2_0_2 != 16'h0 | io_mat2_0_3 != 16'h0 | io_mat2_0_4
         != 16'h0 | io_mat2_0_5 != 16'h0 | io_mat2_0_6 != 16'h0 | io_mat2_0_7 != 16'h0; // @[MatrixPRE-Processor.scala 23:16]
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 21:22]
      reg_1 <= 1'h0; // @[MatrixPRE-Processor.scala 21:22]
    end else begin
      reg_1 <= io_mat2_1_0 != 16'h0 | io_mat2_1_1 != 16'h0 | io_mat2_1_2 != 16'h0 | io_mat2_1_3 != 16'h0 | io_mat2_1_4
         != 16'h0 | io_mat2_1_5 != 16'h0 | io_mat2_1_6 != 16'h0 | io_mat2_1_7 != 16'h0; // @[MatrixPRE-Processor.scala 23:16]
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 21:22]
      reg_2 <= 1'h0; // @[MatrixPRE-Processor.scala 21:22]
    end else begin
      reg_2 <= io_mat2_2_0 != 16'h0 | io_mat2_2_1 != 16'h0 | io_mat2_2_2 != 16'h0 | io_mat2_2_3 != 16'h0 | io_mat2_2_4
         != 16'h0 | io_mat2_2_5 != 16'h0 | io_mat2_2_6 != 16'h0 | io_mat2_2_7 != 16'h0; // @[MatrixPRE-Processor.scala 23:16]
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 21:22]
      reg_3 <= 1'h0; // @[MatrixPRE-Processor.scala 21:22]
    end else begin
      reg_3 <= io_mat2_3_0 != 16'h0 | io_mat2_3_1 != 16'h0 | io_mat2_3_2 != 16'h0 | io_mat2_3_3 != 16'h0 | io_mat2_3_4
         != 16'h0 | io_mat2_3_5 != 16'h0 | io_mat2_3_6 != 16'h0 | io_mat2_3_7 != 16'h0; // @[MatrixPRE-Processor.scala 23:16]
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 21:22]
      reg_4 <= 1'h0; // @[MatrixPRE-Processor.scala 21:22]
    end else begin
      reg_4 <= io_mat2_4_0 != 16'h0 | io_mat2_4_1 != 16'h0 | io_mat2_4_2 != 16'h0 | io_mat2_4_3 != 16'h0 | io_mat2_4_4
         != 16'h0 | io_mat2_4_5 != 16'h0 | io_mat2_4_6 != 16'h0 | io_mat2_4_7 != 16'h0; // @[MatrixPRE-Processor.scala 23:16]
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 21:22]
      reg_5 <= 1'h0; // @[MatrixPRE-Processor.scala 21:22]
    end else begin
      reg_5 <= io_mat2_5_0 != 16'h0 | io_mat2_5_1 != 16'h0 | io_mat2_5_2 != 16'h0 | io_mat2_5_3 != 16'h0 | io_mat2_5_4
         != 16'h0 | io_mat2_5_5 != 16'h0 | io_mat2_5_6 != 16'h0 | io_mat2_5_7 != 16'h0; // @[MatrixPRE-Processor.scala 23:16]
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 21:22]
      reg_6 <= 1'h0; // @[MatrixPRE-Processor.scala 21:22]
    end else begin
      reg_6 <= io_mat2_6_0 != 16'h0 | io_mat2_6_1 != 16'h0 | io_mat2_6_2 != 16'h0 | io_mat2_6_3 != 16'h0 | io_mat2_6_4
         != 16'h0 | io_mat2_6_5 != 16'h0 | io_mat2_6_6 != 16'h0 | io_mat2_6_7 != 16'h0; // @[MatrixPRE-Processor.scala 23:16]
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 21:22]
      reg_7 <= 1'h0; // @[MatrixPRE-Processor.scala 21:22]
    end else begin
      reg_7 <= io_mat2_7_0 != 16'h0 | io_mat2_7_1 != 16'h0 | io_mat2_7_2 != 16'h0 | io_mat2_7_3 != 16'h0 | io_mat2_7_4
         != 16'h0 | io_mat2_7_5 != 16'h0 | io_mat2_7_6 != 16'h0 | io_mat2_7_7 != 16'h0; // @[MatrixPRE-Processor.scala 23:16]
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 28:20]
      i <= 3'h0; // @[MatrixPRE-Processor.scala 28:20]
    end else begin
      i <= _i_T_1;
    end
    if (reset) begin // @[MatrixPRE-Processor.scala 29:20]
      j <= 3'h0; // @[MatrixPRE-Processor.scala 29:20]
    end else if (i == 3'h7) begin // @[MatrixPRE-Processor.scala 42:28]
      j <= _j_T_1; // @[MatrixPRE-Processor.scala 43:11]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  matReg1_0_0 = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  matReg1_0_1 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  matReg1_0_2 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  matReg1_0_3 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  matReg1_0_4 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  matReg1_0_5 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  matReg1_0_6 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  matReg1_0_7 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  matReg1_1_0 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  matReg1_1_1 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  matReg1_1_2 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  matReg1_1_3 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  matReg1_1_4 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  matReg1_1_5 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  matReg1_1_6 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  matReg1_1_7 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  matReg1_2_0 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  matReg1_2_1 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  matReg1_2_2 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  matReg1_2_3 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  matReg1_2_4 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  matReg1_2_5 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  matReg1_2_6 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  matReg1_2_7 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  matReg1_3_0 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  matReg1_3_1 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  matReg1_3_2 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  matReg1_3_3 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  matReg1_3_4 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  matReg1_3_5 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  matReg1_3_6 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  matReg1_3_7 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  matReg1_4_0 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  matReg1_4_1 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  matReg1_4_2 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  matReg1_4_3 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  matReg1_4_4 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  matReg1_4_5 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  matReg1_4_6 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  matReg1_4_7 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  matReg1_5_0 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  matReg1_5_1 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  matReg1_5_2 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  matReg1_5_3 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  matReg1_5_4 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  matReg1_5_5 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  matReg1_5_6 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  matReg1_5_7 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  matReg1_6_0 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  matReg1_6_1 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  matReg1_6_2 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  matReg1_6_3 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  matReg1_6_4 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  matReg1_6_5 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  matReg1_6_6 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  matReg1_6_7 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  matReg1_7_0 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  matReg1_7_1 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  matReg1_7_2 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  matReg1_7_3 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  matReg1_7_4 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  matReg1_7_5 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  matReg1_7_6 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  matReg1_7_7 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  reg_0 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  reg_1 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  reg_2 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  reg_3 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  reg_4 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  reg_5 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  reg_6 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  reg_7 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  i = _RAND_72[2:0];
  _RAND_73 = {1{`RANDOM}};
  j = _RAND_73[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Muxes(
  input         clock,
  input         reset,
  input  [15:0] io_mat1_0_0,
  input  [15:0] io_mat1_0_1,
  input  [15:0] io_mat1_0_2,
  input  [15:0] io_mat1_0_3,
  input  [15:0] io_mat1_0_4,
  input  [15:0] io_mat1_0_5,
  input  [15:0] io_mat1_0_6,
  input  [15:0] io_mat1_0_7,
  input  [15:0] io_mat1_1_0,
  input  [15:0] io_mat1_1_1,
  input  [15:0] io_mat1_1_2,
  input  [15:0] io_mat1_1_3,
  input  [15:0] io_mat1_1_4,
  input  [15:0] io_mat1_1_5,
  input  [15:0] io_mat1_1_6,
  input  [15:0] io_mat1_1_7,
  input  [15:0] io_mat1_2_0,
  input  [15:0] io_mat1_2_1,
  input  [15:0] io_mat1_2_2,
  input  [15:0] io_mat1_2_3,
  input  [15:0] io_mat1_2_4,
  input  [15:0] io_mat1_2_5,
  input  [15:0] io_mat1_2_6,
  input  [15:0] io_mat1_2_7,
  input  [15:0] io_mat1_3_0,
  input  [15:0] io_mat1_3_1,
  input  [15:0] io_mat1_3_2,
  input  [15:0] io_mat1_3_3,
  input  [15:0] io_mat1_3_4,
  input  [15:0] io_mat1_3_5,
  input  [15:0] io_mat1_3_6,
  input  [15:0] io_mat1_3_7,
  input  [15:0] io_mat1_4_0,
  input  [15:0] io_mat1_4_1,
  input  [15:0] io_mat1_4_2,
  input  [15:0] io_mat1_4_3,
  input  [15:0] io_mat1_4_4,
  input  [15:0] io_mat1_4_5,
  input  [15:0] io_mat1_4_6,
  input  [15:0] io_mat1_4_7,
  input  [15:0] io_mat1_5_0,
  input  [15:0] io_mat1_5_1,
  input  [15:0] io_mat1_5_2,
  input  [15:0] io_mat1_5_3,
  input  [15:0] io_mat1_5_4,
  input  [15:0] io_mat1_5_5,
  input  [15:0] io_mat1_5_6,
  input  [15:0] io_mat1_5_7,
  input  [15:0] io_mat1_6_0,
  input  [15:0] io_mat1_6_1,
  input  [15:0] io_mat1_6_2,
  input  [15:0] io_mat1_6_3,
  input  [15:0] io_mat1_6_4,
  input  [15:0] io_mat1_6_5,
  input  [15:0] io_mat1_6_6,
  input  [15:0] io_mat1_6_7,
  input  [15:0] io_mat1_7_0,
  input  [15:0] io_mat1_7_1,
  input  [15:0] io_mat1_7_2,
  input  [15:0] io_mat1_7_3,
  input  [15:0] io_mat1_7_4,
  input  [15:0] io_mat1_7_5,
  input  [15:0] io_mat1_7_6,
  input  [15:0] io_mat1_7_7,
  input  [15:0] io_mat2_0,
  input  [15:0] io_mat2_1,
  input  [15:0] io_mat2_2,
  input  [15:0] io_mat2_3,
  input  [15:0] io_mat2_4,
  input  [15:0] io_mat2_5,
  input  [15:0] io_mat2_6,
  input  [15:0] io_mat2_7,
  input  [15:0] io_counterMatrix1_0_0,
  input  [15:0] io_counterMatrix1_0_1,
  input  [15:0] io_counterMatrix1_0_2,
  input  [15:0] io_counterMatrix1_0_3,
  input  [15:0] io_counterMatrix1_0_4,
  input  [15:0] io_counterMatrix1_0_5,
  input  [15:0] io_counterMatrix1_0_6,
  input  [15:0] io_counterMatrix1_0_7,
  input  [15:0] io_counterMatrix1_1_0,
  input  [15:0] io_counterMatrix1_1_1,
  input  [15:0] io_counterMatrix1_1_2,
  input  [15:0] io_counterMatrix1_1_3,
  input  [15:0] io_counterMatrix1_1_4,
  input  [15:0] io_counterMatrix1_1_5,
  input  [15:0] io_counterMatrix1_1_6,
  input  [15:0] io_counterMatrix1_1_7,
  input  [15:0] io_counterMatrix1_2_0,
  input  [15:0] io_counterMatrix1_2_1,
  input  [15:0] io_counterMatrix1_2_2,
  input  [15:0] io_counterMatrix1_2_3,
  input  [15:0] io_counterMatrix1_2_4,
  input  [15:0] io_counterMatrix1_2_5,
  input  [15:0] io_counterMatrix1_2_6,
  input  [15:0] io_counterMatrix1_2_7,
  input  [15:0] io_counterMatrix1_3_0,
  input  [15:0] io_counterMatrix1_3_1,
  input  [15:0] io_counterMatrix1_3_2,
  input  [15:0] io_counterMatrix1_3_3,
  input  [15:0] io_counterMatrix1_3_4,
  input  [15:0] io_counterMatrix1_3_5,
  input  [15:0] io_counterMatrix1_3_6,
  input  [15:0] io_counterMatrix1_3_7,
  input  [15:0] io_counterMatrix1_4_0,
  input  [15:0] io_counterMatrix1_4_1,
  input  [15:0] io_counterMatrix1_4_2,
  input  [15:0] io_counterMatrix1_4_3,
  input  [15:0] io_counterMatrix1_4_4,
  input  [15:0] io_counterMatrix1_4_5,
  input  [15:0] io_counterMatrix1_4_6,
  input  [15:0] io_counterMatrix1_4_7,
  input  [15:0] io_counterMatrix1_5_0,
  input  [15:0] io_counterMatrix1_5_1,
  input  [15:0] io_counterMatrix1_5_2,
  input  [15:0] io_counterMatrix1_5_3,
  input  [15:0] io_counterMatrix1_5_4,
  input  [15:0] io_counterMatrix1_5_5,
  input  [15:0] io_counterMatrix1_5_6,
  input  [15:0] io_counterMatrix1_5_7,
  input  [15:0] io_counterMatrix1_6_0,
  input  [15:0] io_counterMatrix1_6_1,
  input  [15:0] io_counterMatrix1_6_2,
  input  [15:0] io_counterMatrix1_6_3,
  input  [15:0] io_counterMatrix1_6_4,
  input  [15:0] io_counterMatrix1_6_5,
  input  [15:0] io_counterMatrix1_6_6,
  input  [15:0] io_counterMatrix1_6_7,
  input  [15:0] io_counterMatrix1_7_0,
  input  [15:0] io_counterMatrix1_7_1,
  input  [15:0] io_counterMatrix1_7_2,
  input  [15:0] io_counterMatrix1_7_3,
  input  [15:0] io_counterMatrix1_7_4,
  input  [15:0] io_counterMatrix1_7_5,
  input  [15:0] io_counterMatrix1_7_6,
  input  [15:0] io_counterMatrix1_7_7,
  input  [15:0] io_counterMatrix2_0,
  input  [15:0] io_counterMatrix2_1,
  input  [15:0] io_counterMatrix2_2,
  input  [15:0] io_counterMatrix2_3,
  input  [15:0] io_counterMatrix2_4,
  input  [15:0] io_counterMatrix2_5,
  input  [15:0] io_counterMatrix2_6,
  input  [15:0] io_counterMatrix2_7,
  output [3:0]  io_i_mux_bus_0,
  output [3:0]  io_i_mux_bus_1,
  output [3:0]  io_i_mux_bus_2,
  output [3:0]  io_i_mux_bus_3,
  output [15:0] io_Source_0,
  output [15:0] io_Source_1,
  output [15:0] io_Source_2,
  output [15:0] io_Source_3,
  output        io_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
`endif // RANDOMIZE_REG_INIT
  reg [15:0] prevStationary_matrix_0_0; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_0_1; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_0_2; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_0_3; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_0_4; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_0_5; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_0_6; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_0_7; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_1_0; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_1_1; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_1_2; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_1_3; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_1_4; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_1_5; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_1_6; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_1_7; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_2_0; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_2_1; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_2_2; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_2_3; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_2_4; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_2_5; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_2_6; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_2_7; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_3_0; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_3_1; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_3_2; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_3_3; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_3_4; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_3_5; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_3_6; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_3_7; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_4_0; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_4_1; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_4_2; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_4_3; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_4_4; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_4_5; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_4_6; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_4_7; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_5_0; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_5_1; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_5_2; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_5_3; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_5_4; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_5_5; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_5_6; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_5_7; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_6_0; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_6_1; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_6_2; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_6_3; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_6_4; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_6_5; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_6_6; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_6_7; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_7_0; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_7_1; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_7_2; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_7_3; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_7_4; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_7_5; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_7_6; // @[Muxes.scala 19:40]
  reg [15:0] prevStationary_matrix_7_7; // @[Muxes.scala 19:40]
  reg [15:0] prevStreaming_matrix_0; // @[Muxes.scala 20:39]
  reg [15:0] prevStreaming_matrix_1; // @[Muxes.scala 20:39]
  reg [15:0] prevStreaming_matrix_2; // @[Muxes.scala 20:39]
  reg [15:0] prevStreaming_matrix_3; // @[Muxes.scala 20:39]
  reg [15:0] prevStreaming_matrix_4; // @[Muxes.scala 20:39]
  reg [15:0] prevStreaming_matrix_5; // @[Muxes.scala 20:39]
  reg [15:0] prevStreaming_matrix_6; // @[Muxes.scala 20:39]
  reg [15:0] prevStreaming_matrix_7; // @[Muxes.scala 20:39]
  reg  matricesAreEqual; // @[Muxes.scala 21:31]
  reg  jValid; // @[Muxes.scala 27:25]
  reg [31:0] i; // @[Muxes.scala 28:20]
  reg [31:0] j; // @[Muxes.scala 29:20]
  reg [31:0] k; // @[Muxes.scala 30:20]
  reg [31:0] counter; // @[Muxes.scala 31:26]
  reg [3:0] mux_0; // @[Muxes.scala 32:22]
  reg [3:0] mux_1; // @[Muxes.scala 32:22]
  reg [3:0] mux_2; // @[Muxes.scala 32:22]
  reg [3:0] mux_3; // @[Muxes.scala 32:22]
  reg [15:0] src_0; // @[Muxes.scala 33:22]
  reg [15:0] src_1; // @[Muxes.scala 33:22]
  reg [15:0] src_2; // @[Muxes.scala 33:22]
  reg [15:0] src_3; // @[Muxes.scala 33:22]
  reg [15:0] dest_0; // @[Muxes.scala 34:23]
  reg [15:0] dest_1; // @[Muxes.scala 34:23]
  reg [15:0] dest_2; // @[Muxes.scala 34:23]
  reg [15:0] dest_3; // @[Muxes.scala 34:23]
  wire  _GEN_0 = io_mat1_0_0 != prevStationary_matrix_0_0 ? 1'h0 : 1'h1; // @[Muxes.scala 22:22 45:61 46:28]
  wire  _GEN_1 = io_mat1_0_1 != prevStationary_matrix_0_1 ? 1'h0 : _GEN_0; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_2 = io_mat1_0_2 != prevStationary_matrix_0_2 ? 1'h0 : _GEN_1; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_3 = io_mat1_0_3 != prevStationary_matrix_0_3 ? 1'h0 : _GEN_2; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_4 = io_mat1_0_4 != prevStationary_matrix_0_4 ? 1'h0 : _GEN_3; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_5 = io_mat1_0_5 != prevStationary_matrix_0_5 ? 1'h0 : _GEN_4; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_6 = io_mat1_0_6 != prevStationary_matrix_0_6 ? 1'h0 : _GEN_5; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_7 = io_mat1_0_7 != prevStationary_matrix_0_7 ? 1'h0 : _GEN_6; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_8 = io_mat2_0 != prevStreaming_matrix_0 ? 1'h0 : _GEN_7; // @[Muxes.scala 49:51 50:26]
  wire  _GEN_9 = io_mat1_1_0 != prevStationary_matrix_1_0 ? 1'h0 : _GEN_8; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_10 = io_mat1_1_1 != prevStationary_matrix_1_1 ? 1'h0 : _GEN_9; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_11 = io_mat1_1_2 != prevStationary_matrix_1_2 ? 1'h0 : _GEN_10; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_12 = io_mat1_1_3 != prevStationary_matrix_1_3 ? 1'h0 : _GEN_11; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_13 = io_mat1_1_4 != prevStationary_matrix_1_4 ? 1'h0 : _GEN_12; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_14 = io_mat1_1_5 != prevStationary_matrix_1_5 ? 1'h0 : _GEN_13; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_15 = io_mat1_1_6 != prevStationary_matrix_1_6 ? 1'h0 : _GEN_14; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_16 = io_mat1_1_7 != prevStationary_matrix_1_7 ? 1'h0 : _GEN_15; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_17 = io_mat2_1 != prevStreaming_matrix_1 ? 1'h0 : _GEN_16; // @[Muxes.scala 49:51 50:26]
  wire  _GEN_18 = io_mat1_2_0 != prevStationary_matrix_2_0 ? 1'h0 : _GEN_17; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_19 = io_mat1_2_1 != prevStationary_matrix_2_1 ? 1'h0 : _GEN_18; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_20 = io_mat1_2_2 != prevStationary_matrix_2_2 ? 1'h0 : _GEN_19; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_21 = io_mat1_2_3 != prevStationary_matrix_2_3 ? 1'h0 : _GEN_20; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_22 = io_mat1_2_4 != prevStationary_matrix_2_4 ? 1'h0 : _GEN_21; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_23 = io_mat1_2_5 != prevStationary_matrix_2_5 ? 1'h0 : _GEN_22; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_24 = io_mat1_2_6 != prevStationary_matrix_2_6 ? 1'h0 : _GEN_23; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_25 = io_mat1_2_7 != prevStationary_matrix_2_7 ? 1'h0 : _GEN_24; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_26 = io_mat2_2 != prevStreaming_matrix_2 ? 1'h0 : _GEN_25; // @[Muxes.scala 49:51 50:26]
  wire  _GEN_27 = io_mat1_3_0 != prevStationary_matrix_3_0 ? 1'h0 : _GEN_26; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_28 = io_mat1_3_1 != prevStationary_matrix_3_1 ? 1'h0 : _GEN_27; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_29 = io_mat1_3_2 != prevStationary_matrix_3_2 ? 1'h0 : _GEN_28; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_30 = io_mat1_3_3 != prevStationary_matrix_3_3 ? 1'h0 : _GEN_29; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_31 = io_mat1_3_4 != prevStationary_matrix_3_4 ? 1'h0 : _GEN_30; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_32 = io_mat1_3_5 != prevStationary_matrix_3_5 ? 1'h0 : _GEN_31; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_33 = io_mat1_3_6 != prevStationary_matrix_3_6 ? 1'h0 : _GEN_32; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_34 = io_mat1_3_7 != prevStationary_matrix_3_7 ? 1'h0 : _GEN_33; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_35 = io_mat2_3 != prevStreaming_matrix_3 ? 1'h0 : _GEN_34; // @[Muxes.scala 49:51 50:26]
  wire  _GEN_36 = io_mat1_4_0 != prevStationary_matrix_4_0 ? 1'h0 : _GEN_35; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_37 = io_mat1_4_1 != prevStationary_matrix_4_1 ? 1'h0 : _GEN_36; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_38 = io_mat1_4_2 != prevStationary_matrix_4_2 ? 1'h0 : _GEN_37; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_39 = io_mat1_4_3 != prevStationary_matrix_4_3 ? 1'h0 : _GEN_38; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_40 = io_mat1_4_4 != prevStationary_matrix_4_4 ? 1'h0 : _GEN_39; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_41 = io_mat1_4_5 != prevStationary_matrix_4_5 ? 1'h0 : _GEN_40; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_42 = io_mat1_4_6 != prevStationary_matrix_4_6 ? 1'h0 : _GEN_41; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_43 = io_mat1_4_7 != prevStationary_matrix_4_7 ? 1'h0 : _GEN_42; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_44 = io_mat2_4 != prevStreaming_matrix_4 ? 1'h0 : _GEN_43; // @[Muxes.scala 49:51 50:26]
  wire  _GEN_45 = io_mat1_5_0 != prevStationary_matrix_5_0 ? 1'h0 : _GEN_44; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_46 = io_mat1_5_1 != prevStationary_matrix_5_1 ? 1'h0 : _GEN_45; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_47 = io_mat1_5_2 != prevStationary_matrix_5_2 ? 1'h0 : _GEN_46; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_48 = io_mat1_5_3 != prevStationary_matrix_5_3 ? 1'h0 : _GEN_47; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_49 = io_mat1_5_4 != prevStationary_matrix_5_4 ? 1'h0 : _GEN_48; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_50 = io_mat1_5_5 != prevStationary_matrix_5_5 ? 1'h0 : _GEN_49; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_51 = io_mat1_5_6 != prevStationary_matrix_5_6 ? 1'h0 : _GEN_50; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_52 = io_mat1_5_7 != prevStationary_matrix_5_7 ? 1'h0 : _GEN_51; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_53 = io_mat2_5 != prevStreaming_matrix_5 ? 1'h0 : _GEN_52; // @[Muxes.scala 49:51 50:26]
  wire  _GEN_54 = io_mat1_6_0 != prevStationary_matrix_6_0 ? 1'h0 : _GEN_53; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_55 = io_mat1_6_1 != prevStationary_matrix_6_1 ? 1'h0 : _GEN_54; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_56 = io_mat1_6_2 != prevStationary_matrix_6_2 ? 1'h0 : _GEN_55; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_57 = io_mat1_6_3 != prevStationary_matrix_6_3 ? 1'h0 : _GEN_56; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_58 = io_mat1_6_4 != prevStationary_matrix_6_4 ? 1'h0 : _GEN_57; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_59 = io_mat1_6_5 != prevStationary_matrix_6_5 ? 1'h0 : _GEN_58; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_60 = io_mat1_6_6 != prevStationary_matrix_6_6 ? 1'h0 : _GEN_59; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_61 = io_mat1_6_7 != prevStationary_matrix_6_7 ? 1'h0 : _GEN_60; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_62 = io_mat2_6 != prevStreaming_matrix_6 ? 1'h0 : _GEN_61; // @[Muxes.scala 49:51 50:26]
  wire  _GEN_63 = io_mat1_7_0 != prevStationary_matrix_7_0 ? 1'h0 : _GEN_62; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_64 = io_mat1_7_1 != prevStationary_matrix_7_1 ? 1'h0 : _GEN_63; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_65 = io_mat1_7_2 != prevStationary_matrix_7_2 ? 1'h0 : _GEN_64; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_66 = io_mat1_7_3 != prevStationary_matrix_7_3 ? 1'h0 : _GEN_65; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_67 = io_mat1_7_4 != prevStationary_matrix_7_4 ? 1'h0 : _GEN_66; // @[Muxes.scala 45:61 46:28]
  wire  _GEN_596 = 3'h0 == j[2:0]; // @[Muxes.scala 54:{36,36}]
  wire  _GEN_597 = 3'h1 == i[2:0]; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_73 = 3'h0 == j[2:0] & 3'h1 == i[2:0] ? io_counterMatrix1_0_1 : io_counterMatrix1_0_0; // @[Muxes.scala 54:{36,36}]
  wire  _GEN_599 = 3'h2 == i[2:0]; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_74 = 3'h0 == j[2:0] & 3'h2 == i[2:0] ? io_counterMatrix1_0_2 : _GEN_73; // @[Muxes.scala 54:{36,36}]
  wire  _GEN_601 = 3'h3 == i[2:0]; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_75 = 3'h0 == j[2:0] & 3'h3 == i[2:0] ? io_counterMatrix1_0_3 : _GEN_74; // @[Muxes.scala 54:{36,36}]
  wire  _GEN_603 = 3'h4 == i[2:0]; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_76 = 3'h0 == j[2:0] & 3'h4 == i[2:0] ? io_counterMatrix1_0_4 : _GEN_75; // @[Muxes.scala 54:{36,36}]
  wire  _GEN_605 = 3'h5 == i[2:0]; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_77 = 3'h0 == j[2:0] & 3'h5 == i[2:0] ? io_counterMatrix1_0_5 : _GEN_76; // @[Muxes.scala 54:{36,36}]
  wire  _GEN_607 = 3'h6 == i[2:0]; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_78 = 3'h0 == j[2:0] & 3'h6 == i[2:0] ? io_counterMatrix1_0_6 : _GEN_77; // @[Muxes.scala 54:{36,36}]
  wire  _GEN_609 = 3'h7 == i[2:0]; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_79 = 3'h0 == j[2:0] & 3'h7 == i[2:0] ? io_counterMatrix1_0_7 : _GEN_78; // @[Muxes.scala 54:{36,36}]
  wire  _GEN_610 = 3'h1 == j[2:0]; // @[Muxes.scala 54:{36,36}]
  wire  _GEN_611 = 3'h0 == i[2:0]; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_80 = 3'h1 == j[2:0] & 3'h0 == i[2:0] ? io_counterMatrix1_1_0 : _GEN_79; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_81 = 3'h1 == j[2:0] & 3'h1 == i[2:0] ? io_counterMatrix1_1_1 : _GEN_80; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_82 = 3'h1 == j[2:0] & 3'h2 == i[2:0] ? io_counterMatrix1_1_2 : _GEN_81; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_83 = 3'h1 == j[2:0] & 3'h3 == i[2:0] ? io_counterMatrix1_1_3 : _GEN_82; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_84 = 3'h1 == j[2:0] & 3'h4 == i[2:0] ? io_counterMatrix1_1_4 : _GEN_83; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_85 = 3'h1 == j[2:0] & 3'h5 == i[2:0] ? io_counterMatrix1_1_5 : _GEN_84; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_86 = 3'h1 == j[2:0] & 3'h6 == i[2:0] ? io_counterMatrix1_1_6 : _GEN_85; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_87 = 3'h1 == j[2:0] & 3'h7 == i[2:0] ? io_counterMatrix1_1_7 : _GEN_86; // @[Muxes.scala 54:{36,36}]
  wire  _GEN_626 = 3'h2 == j[2:0]; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_88 = 3'h2 == j[2:0] & 3'h0 == i[2:0] ? io_counterMatrix1_2_0 : _GEN_87; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_89 = 3'h2 == j[2:0] & 3'h1 == i[2:0] ? io_counterMatrix1_2_1 : _GEN_88; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_90 = 3'h2 == j[2:0] & 3'h2 == i[2:0] ? io_counterMatrix1_2_2 : _GEN_89; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_91 = 3'h2 == j[2:0] & 3'h3 == i[2:0] ? io_counterMatrix1_2_3 : _GEN_90; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_92 = 3'h2 == j[2:0] & 3'h4 == i[2:0] ? io_counterMatrix1_2_4 : _GEN_91; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_93 = 3'h2 == j[2:0] & 3'h5 == i[2:0] ? io_counterMatrix1_2_5 : _GEN_92; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_94 = 3'h2 == j[2:0] & 3'h6 == i[2:0] ? io_counterMatrix1_2_6 : _GEN_93; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_95 = 3'h2 == j[2:0] & 3'h7 == i[2:0] ? io_counterMatrix1_2_7 : _GEN_94; // @[Muxes.scala 54:{36,36}]
  wire  _GEN_642 = 3'h3 == j[2:0]; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_96 = 3'h3 == j[2:0] & 3'h0 == i[2:0] ? io_counterMatrix1_3_0 : _GEN_95; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_97 = 3'h3 == j[2:0] & 3'h1 == i[2:0] ? io_counterMatrix1_3_1 : _GEN_96; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_98 = 3'h3 == j[2:0] & 3'h2 == i[2:0] ? io_counterMatrix1_3_2 : _GEN_97; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_99 = 3'h3 == j[2:0] & 3'h3 == i[2:0] ? io_counterMatrix1_3_3 : _GEN_98; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_100 = 3'h3 == j[2:0] & 3'h4 == i[2:0] ? io_counterMatrix1_3_4 : _GEN_99; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_101 = 3'h3 == j[2:0] & 3'h5 == i[2:0] ? io_counterMatrix1_3_5 : _GEN_100; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_102 = 3'h3 == j[2:0] & 3'h6 == i[2:0] ? io_counterMatrix1_3_6 : _GEN_101; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_103 = 3'h3 == j[2:0] & 3'h7 == i[2:0] ? io_counterMatrix1_3_7 : _GEN_102; // @[Muxes.scala 54:{36,36}]
  wire  _GEN_658 = 3'h4 == j[2:0]; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_104 = 3'h4 == j[2:0] & 3'h0 == i[2:0] ? io_counterMatrix1_4_0 : _GEN_103; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_105 = 3'h4 == j[2:0] & 3'h1 == i[2:0] ? io_counterMatrix1_4_1 : _GEN_104; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_106 = 3'h4 == j[2:0] & 3'h2 == i[2:0] ? io_counterMatrix1_4_2 : _GEN_105; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_107 = 3'h4 == j[2:0] & 3'h3 == i[2:0] ? io_counterMatrix1_4_3 : _GEN_106; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_108 = 3'h4 == j[2:0] & 3'h4 == i[2:0] ? io_counterMatrix1_4_4 : _GEN_107; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_109 = 3'h4 == j[2:0] & 3'h5 == i[2:0] ? io_counterMatrix1_4_5 : _GEN_108; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_110 = 3'h4 == j[2:0] & 3'h6 == i[2:0] ? io_counterMatrix1_4_6 : _GEN_109; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_111 = 3'h4 == j[2:0] & 3'h7 == i[2:0] ? io_counterMatrix1_4_7 : _GEN_110; // @[Muxes.scala 54:{36,36}]
  wire  _GEN_674 = 3'h5 == j[2:0]; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_112 = 3'h5 == j[2:0] & 3'h0 == i[2:0] ? io_counterMatrix1_5_0 : _GEN_111; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_113 = 3'h5 == j[2:0] & 3'h1 == i[2:0] ? io_counterMatrix1_5_1 : _GEN_112; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_114 = 3'h5 == j[2:0] & 3'h2 == i[2:0] ? io_counterMatrix1_5_2 : _GEN_113; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_115 = 3'h5 == j[2:0] & 3'h3 == i[2:0] ? io_counterMatrix1_5_3 : _GEN_114; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_116 = 3'h5 == j[2:0] & 3'h4 == i[2:0] ? io_counterMatrix1_5_4 : _GEN_115; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_117 = 3'h5 == j[2:0] & 3'h5 == i[2:0] ? io_counterMatrix1_5_5 : _GEN_116; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_118 = 3'h5 == j[2:0] & 3'h6 == i[2:0] ? io_counterMatrix1_5_6 : _GEN_117; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_119 = 3'h5 == j[2:0] & 3'h7 == i[2:0] ? io_counterMatrix1_5_7 : _GEN_118; // @[Muxes.scala 54:{36,36}]
  wire  _GEN_690 = 3'h6 == j[2:0]; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_120 = 3'h6 == j[2:0] & 3'h0 == i[2:0] ? io_counterMatrix1_6_0 : _GEN_119; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_121 = 3'h6 == j[2:0] & 3'h1 == i[2:0] ? io_counterMatrix1_6_1 : _GEN_120; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_122 = 3'h6 == j[2:0] & 3'h2 == i[2:0] ? io_counterMatrix1_6_2 : _GEN_121; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_123 = 3'h6 == j[2:0] & 3'h3 == i[2:0] ? io_counterMatrix1_6_3 : _GEN_122; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_124 = 3'h6 == j[2:0] & 3'h4 == i[2:0] ? io_counterMatrix1_6_4 : _GEN_123; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_125 = 3'h6 == j[2:0] & 3'h5 == i[2:0] ? io_counterMatrix1_6_5 : _GEN_124; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_126 = 3'h6 == j[2:0] & 3'h6 == i[2:0] ? io_counterMatrix1_6_6 : _GEN_125; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_127 = 3'h6 == j[2:0] & 3'h7 == i[2:0] ? io_counterMatrix1_6_7 : _GEN_126; // @[Muxes.scala 54:{36,36}]
  wire  _GEN_706 = 3'h7 == j[2:0]; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_128 = 3'h7 == j[2:0] & 3'h0 == i[2:0] ? io_counterMatrix1_7_0 : _GEN_127; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_129 = 3'h7 == j[2:0] & 3'h1 == i[2:0] ? io_counterMatrix1_7_1 : _GEN_128; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_130 = 3'h7 == j[2:0] & 3'h2 == i[2:0] ? io_counterMatrix1_7_2 : _GEN_129; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_131 = 3'h7 == j[2:0] & 3'h3 == i[2:0] ? io_counterMatrix1_7_3 : _GEN_130; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_132 = 3'h7 == j[2:0] & 3'h4 == i[2:0] ? io_counterMatrix1_7_4 : _GEN_131; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_133 = 3'h7 == j[2:0] & 3'h5 == i[2:0] ? io_counterMatrix1_7_5 : _GEN_132; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_134 = 3'h7 == j[2:0] & 3'h6 == i[2:0] ? io_counterMatrix1_7_6 : _GEN_133; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_135 = 3'h7 == j[2:0] & 3'h7 == i[2:0] ? io_counterMatrix1_7_7 : _GEN_134; // @[Muxes.scala 54:{36,36}]
  wire [15:0] _GEN_137 = 3'h1 == i[2:0] ? io_mat2_1 : io_mat2_0; // @[Muxes.scala 54:{60,60}]
  wire [15:0] _GEN_138 = 3'h2 == i[2:0] ? io_mat2_2 : _GEN_137; // @[Muxes.scala 54:{60,60}]
  wire [15:0] _GEN_139 = 3'h3 == i[2:0] ? io_mat2_3 : _GEN_138; // @[Muxes.scala 54:{60,60}]
  wire [15:0] _GEN_140 = 3'h4 == i[2:0] ? io_mat2_4 : _GEN_139; // @[Muxes.scala 54:{60,60}]
  wire [15:0] _GEN_141 = 3'h5 == i[2:0] ? io_mat2_5 : _GEN_140; // @[Muxes.scala 54:{60,60}]
  wire [15:0] _GEN_142 = 3'h6 == i[2:0] ? io_mat2_6 : _GEN_141; // @[Muxes.scala 54:{60,60}]
  wire [15:0] _GEN_143 = 3'h7 == i[2:0] ? io_mat2_7 : _GEN_142; // @[Muxes.scala 54:{60,60}]
  wire [15:0] _GEN_209 = 3'h1 == i[2:0] ? io_counterMatrix2_1 : io_counterMatrix2_0; // @[Muxes.scala 56:{38,38}]
  wire [15:0] _GEN_210 = 3'h2 == i[2:0] ? io_counterMatrix2_2 : _GEN_209; // @[Muxes.scala 56:{38,38}]
  wire [15:0] _GEN_211 = 3'h3 == i[2:0] ? io_counterMatrix2_3 : _GEN_210; // @[Muxes.scala 56:{38,38}]
  wire [15:0] _GEN_212 = 3'h4 == i[2:0] ? io_counterMatrix2_4 : _GEN_211; // @[Muxes.scala 56:{38,38}]
  wire [15:0] _GEN_213 = 3'h5 == i[2:0] ? io_counterMatrix2_5 : _GEN_212; // @[Muxes.scala 56:{38,38}]
  wire [15:0] _GEN_214 = 3'h6 == i[2:0] ? io_counterMatrix2_6 : _GEN_213; // @[Muxes.scala 56:{38,38}]
  wire [15:0] _GEN_215 = 3'h7 == i[2:0] ? io_counterMatrix2_7 : _GEN_214; // @[Muxes.scala 56:{38,38}]
  wire [15:0] _mux_T_2 = _GEN_215 - 16'h1; // @[Muxes.scala 57:51]
  wire [15:0] _mux_T_6 = _GEN_135 - 16'h1; // @[Muxes.scala 57:85]
  wire [15:0] _mux_T_8 = _mux_T_2 - _mux_T_6; // @[Muxes.scala 57:58]
  wire [3:0] _GEN_288 = 2'h0 == counter[1:0] ? _mux_T_8[3:0] : mux_0; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_289 = 2'h1 == counter[1:0] ? _mux_T_8[3:0] : mux_1; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_290 = 2'h2 == counter[1:0] ? _mux_T_8[3:0] : mux_2; // @[Muxes.scala 32:22 57:{24,24}]
  wire [3:0] _GEN_291 = 2'h3 == counter[1:0] ? _mux_T_8[3:0] : mux_3; // @[Muxes.scala 32:22 57:{24,24}]
  wire [15:0] _GEN_292 = 2'h0 == counter[1:0] ? _GEN_143 : src_0; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_293 = 2'h1 == counter[1:0] ? _GEN_143 : src_1; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_294 = 2'h2 == counter[1:0] ? _GEN_143 : src_2; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_295 = 2'h3 == counter[1:0] ? _GEN_143 : src_3; // @[Muxes.scala 33:22 58:{24,24}]
  wire [15:0] _GEN_309 = _GEN_596 & _GEN_597 ? io_mat1_0_1 : io_mat1_0_0; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_310 = _GEN_596 & _GEN_599 ? io_mat1_0_2 : _GEN_309; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_311 = _GEN_596 & _GEN_601 ? io_mat1_0_3 : _GEN_310; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_312 = _GEN_596 & _GEN_603 ? io_mat1_0_4 : _GEN_311; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_313 = _GEN_596 & _GEN_605 ? io_mat1_0_5 : _GEN_312; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_314 = _GEN_596 & _GEN_607 ? io_mat1_0_6 : _GEN_313; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_315 = _GEN_596 & _GEN_609 ? io_mat1_0_7 : _GEN_314; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_316 = _GEN_610 & _GEN_611 ? io_mat1_1_0 : _GEN_315; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_317 = _GEN_610 & _GEN_597 ? io_mat1_1_1 : _GEN_316; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_318 = _GEN_610 & _GEN_599 ? io_mat1_1_2 : _GEN_317; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_319 = _GEN_610 & _GEN_601 ? io_mat1_1_3 : _GEN_318; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_320 = _GEN_610 & _GEN_603 ? io_mat1_1_4 : _GEN_319; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_321 = _GEN_610 & _GEN_605 ? io_mat1_1_5 : _GEN_320; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_322 = _GEN_610 & _GEN_607 ? io_mat1_1_6 : _GEN_321; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_323 = _GEN_610 & _GEN_609 ? io_mat1_1_7 : _GEN_322; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_324 = _GEN_626 & _GEN_611 ? io_mat1_2_0 : _GEN_323; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_325 = _GEN_626 & _GEN_597 ? io_mat1_2_1 : _GEN_324; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_326 = _GEN_626 & _GEN_599 ? io_mat1_2_2 : _GEN_325; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_327 = _GEN_626 & _GEN_601 ? io_mat1_2_3 : _GEN_326; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_328 = _GEN_626 & _GEN_603 ? io_mat1_2_4 : _GEN_327; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_329 = _GEN_626 & _GEN_605 ? io_mat1_2_5 : _GEN_328; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_330 = _GEN_626 & _GEN_607 ? io_mat1_2_6 : _GEN_329; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_331 = _GEN_626 & _GEN_609 ? io_mat1_2_7 : _GEN_330; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_332 = _GEN_642 & _GEN_611 ? io_mat1_3_0 : _GEN_331; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_333 = _GEN_642 & _GEN_597 ? io_mat1_3_1 : _GEN_332; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_334 = _GEN_642 & _GEN_599 ? io_mat1_3_2 : _GEN_333; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_335 = _GEN_642 & _GEN_601 ? io_mat1_3_3 : _GEN_334; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_336 = _GEN_642 & _GEN_603 ? io_mat1_3_4 : _GEN_335; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_337 = _GEN_642 & _GEN_605 ? io_mat1_3_5 : _GEN_336; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_338 = _GEN_642 & _GEN_607 ? io_mat1_3_6 : _GEN_337; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_339 = _GEN_642 & _GEN_609 ? io_mat1_3_7 : _GEN_338; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_340 = _GEN_658 & _GEN_611 ? io_mat1_4_0 : _GEN_339; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_341 = _GEN_658 & _GEN_597 ? io_mat1_4_1 : _GEN_340; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_342 = _GEN_658 & _GEN_599 ? io_mat1_4_2 : _GEN_341; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_343 = _GEN_658 & _GEN_601 ? io_mat1_4_3 : _GEN_342; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_344 = _GEN_658 & _GEN_603 ? io_mat1_4_4 : _GEN_343; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_345 = _GEN_658 & _GEN_605 ? io_mat1_4_5 : _GEN_344; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_346 = _GEN_658 & _GEN_607 ? io_mat1_4_6 : _GEN_345; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_347 = _GEN_658 & _GEN_609 ? io_mat1_4_7 : _GEN_346; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_348 = _GEN_674 & _GEN_611 ? io_mat1_5_0 : _GEN_347; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_349 = _GEN_674 & _GEN_597 ? io_mat1_5_1 : _GEN_348; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_350 = _GEN_674 & _GEN_599 ? io_mat1_5_2 : _GEN_349; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_351 = _GEN_674 & _GEN_601 ? io_mat1_5_3 : _GEN_350; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_352 = _GEN_674 & _GEN_603 ? io_mat1_5_4 : _GEN_351; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_353 = _GEN_674 & _GEN_605 ? io_mat1_5_5 : _GEN_352; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_354 = _GEN_674 & _GEN_607 ? io_mat1_5_6 : _GEN_353; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_355 = _GEN_674 & _GEN_609 ? io_mat1_5_7 : _GEN_354; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_356 = _GEN_690 & _GEN_611 ? io_mat1_6_0 : _GEN_355; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_357 = _GEN_690 & _GEN_597 ? io_mat1_6_1 : _GEN_356; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_358 = _GEN_690 & _GEN_599 ? io_mat1_6_2 : _GEN_357; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_359 = _GEN_690 & _GEN_601 ? io_mat1_6_3 : _GEN_358; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_360 = _GEN_690 & _GEN_603 ? io_mat1_6_4 : _GEN_359; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_361 = _GEN_690 & _GEN_605 ? io_mat1_6_5 : _GEN_360; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_362 = _GEN_690 & _GEN_607 ? io_mat1_6_6 : _GEN_361; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_363 = _GEN_690 & _GEN_609 ? io_mat1_6_7 : _GEN_362; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_364 = _GEN_706 & _GEN_611 ? io_mat1_7_0 : _GEN_363; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_365 = _GEN_706 & _GEN_597 ? io_mat1_7_1 : _GEN_364; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_366 = _GEN_706 & _GEN_599 ? io_mat1_7_2 : _GEN_365; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_367 = _GEN_706 & _GEN_601 ? io_mat1_7_3 : _GEN_366; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_368 = _GEN_706 & _GEN_603 ? io_mat1_7_4 : _GEN_367; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_369 = _GEN_706 & _GEN_605 ? io_mat1_7_5 : _GEN_368; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_370 = _GEN_706 & _GEN_607 ? io_mat1_7_6 : _GEN_369; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_371 = _GEN_706 & _GEN_609 ? io_mat1_7_7 : _GEN_370; // @[Muxes.scala 59:{25,25}]
  wire [15:0] _GEN_304 = 2'h0 == counter[1:0] ? _GEN_371 : dest_0; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_305 = 2'h1 == counter[1:0] ? _GEN_371 : dest_1; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_306 = 2'h2 == counter[1:0] ? _GEN_371 : dest_2; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _GEN_307 = 2'h3 == counter[1:0] ? _GEN_371 : dest_3; // @[Muxes.scala 34:23 59:{25,25}]
  wire [15:0] _mux_T_17 = _mux_T_6 - _mux_T_2; // @[Muxes.scala 61:61]
  wire [3:0] _GEN_444 = 2'h0 == counter[1:0] ? _mux_T_17[3:0] : mux_0; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_445 = 2'h1 == counter[1:0] ? _mux_T_17[3:0] : mux_1; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_446 = 2'h2 == counter[1:0] ? _mux_T_17[3:0] : mux_2; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_447 = 2'h3 == counter[1:0] ? _mux_T_17[3:0] : mux_3; // @[Muxes.scala 32:22 61:{24,24}]
  wire [3:0] _GEN_528 = _GEN_135 <= _GEN_215 ? _GEN_288 : _GEN_444; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_529 = _GEN_135 <= _GEN_215 ? _GEN_289 : _GEN_445; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_530 = _GEN_135 <= _GEN_215 ? _GEN_290 : _GEN_446; // @[Muxes.scala 56:62]
  wire [3:0] _GEN_531 = _GEN_135 <= _GEN_215 ? _GEN_291 : _GEN_447; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_532 = _GEN_135 <= _GEN_215 ? _GEN_292 : _GEN_292; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_533 = _GEN_135 <= _GEN_215 ? _GEN_293 : _GEN_293; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_534 = _GEN_135 <= _GEN_215 ? _GEN_294 : _GEN_294; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_535 = _GEN_135 <= _GEN_215 ? _GEN_295 : _GEN_295; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_536 = _GEN_135 <= _GEN_215 ? _GEN_304 : _GEN_304; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_537 = _GEN_135 <= _GEN_215 ? _GEN_305 : _GEN_305; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_538 = _GEN_135 <= _GEN_215 ? _GEN_306 : _GEN_306; // @[Muxes.scala 56:62]
  wire [15:0] _GEN_539 = _GEN_135 <= _GEN_215 ? _GEN_307 : _GEN_307; // @[Muxes.scala 56:62]
  wire  _T_88 = ~jValid; // @[Muxes.scala 66:15]
  wire  _T_89 = j == 32'h7; // @[Muxes.scala 68:22]
  wire  _T_90 = i == 32'h7; // @[Muxes.scala 68:56]
  wire  _T_91 = j == 32'h7 & i == 32'h7; // @[Muxes.scala 68:50]
  wire [31:0] _counter_T_1 = counter + 32'h1; // @[Muxes.scala 69:30]
  wire [31:0] _GEN_540 = ~(j == 32'h7 & i == 32'h7) ? _counter_T_1 : counter; // @[Muxes.scala 68:85 69:19 31:26]
  wire [31:0] _GEN_541 = ~jValid ? _GEN_540 : counter; // @[Muxes.scala 66:24 31:26]
  wire [3:0] _GEN_542 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_528 : mux_0; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_543 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_529 : mux_1; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_544 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_530 : mux_2; // @[Muxes.scala 32:22 54:70]
  wire [3:0] _GEN_545 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_531 : mux_3; // @[Muxes.scala 32:22 54:70]
  wire [15:0] _GEN_546 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_532 : src_0; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_547 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_533 : src_1; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_548 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_534 : src_2; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_549 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_535 : src_3; // @[Muxes.scala 33:22 54:70]
  wire [15:0] _GEN_550 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_536 : dest_0; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_551 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_537 : dest_1; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_552 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_538 : dest_2; // @[Muxes.scala 34:23 54:70]
  wire [15:0] _GEN_553 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_539 : dest_3; // @[Muxes.scala 34:23 54:70]
  wire [31:0] _GEN_554 = _GEN_135 != 16'h0 & _GEN_143 != 16'h0 ? _GEN_541 : counter; // @[Muxes.scala 31:26 54:70]
  wire [31:0] _j_T_1 = j + 32'h1; // @[Muxes.scala 79:16]
  wire [31:0] _i_T_1 = i + 32'h1; // @[Muxes.scala 85:18]
  wire [31:0] _GEN_555 = i < 32'h7 ? _i_T_1 : i; // @[Muxes.scala 84:42 85:13 28:20]
  wire  _GEN_556 = _T_91 | jValid; // @[Muxes.scala 80:83 81:16 27:25]
  reg [31:0] jNext; // @[Muxes.scala 105:24]
  wire [31:0] _k_T_1 = k + 32'h1; // @[Muxes.scala 114:14]
  assign io_i_mux_bus_0 = mux_0; // @[Muxes.scala 35:18]
  assign io_i_mux_bus_1 = mux_1; // @[Muxes.scala 35:18]
  assign io_i_mux_bus_2 = mux_2; // @[Muxes.scala 35:18]
  assign io_i_mux_bus_3 = mux_3; // @[Muxes.scala 35:18]
  assign io_Source_0 = src_0; // @[Muxes.scala 36:15]
  assign io_Source_1 = src_1; // @[Muxes.scala 36:15]
  assign io_Source_2 = src_2; // @[Muxes.scala 36:15]
  assign io_Source_3 = src_3; // @[Muxes.scala 36:15]
  assign io_valid = k != 32'h0 & _T_89 & _T_90 & jNext == 32'h6; // @[Muxes.scala 108:86]
  always @(posedge clock) begin
    prevStationary_matrix_0_0 <= io_mat1_0_0; // @[Muxes.scala 19:40]
    prevStationary_matrix_0_1 <= io_mat1_0_1; // @[Muxes.scala 19:40]
    prevStationary_matrix_0_2 <= io_mat1_0_2; // @[Muxes.scala 19:40]
    prevStationary_matrix_0_3 <= io_mat1_0_3; // @[Muxes.scala 19:40]
    prevStationary_matrix_0_4 <= io_mat1_0_4; // @[Muxes.scala 19:40]
    prevStationary_matrix_0_5 <= io_mat1_0_5; // @[Muxes.scala 19:40]
    prevStationary_matrix_0_6 <= io_mat1_0_6; // @[Muxes.scala 19:40]
    prevStationary_matrix_0_7 <= io_mat1_0_7; // @[Muxes.scala 19:40]
    prevStationary_matrix_1_0 <= io_mat1_1_0; // @[Muxes.scala 19:40]
    prevStationary_matrix_1_1 <= io_mat1_1_1; // @[Muxes.scala 19:40]
    prevStationary_matrix_1_2 <= io_mat1_1_2; // @[Muxes.scala 19:40]
    prevStationary_matrix_1_3 <= io_mat1_1_3; // @[Muxes.scala 19:40]
    prevStationary_matrix_1_4 <= io_mat1_1_4; // @[Muxes.scala 19:40]
    prevStationary_matrix_1_5 <= io_mat1_1_5; // @[Muxes.scala 19:40]
    prevStationary_matrix_1_6 <= io_mat1_1_6; // @[Muxes.scala 19:40]
    prevStationary_matrix_1_7 <= io_mat1_1_7; // @[Muxes.scala 19:40]
    prevStationary_matrix_2_0 <= io_mat1_2_0; // @[Muxes.scala 19:40]
    prevStationary_matrix_2_1 <= io_mat1_2_1; // @[Muxes.scala 19:40]
    prevStationary_matrix_2_2 <= io_mat1_2_2; // @[Muxes.scala 19:40]
    prevStationary_matrix_2_3 <= io_mat1_2_3; // @[Muxes.scala 19:40]
    prevStationary_matrix_2_4 <= io_mat1_2_4; // @[Muxes.scala 19:40]
    prevStationary_matrix_2_5 <= io_mat1_2_5; // @[Muxes.scala 19:40]
    prevStationary_matrix_2_6 <= io_mat1_2_6; // @[Muxes.scala 19:40]
    prevStationary_matrix_2_7 <= io_mat1_2_7; // @[Muxes.scala 19:40]
    prevStationary_matrix_3_0 <= io_mat1_3_0; // @[Muxes.scala 19:40]
    prevStationary_matrix_3_1 <= io_mat1_3_1; // @[Muxes.scala 19:40]
    prevStationary_matrix_3_2 <= io_mat1_3_2; // @[Muxes.scala 19:40]
    prevStationary_matrix_3_3 <= io_mat1_3_3; // @[Muxes.scala 19:40]
    prevStationary_matrix_3_4 <= io_mat1_3_4; // @[Muxes.scala 19:40]
    prevStationary_matrix_3_5 <= io_mat1_3_5; // @[Muxes.scala 19:40]
    prevStationary_matrix_3_6 <= io_mat1_3_6; // @[Muxes.scala 19:40]
    prevStationary_matrix_3_7 <= io_mat1_3_7; // @[Muxes.scala 19:40]
    prevStationary_matrix_4_0 <= io_mat1_4_0; // @[Muxes.scala 19:40]
    prevStationary_matrix_4_1 <= io_mat1_4_1; // @[Muxes.scala 19:40]
    prevStationary_matrix_4_2 <= io_mat1_4_2; // @[Muxes.scala 19:40]
    prevStationary_matrix_4_3 <= io_mat1_4_3; // @[Muxes.scala 19:40]
    prevStationary_matrix_4_4 <= io_mat1_4_4; // @[Muxes.scala 19:40]
    prevStationary_matrix_4_5 <= io_mat1_4_5; // @[Muxes.scala 19:40]
    prevStationary_matrix_4_6 <= io_mat1_4_6; // @[Muxes.scala 19:40]
    prevStationary_matrix_4_7 <= io_mat1_4_7; // @[Muxes.scala 19:40]
    prevStationary_matrix_5_0 <= io_mat1_5_0; // @[Muxes.scala 19:40]
    prevStationary_matrix_5_1 <= io_mat1_5_1; // @[Muxes.scala 19:40]
    prevStationary_matrix_5_2 <= io_mat1_5_2; // @[Muxes.scala 19:40]
    prevStationary_matrix_5_3 <= io_mat1_5_3; // @[Muxes.scala 19:40]
    prevStationary_matrix_5_4 <= io_mat1_5_4; // @[Muxes.scala 19:40]
    prevStationary_matrix_5_5 <= io_mat1_5_5; // @[Muxes.scala 19:40]
    prevStationary_matrix_5_6 <= io_mat1_5_6; // @[Muxes.scala 19:40]
    prevStationary_matrix_5_7 <= io_mat1_5_7; // @[Muxes.scala 19:40]
    prevStationary_matrix_6_0 <= io_mat1_6_0; // @[Muxes.scala 19:40]
    prevStationary_matrix_6_1 <= io_mat1_6_1; // @[Muxes.scala 19:40]
    prevStationary_matrix_6_2 <= io_mat1_6_2; // @[Muxes.scala 19:40]
    prevStationary_matrix_6_3 <= io_mat1_6_3; // @[Muxes.scala 19:40]
    prevStationary_matrix_6_4 <= io_mat1_6_4; // @[Muxes.scala 19:40]
    prevStationary_matrix_6_5 <= io_mat1_6_5; // @[Muxes.scala 19:40]
    prevStationary_matrix_6_6 <= io_mat1_6_6; // @[Muxes.scala 19:40]
    prevStationary_matrix_6_7 <= io_mat1_6_7; // @[Muxes.scala 19:40]
    prevStationary_matrix_7_0 <= io_mat1_7_0; // @[Muxes.scala 19:40]
    prevStationary_matrix_7_1 <= io_mat1_7_1; // @[Muxes.scala 19:40]
    prevStationary_matrix_7_2 <= io_mat1_7_2; // @[Muxes.scala 19:40]
    prevStationary_matrix_7_3 <= io_mat1_7_3; // @[Muxes.scala 19:40]
    prevStationary_matrix_7_4 <= io_mat1_7_4; // @[Muxes.scala 19:40]
    prevStationary_matrix_7_5 <= io_mat1_7_5; // @[Muxes.scala 19:40]
    prevStationary_matrix_7_6 <= io_mat1_7_6; // @[Muxes.scala 19:40]
    prevStationary_matrix_7_7 <= io_mat1_7_7; // @[Muxes.scala 19:40]
    prevStreaming_matrix_0 <= io_mat2_0; // @[Muxes.scala 20:39]
    prevStreaming_matrix_1 <= io_mat2_1; // @[Muxes.scala 20:39]
    prevStreaming_matrix_2 <= io_mat2_2; // @[Muxes.scala 20:39]
    prevStreaming_matrix_3 <= io_mat2_3; // @[Muxes.scala 20:39]
    prevStreaming_matrix_4 <= io_mat2_4; // @[Muxes.scala 20:39]
    prevStreaming_matrix_5 <= io_mat2_5; // @[Muxes.scala 20:39]
    prevStreaming_matrix_6 <= io_mat2_6; // @[Muxes.scala 20:39]
    prevStreaming_matrix_7 <= io_mat2_7; // @[Muxes.scala 20:39]
    if (io_mat2_7 != prevStreaming_matrix_7) begin // @[Muxes.scala 49:51]
      matricesAreEqual <= 1'h0; // @[Muxes.scala 50:26]
    end else if (io_mat1_7_7 != prevStationary_matrix_7_7) begin // @[Muxes.scala 45:61]
      matricesAreEqual <= 1'h0; // @[Muxes.scala 46:28]
    end else if (io_mat1_7_6 != prevStationary_matrix_7_6) begin // @[Muxes.scala 45:61]
      matricesAreEqual <= 1'h0; // @[Muxes.scala 46:28]
    end else if (io_mat1_7_5 != prevStationary_matrix_7_5) begin // @[Muxes.scala 45:61]
      matricesAreEqual <= 1'h0; // @[Muxes.scala 46:28]
    end else begin
      matricesAreEqual <= _GEN_67;
    end
    if (reset) begin // @[Muxes.scala 27:25]
      jValid <= 1'h0; // @[Muxes.scala 27:25]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      if (!(j < 32'h7)) begin // @[Muxes.scala 78:40]
        jValid <= _GEN_556;
      end
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      jValid <= 1'h0; // @[Muxes.scala 93:14]
    end
    if (reset) begin // @[Muxes.scala 28:20]
      i <= 32'h0; // @[Muxes.scala 28:20]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      if (!(j < 32'h7)) begin // @[Muxes.scala 78:40]
        if (!(_T_91)) begin // @[Muxes.scala 80:83]
          i <= _GEN_555;
        end
      end
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      i <= 32'h0; // @[Muxes.scala 91:9]
    end
    if (reset) begin // @[Muxes.scala 29:20]
      j <= 32'h0; // @[Muxes.scala 29:20]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      if (j < 32'h7) begin // @[Muxes.scala 78:40]
        j <= _j_T_1; // @[Muxes.scala 79:11]
      end else if (!(_T_91)) begin // @[Muxes.scala 80:83]
        j <= 32'h0; // @[Muxes.scala 83:11]
      end
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      j <= 32'h0; // @[Muxes.scala 92:9]
    end
    if (reset) begin // @[Muxes.scala 30:20]
      k <= 32'h0; // @[Muxes.scala 30:20]
    end else if (_T_90 & _T_89) begin // @[Muxes.scala 113:76]
      k <= _k_T_1; // @[Muxes.scala 114:9]
    end
    if (reset) begin // @[Muxes.scala 31:26]
      counter <= 32'h0; // @[Muxes.scala 31:26]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      counter <= _GEN_554;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      counter <= 32'h0; // @[Muxes.scala 94:15]
    end else begin
      counter <= _GEN_554;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_0 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_0 <= _GEN_542;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_0 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_0 <= _GEN_542;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_1 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_1 <= _GEN_543;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_1 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_1 <= _GEN_543;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_2 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_2 <= _GEN_544;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_2 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_2 <= _GEN_544;
    end
    if (reset) begin // @[Muxes.scala 32:22]
      mux_3 <= 4'h0; // @[Muxes.scala 32:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      mux_3 <= _GEN_545;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      mux_3 <= 4'h0; // @[Muxes.scala 99:16]
    end else begin
      mux_3 <= _GEN_545;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_0 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_0 <= _GEN_546;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_0 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_0 <= _GEN_546;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_1 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_1 <= _GEN_547;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_1 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_1 <= _GEN_547;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_2 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_2 <= _GEN_548;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_2 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_2 <= _GEN_548;
    end
    if (reset) begin // @[Muxes.scala 33:22]
      src_3 <= 16'h0; // @[Muxes.scala 33:22]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      src_3 <= _GEN_549;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      src_3 <= 16'h0; // @[Muxes.scala 97:16]
    end else begin
      src_3 <= _GEN_549;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_0 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_0 <= _GEN_550;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_0 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_0 <= _GEN_550;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_1 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_1 <= _GEN_551;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_1 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_1 <= _GEN_551;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_2 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_2 <= _GEN_552;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_2 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_2 <= _GEN_552;
    end
    if (reset) begin // @[Muxes.scala 34:23]
      dest_3 <= 16'h0; // @[Muxes.scala 34:23]
    end else if (_T_88) begin // @[Muxes.scala 76:29]
      dest_3 <= _GEN_553;
    end else if (jValid & ~matricesAreEqual) begin // @[Muxes.scala 89:64]
      dest_3 <= 16'h0; // @[Muxes.scala 98:17]
    end else begin
      dest_3 <= _GEN_553;
    end
    if (reset) begin // @[Muxes.scala 105:24]
      jNext <= 32'h0; // @[Muxes.scala 105:24]
    end else begin
      jNext <= j; // @[Muxes.scala 106:11]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  prevStationary_matrix_0_0 = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  prevStationary_matrix_0_1 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  prevStationary_matrix_0_2 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  prevStationary_matrix_0_3 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  prevStationary_matrix_0_4 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  prevStationary_matrix_0_5 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  prevStationary_matrix_0_6 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  prevStationary_matrix_0_7 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  prevStationary_matrix_1_0 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  prevStationary_matrix_1_1 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  prevStationary_matrix_1_2 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  prevStationary_matrix_1_3 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  prevStationary_matrix_1_4 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  prevStationary_matrix_1_5 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  prevStationary_matrix_1_6 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  prevStationary_matrix_1_7 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  prevStationary_matrix_2_0 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  prevStationary_matrix_2_1 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  prevStationary_matrix_2_2 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  prevStationary_matrix_2_3 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  prevStationary_matrix_2_4 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  prevStationary_matrix_2_5 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  prevStationary_matrix_2_6 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  prevStationary_matrix_2_7 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  prevStationary_matrix_3_0 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  prevStationary_matrix_3_1 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  prevStationary_matrix_3_2 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  prevStationary_matrix_3_3 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  prevStationary_matrix_3_4 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  prevStationary_matrix_3_5 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  prevStationary_matrix_3_6 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  prevStationary_matrix_3_7 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  prevStationary_matrix_4_0 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  prevStationary_matrix_4_1 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  prevStationary_matrix_4_2 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  prevStationary_matrix_4_3 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  prevStationary_matrix_4_4 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  prevStationary_matrix_4_5 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  prevStationary_matrix_4_6 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  prevStationary_matrix_4_7 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  prevStationary_matrix_5_0 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  prevStationary_matrix_5_1 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  prevStationary_matrix_5_2 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  prevStationary_matrix_5_3 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  prevStationary_matrix_5_4 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  prevStationary_matrix_5_5 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  prevStationary_matrix_5_6 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  prevStationary_matrix_5_7 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  prevStationary_matrix_6_0 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  prevStationary_matrix_6_1 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  prevStationary_matrix_6_2 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  prevStationary_matrix_6_3 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  prevStationary_matrix_6_4 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  prevStationary_matrix_6_5 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  prevStationary_matrix_6_6 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  prevStationary_matrix_6_7 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  prevStationary_matrix_7_0 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  prevStationary_matrix_7_1 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  prevStationary_matrix_7_2 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  prevStationary_matrix_7_3 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  prevStationary_matrix_7_4 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  prevStationary_matrix_7_5 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  prevStationary_matrix_7_6 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  prevStationary_matrix_7_7 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  prevStreaming_matrix_0 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  prevStreaming_matrix_1 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  prevStreaming_matrix_2 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  prevStreaming_matrix_3 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  prevStreaming_matrix_4 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  prevStreaming_matrix_5 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  prevStreaming_matrix_6 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  prevStreaming_matrix_7 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  matricesAreEqual = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  jValid = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  i = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  j = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  k = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  counter = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  mux_0 = _RAND_78[3:0];
  _RAND_79 = {1{`RANDOM}};
  mux_1 = _RAND_79[3:0];
  _RAND_80 = {1{`RANDOM}};
  mux_2 = _RAND_80[3:0];
  _RAND_81 = {1{`RANDOM}};
  mux_3 = _RAND_81[3:0];
  _RAND_82 = {1{`RANDOM}};
  src_0 = _RAND_82[15:0];
  _RAND_83 = {1{`RANDOM}};
  src_1 = _RAND_83[15:0];
  _RAND_84 = {1{`RANDOM}};
  src_2 = _RAND_84[15:0];
  _RAND_85 = {1{`RANDOM}};
  src_3 = _RAND_85[15:0];
  _RAND_86 = {1{`RANDOM}};
  dest_0 = _RAND_86[15:0];
  _RAND_87 = {1{`RANDOM}};
  dest_1 = _RAND_87[15:0];
  _RAND_88 = {1{`RANDOM}};
  dest_2 = _RAND_88[15:0];
  _RAND_89 = {1{`RANDOM}};
  dest_3 = _RAND_89[15:0];
  _RAND_90 = {1{`RANDOM}};
  jNext = _RAND_90[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SourceDestination(
  input         clock,
  input         reset,
  input  [15:0] io_Stationary_matrix_0_0,
  input  [15:0] io_Stationary_matrix_0_1,
  input  [15:0] io_Stationary_matrix_0_2,
  input  [15:0] io_Stationary_matrix_0_3,
  input  [15:0] io_Stationary_matrix_0_4,
  input  [15:0] io_Stationary_matrix_0_5,
  input  [15:0] io_Stationary_matrix_0_6,
  input  [15:0] io_Stationary_matrix_0_7,
  input  [15:0] io_Stationary_matrix_1_0,
  input  [15:0] io_Stationary_matrix_1_1,
  input  [15:0] io_Stationary_matrix_1_2,
  input  [15:0] io_Stationary_matrix_1_3,
  input  [15:0] io_Stationary_matrix_1_4,
  input  [15:0] io_Stationary_matrix_1_5,
  input  [15:0] io_Stationary_matrix_1_6,
  input  [15:0] io_Stationary_matrix_1_7,
  input  [15:0] io_Stationary_matrix_2_0,
  input  [15:0] io_Stationary_matrix_2_1,
  input  [15:0] io_Stationary_matrix_2_2,
  input  [15:0] io_Stationary_matrix_2_3,
  input  [15:0] io_Stationary_matrix_2_4,
  input  [15:0] io_Stationary_matrix_2_5,
  input  [15:0] io_Stationary_matrix_2_6,
  input  [15:0] io_Stationary_matrix_2_7,
  input  [15:0] io_Stationary_matrix_3_0,
  input  [15:0] io_Stationary_matrix_3_1,
  input  [15:0] io_Stationary_matrix_3_2,
  input  [15:0] io_Stationary_matrix_3_3,
  input  [15:0] io_Stationary_matrix_3_4,
  input  [15:0] io_Stationary_matrix_3_5,
  input  [15:0] io_Stationary_matrix_3_6,
  input  [15:0] io_Stationary_matrix_3_7,
  input  [15:0] io_Stationary_matrix_4_0,
  input  [15:0] io_Stationary_matrix_4_1,
  input  [15:0] io_Stationary_matrix_4_2,
  input  [15:0] io_Stationary_matrix_4_3,
  input  [15:0] io_Stationary_matrix_4_4,
  input  [15:0] io_Stationary_matrix_4_5,
  input  [15:0] io_Stationary_matrix_4_6,
  input  [15:0] io_Stationary_matrix_4_7,
  input  [15:0] io_Stationary_matrix_5_0,
  input  [15:0] io_Stationary_matrix_5_1,
  input  [15:0] io_Stationary_matrix_5_2,
  input  [15:0] io_Stationary_matrix_5_3,
  input  [15:0] io_Stationary_matrix_5_4,
  input  [15:0] io_Stationary_matrix_5_5,
  input  [15:0] io_Stationary_matrix_5_6,
  input  [15:0] io_Stationary_matrix_5_7,
  input  [15:0] io_Stationary_matrix_6_0,
  input  [15:0] io_Stationary_matrix_6_1,
  input  [15:0] io_Stationary_matrix_6_2,
  input  [15:0] io_Stationary_matrix_6_3,
  input  [15:0] io_Stationary_matrix_6_4,
  input  [15:0] io_Stationary_matrix_6_5,
  input  [15:0] io_Stationary_matrix_6_6,
  input  [15:0] io_Stationary_matrix_6_7,
  input  [15:0] io_Stationary_matrix_7_0,
  input  [15:0] io_Stationary_matrix_7_1,
  input  [15:0] io_Stationary_matrix_7_2,
  input  [15:0] io_Stationary_matrix_7_3,
  input  [15:0] io_Stationary_matrix_7_4,
  input  [15:0] io_Stationary_matrix_7_5,
  input  [15:0] io_Stationary_matrix_7_6,
  input  [15:0] io_Stationary_matrix_7_7,
  input  [15:0] io_Streaming_matrix_0,
  input  [15:0] io_Streaming_matrix_1,
  input  [15:0] io_Streaming_matrix_2,
  input  [15:0] io_Streaming_matrix_3,
  input  [15:0] io_Streaming_matrix_4,
  input  [15:0] io_Streaming_matrix_5,
  input  [15:0] io_Streaming_matrix_6,
  input  [15:0] io_Streaming_matrix_7,
  output [15:0] io_counterMatrix1_bits_0_0,
  output [15:0] io_counterMatrix1_bits_0_1,
  output [15:0] io_counterMatrix1_bits_0_2,
  output [15:0] io_counterMatrix1_bits_0_3,
  output [15:0] io_counterMatrix1_bits_0_4,
  output [15:0] io_counterMatrix1_bits_0_5,
  output [15:0] io_counterMatrix1_bits_0_6,
  output [15:0] io_counterMatrix1_bits_0_7,
  output [15:0] io_counterMatrix1_bits_1_0,
  output [15:0] io_counterMatrix1_bits_1_1,
  output [15:0] io_counterMatrix1_bits_1_2,
  output [15:0] io_counterMatrix1_bits_1_3,
  output [15:0] io_counterMatrix1_bits_1_4,
  output [15:0] io_counterMatrix1_bits_1_5,
  output [15:0] io_counterMatrix1_bits_1_6,
  output [15:0] io_counterMatrix1_bits_1_7,
  output [15:0] io_counterMatrix1_bits_2_0,
  output [15:0] io_counterMatrix1_bits_2_1,
  output [15:0] io_counterMatrix1_bits_2_2,
  output [15:0] io_counterMatrix1_bits_2_3,
  output [15:0] io_counterMatrix1_bits_2_4,
  output [15:0] io_counterMatrix1_bits_2_5,
  output [15:0] io_counterMatrix1_bits_2_6,
  output [15:0] io_counterMatrix1_bits_2_7,
  output [15:0] io_counterMatrix1_bits_3_0,
  output [15:0] io_counterMatrix1_bits_3_1,
  output [15:0] io_counterMatrix1_bits_3_2,
  output [15:0] io_counterMatrix1_bits_3_3,
  output [15:0] io_counterMatrix1_bits_3_4,
  output [15:0] io_counterMatrix1_bits_3_5,
  output [15:0] io_counterMatrix1_bits_3_6,
  output [15:0] io_counterMatrix1_bits_3_7,
  output [15:0] io_counterMatrix1_bits_4_0,
  output [15:0] io_counterMatrix1_bits_4_1,
  output [15:0] io_counterMatrix1_bits_4_2,
  output [15:0] io_counterMatrix1_bits_4_3,
  output [15:0] io_counterMatrix1_bits_4_4,
  output [15:0] io_counterMatrix1_bits_4_5,
  output [15:0] io_counterMatrix1_bits_4_6,
  output [15:0] io_counterMatrix1_bits_4_7,
  output [15:0] io_counterMatrix1_bits_5_0,
  output [15:0] io_counterMatrix1_bits_5_1,
  output [15:0] io_counterMatrix1_bits_5_2,
  output [15:0] io_counterMatrix1_bits_5_3,
  output [15:0] io_counterMatrix1_bits_5_4,
  output [15:0] io_counterMatrix1_bits_5_5,
  output [15:0] io_counterMatrix1_bits_5_6,
  output [15:0] io_counterMatrix1_bits_5_7,
  output [15:0] io_counterMatrix1_bits_6_0,
  output [15:0] io_counterMatrix1_bits_6_1,
  output [15:0] io_counterMatrix1_bits_6_2,
  output [15:0] io_counterMatrix1_bits_6_3,
  output [15:0] io_counterMatrix1_bits_6_4,
  output [15:0] io_counterMatrix1_bits_6_5,
  output [15:0] io_counterMatrix1_bits_6_6,
  output [15:0] io_counterMatrix1_bits_6_7,
  output [15:0] io_counterMatrix1_bits_7_0,
  output [15:0] io_counterMatrix1_bits_7_1,
  output [15:0] io_counterMatrix1_bits_7_2,
  output [15:0] io_counterMatrix1_bits_7_3,
  output [15:0] io_counterMatrix1_bits_7_4,
  output [15:0] io_counterMatrix1_bits_7_5,
  output [15:0] io_counterMatrix1_bits_7_6,
  output [15:0] io_counterMatrix1_bits_7_7,
  output [15:0] io_counterMatrix2_bits_0,
  output [15:0] io_counterMatrix2_bits_1,
  output [15:0] io_counterMatrix2_bits_2,
  output [15:0] io_counterMatrix2_bits_3,
  output [15:0] io_counterMatrix2_bits_4,
  output [15:0] io_counterMatrix2_bits_5,
  output [15:0] io_counterMatrix2_bits_6,
  output [15:0] io_counterMatrix2_bits_7,
  output        io_valid,
  input         io_start
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
`endif // RANDOMIZE_REG_INIT
  reg [15:0] prevStationary_matrix_0_0; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_0_1; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_0_2; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_0_3; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_0_4; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_0_5; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_0_6; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_0_7; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_1_0; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_1_1; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_1_2; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_1_3; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_1_4; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_1_5; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_1_6; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_1_7; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_2_0; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_2_1; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_2_2; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_2_3; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_2_4; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_2_5; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_2_6; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_2_7; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_3_0; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_3_1; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_3_2; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_3_3; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_3_4; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_3_5; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_3_6; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_3_7; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_4_0; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_4_1; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_4_2; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_4_3; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_4_4; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_4_5; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_4_6; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_4_7; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_5_0; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_5_1; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_5_2; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_5_3; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_5_4; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_5_5; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_5_6; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_5_7; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_6_0; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_6_1; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_6_2; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_6_3; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_6_4; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_6_5; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_6_6; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_6_7; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_7_0; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_7_1; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_7_2; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_7_3; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_7_4; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_7_5; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_7_6; // @[SourceDestination.scala 15:40]
  reg [15:0] prevStationary_matrix_7_7; // @[SourceDestination.scala 15:40]
  reg  matricesAreEqual; // @[SourceDestination.scala 16:31]
  reg [15:0] counterRegs1_0_0; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_0_1; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_0_2; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_0_3; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_0_4; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_0_5; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_0_6; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_0_7; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_1_0; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_1_1; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_1_2; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_1_3; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_1_4; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_1_5; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_1_6; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_1_7; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_2_0; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_2_1; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_2_2; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_2_3; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_2_4; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_2_5; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_2_6; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_2_7; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_3_0; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_3_1; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_3_2; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_3_3; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_3_4; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_3_5; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_3_6; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_3_7; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_4_0; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_4_1; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_4_2; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_4_3; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_4_4; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_4_5; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_4_6; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_4_7; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_5_0; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_5_1; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_5_2; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_5_3; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_5_4; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_5_5; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_5_6; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_5_7; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_6_0; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_6_1; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_6_2; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_6_3; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_6_4; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_6_5; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_6_6; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_6_7; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_7_0; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_7_1; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_7_2; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_7_3; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_7_4; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_7_5; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_7_6; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs1_7_7; // @[SourceDestination.scala 17:31]
  reg [15:0] counterRegs2_0; // @[SourceDestination.scala 18:31]
  reg [15:0] counterRegs2_1; // @[SourceDestination.scala 18:31]
  reg [15:0] counterRegs2_2; // @[SourceDestination.scala 18:31]
  reg [15:0] counterRegs2_3; // @[SourceDestination.scala 18:31]
  reg [15:0] counterRegs2_4; // @[SourceDestination.scala 18:31]
  reg [15:0] counterRegs2_5; // @[SourceDestination.scala 18:31]
  reg [15:0] counterRegs2_6; // @[SourceDestination.scala 18:31]
  reg [15:0] counterRegs2_7; // @[SourceDestination.scala 18:31]
  reg [31:0] i; // @[SourceDestination.scala 20:20]
  reg [31:0] j; // @[SourceDestination.scala 21:20]
  reg  jValid; // @[SourceDestination.scala 25:21]
  reg [31:0] k; // @[SourceDestination.scala 26:20]
  reg [31:0] counter1; // @[SourceDestination.scala 28:27]
  reg [31:0] counter2; // @[SourceDestination.scala 29:27]
  wire  _reg_i_T_2 = j == 32'h7 & i == 32'h7; // @[SourceDestination.scala 31:57]
  wire  _GEN_0 = io_Stationary_matrix_0_0 != prevStationary_matrix_0_0 ? 1'h0 : 1'h1; // @[SourceDestination.scala 36:22 40:74 41:28]
  wire  _GEN_1 = io_Stationary_matrix_0_1 != prevStationary_matrix_0_1 ? 1'h0 : _GEN_0; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_2 = io_Stationary_matrix_0_2 != prevStationary_matrix_0_2 ? 1'h0 : _GEN_1; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_3 = io_Stationary_matrix_0_3 != prevStationary_matrix_0_3 ? 1'h0 : _GEN_2; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_4 = io_Stationary_matrix_0_4 != prevStationary_matrix_0_4 ? 1'h0 : _GEN_3; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_5 = io_Stationary_matrix_0_5 != prevStationary_matrix_0_5 ? 1'h0 : _GEN_4; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_6 = io_Stationary_matrix_0_6 != prevStationary_matrix_0_6 ? 1'h0 : _GEN_5; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_7 = io_Stationary_matrix_0_7 != prevStationary_matrix_0_7 ? 1'h0 : _GEN_6; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_8 = io_Stationary_matrix_1_0 != prevStationary_matrix_1_0 ? 1'h0 : _GEN_7; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_9 = io_Stationary_matrix_1_1 != prevStationary_matrix_1_1 ? 1'h0 : _GEN_8; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_10 = io_Stationary_matrix_1_2 != prevStationary_matrix_1_2 ? 1'h0 : _GEN_9; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_11 = io_Stationary_matrix_1_3 != prevStationary_matrix_1_3 ? 1'h0 : _GEN_10; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_12 = io_Stationary_matrix_1_4 != prevStationary_matrix_1_4 ? 1'h0 : _GEN_11; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_13 = io_Stationary_matrix_1_5 != prevStationary_matrix_1_5 ? 1'h0 : _GEN_12; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_14 = io_Stationary_matrix_1_6 != prevStationary_matrix_1_6 ? 1'h0 : _GEN_13; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_15 = io_Stationary_matrix_1_7 != prevStationary_matrix_1_7 ? 1'h0 : _GEN_14; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_16 = io_Stationary_matrix_2_0 != prevStationary_matrix_2_0 ? 1'h0 : _GEN_15; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_17 = io_Stationary_matrix_2_1 != prevStationary_matrix_2_1 ? 1'h0 : _GEN_16; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_18 = io_Stationary_matrix_2_2 != prevStationary_matrix_2_2 ? 1'h0 : _GEN_17; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_19 = io_Stationary_matrix_2_3 != prevStationary_matrix_2_3 ? 1'h0 : _GEN_18; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_20 = io_Stationary_matrix_2_4 != prevStationary_matrix_2_4 ? 1'h0 : _GEN_19; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_21 = io_Stationary_matrix_2_5 != prevStationary_matrix_2_5 ? 1'h0 : _GEN_20; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_22 = io_Stationary_matrix_2_6 != prevStationary_matrix_2_6 ? 1'h0 : _GEN_21; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_23 = io_Stationary_matrix_2_7 != prevStationary_matrix_2_7 ? 1'h0 : _GEN_22; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_24 = io_Stationary_matrix_3_0 != prevStationary_matrix_3_0 ? 1'h0 : _GEN_23; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_25 = io_Stationary_matrix_3_1 != prevStationary_matrix_3_1 ? 1'h0 : _GEN_24; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_26 = io_Stationary_matrix_3_2 != prevStationary_matrix_3_2 ? 1'h0 : _GEN_25; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_27 = io_Stationary_matrix_3_3 != prevStationary_matrix_3_3 ? 1'h0 : _GEN_26; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_28 = io_Stationary_matrix_3_4 != prevStationary_matrix_3_4 ? 1'h0 : _GEN_27; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_29 = io_Stationary_matrix_3_5 != prevStationary_matrix_3_5 ? 1'h0 : _GEN_28; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_30 = io_Stationary_matrix_3_6 != prevStationary_matrix_3_6 ? 1'h0 : _GEN_29; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_31 = io_Stationary_matrix_3_7 != prevStationary_matrix_3_7 ? 1'h0 : _GEN_30; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_32 = io_Stationary_matrix_4_0 != prevStationary_matrix_4_0 ? 1'h0 : _GEN_31; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_33 = io_Stationary_matrix_4_1 != prevStationary_matrix_4_1 ? 1'h0 : _GEN_32; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_34 = io_Stationary_matrix_4_2 != prevStationary_matrix_4_2 ? 1'h0 : _GEN_33; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_35 = io_Stationary_matrix_4_3 != prevStationary_matrix_4_3 ? 1'h0 : _GEN_34; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_36 = io_Stationary_matrix_4_4 != prevStationary_matrix_4_4 ? 1'h0 : _GEN_35; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_37 = io_Stationary_matrix_4_5 != prevStationary_matrix_4_5 ? 1'h0 : _GEN_36; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_38 = io_Stationary_matrix_4_6 != prevStationary_matrix_4_6 ? 1'h0 : _GEN_37; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_39 = io_Stationary_matrix_4_7 != prevStationary_matrix_4_7 ? 1'h0 : _GEN_38; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_40 = io_Stationary_matrix_5_0 != prevStationary_matrix_5_0 ? 1'h0 : _GEN_39; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_41 = io_Stationary_matrix_5_1 != prevStationary_matrix_5_1 ? 1'h0 : _GEN_40; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_42 = io_Stationary_matrix_5_2 != prevStationary_matrix_5_2 ? 1'h0 : _GEN_41; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_43 = io_Stationary_matrix_5_3 != prevStationary_matrix_5_3 ? 1'h0 : _GEN_42; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_44 = io_Stationary_matrix_5_4 != prevStationary_matrix_5_4 ? 1'h0 : _GEN_43; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_45 = io_Stationary_matrix_5_5 != prevStationary_matrix_5_5 ? 1'h0 : _GEN_44; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_46 = io_Stationary_matrix_5_6 != prevStationary_matrix_5_6 ? 1'h0 : _GEN_45; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_47 = io_Stationary_matrix_5_7 != prevStationary_matrix_5_7 ? 1'h0 : _GEN_46; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_48 = io_Stationary_matrix_6_0 != prevStationary_matrix_6_0 ? 1'h0 : _GEN_47; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_49 = io_Stationary_matrix_6_1 != prevStationary_matrix_6_1 ? 1'h0 : _GEN_48; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_50 = io_Stationary_matrix_6_2 != prevStationary_matrix_6_2 ? 1'h0 : _GEN_49; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_51 = io_Stationary_matrix_6_3 != prevStationary_matrix_6_3 ? 1'h0 : _GEN_50; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_52 = io_Stationary_matrix_6_4 != prevStationary_matrix_6_4 ? 1'h0 : _GEN_51; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_53 = io_Stationary_matrix_6_5 != prevStationary_matrix_6_5 ? 1'h0 : _GEN_52; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_54 = io_Stationary_matrix_6_6 != prevStationary_matrix_6_6 ? 1'h0 : _GEN_53; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_55 = io_Stationary_matrix_6_7 != prevStationary_matrix_6_7 ? 1'h0 : _GEN_54; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_56 = io_Stationary_matrix_7_0 != prevStationary_matrix_7_0 ? 1'h0 : _GEN_55; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_57 = io_Stationary_matrix_7_1 != prevStationary_matrix_7_1 ? 1'h0 : _GEN_56; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_58 = io_Stationary_matrix_7_2 != prevStationary_matrix_7_2 ? 1'h0 : _GEN_57; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_59 = io_Stationary_matrix_7_3 != prevStationary_matrix_7_3 ? 1'h0 : _GEN_58; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_60 = io_Stationary_matrix_7_4 != prevStationary_matrix_7_4 ? 1'h0 : _GEN_59; // @[SourceDestination.scala 40:74 41:28]
  wire  _GEN_796 = 3'h0 == i[2:0]; // @[SourceDestination.scala 53:{38,38}]
  wire  _GEN_797 = 3'h1 == j[2:0]; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_65 = 3'h0 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_0_1 : io_Stationary_matrix_0_0; // @[SourceDestination.scala 53:{38,38}]
  wire  _GEN_799 = 3'h2 == j[2:0]; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_66 = 3'h0 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_0_2 : _GEN_65; // @[SourceDestination.scala 53:{38,38}]
  wire  _GEN_801 = 3'h3 == j[2:0]; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_67 = 3'h0 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_0_3 : _GEN_66; // @[SourceDestination.scala 53:{38,38}]
  wire  _GEN_803 = 3'h4 == j[2:0]; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_68 = 3'h0 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_0_4 : _GEN_67; // @[SourceDestination.scala 53:{38,38}]
  wire  _GEN_805 = 3'h5 == j[2:0]; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_69 = 3'h0 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_0_5 : _GEN_68; // @[SourceDestination.scala 53:{38,38}]
  wire  _GEN_807 = 3'h6 == j[2:0]; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_70 = 3'h0 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_0_6 : _GEN_69; // @[SourceDestination.scala 53:{38,38}]
  wire  _GEN_809 = 3'h7 == j[2:0]; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_71 = 3'h0 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_0_7 : _GEN_70; // @[SourceDestination.scala 53:{38,38}]
  wire  _GEN_810 = 3'h1 == i[2:0]; // @[SourceDestination.scala 53:{38,38}]
  wire  _GEN_811 = 3'h0 == j[2:0]; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_72 = 3'h1 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_1_0 : _GEN_71; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_73 = 3'h1 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_1_1 : _GEN_72; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_74 = 3'h1 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_1_2 : _GEN_73; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_75 = 3'h1 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_1_3 : _GEN_74; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_76 = 3'h1 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_1_4 : _GEN_75; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_77 = 3'h1 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_1_5 : _GEN_76; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_78 = 3'h1 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_1_6 : _GEN_77; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_79 = 3'h1 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_1_7 : _GEN_78; // @[SourceDestination.scala 53:{38,38}]
  wire  _GEN_826 = 3'h2 == i[2:0]; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_80 = 3'h2 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_2_0 : _GEN_79; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_81 = 3'h2 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_2_1 : _GEN_80; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_82 = 3'h2 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_2_2 : _GEN_81; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_83 = 3'h2 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_2_3 : _GEN_82; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_84 = 3'h2 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_2_4 : _GEN_83; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_85 = 3'h2 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_2_5 : _GEN_84; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_86 = 3'h2 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_2_6 : _GEN_85; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_87 = 3'h2 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_2_7 : _GEN_86; // @[SourceDestination.scala 53:{38,38}]
  wire  _GEN_842 = 3'h3 == i[2:0]; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_88 = 3'h3 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_3_0 : _GEN_87; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_89 = 3'h3 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_3_1 : _GEN_88; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_90 = 3'h3 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_3_2 : _GEN_89; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_91 = 3'h3 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_3_3 : _GEN_90; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_92 = 3'h3 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_3_4 : _GEN_91; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_93 = 3'h3 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_3_5 : _GEN_92; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_94 = 3'h3 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_3_6 : _GEN_93; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_95 = 3'h3 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_3_7 : _GEN_94; // @[SourceDestination.scala 53:{38,38}]
  wire  _GEN_858 = 3'h4 == i[2:0]; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_96 = 3'h4 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_4_0 : _GEN_95; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_97 = 3'h4 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_4_1 : _GEN_96; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_98 = 3'h4 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_4_2 : _GEN_97; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_99 = 3'h4 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_4_3 : _GEN_98; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_100 = 3'h4 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_4_4 : _GEN_99; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_101 = 3'h4 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_4_5 : _GEN_100; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_102 = 3'h4 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_4_6 : _GEN_101; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_103 = 3'h4 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_4_7 : _GEN_102; // @[SourceDestination.scala 53:{38,38}]
  wire  _GEN_874 = 3'h5 == i[2:0]; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_104 = 3'h5 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_5_0 : _GEN_103; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_105 = 3'h5 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_5_1 : _GEN_104; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_106 = 3'h5 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_5_2 : _GEN_105; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_107 = 3'h5 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_5_3 : _GEN_106; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_108 = 3'h5 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_5_4 : _GEN_107; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_109 = 3'h5 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_5_5 : _GEN_108; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_110 = 3'h5 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_5_6 : _GEN_109; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_111 = 3'h5 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_5_7 : _GEN_110; // @[SourceDestination.scala 53:{38,38}]
  wire  _GEN_890 = 3'h6 == i[2:0]; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_112 = 3'h6 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_6_0 : _GEN_111; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_113 = 3'h6 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_6_1 : _GEN_112; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_114 = 3'h6 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_6_2 : _GEN_113; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_115 = 3'h6 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_6_3 : _GEN_114; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_116 = 3'h6 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_6_4 : _GEN_115; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_117 = 3'h6 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_6_5 : _GEN_116; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_118 = 3'h6 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_6_6 : _GEN_117; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_119 = 3'h6 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_6_7 : _GEN_118; // @[SourceDestination.scala 53:{38,38}]
  wire  _GEN_906 = 3'h7 == i[2:0]; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_120 = 3'h7 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_7_0 : _GEN_119; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_121 = 3'h7 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_7_1 : _GEN_120; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_122 = 3'h7 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_7_2 : _GEN_121; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_123 = 3'h7 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_7_3 : _GEN_122; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_124 = 3'h7 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_7_4 : _GEN_123; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_125 = 3'h7 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_7_5 : _GEN_124; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_126 = 3'h7 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_7_6 : _GEN_125; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_127 = 3'h7 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_7_7 : _GEN_126; // @[SourceDestination.scala 53:{38,38}]
  wire [15:0] _GEN_128 = _GEN_796 & _GEN_811 ? counter1[15:0] : counterRegs1_0_0; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_129 = _GEN_796 & _GEN_797 ? counter1[15:0] : counterRegs1_0_1; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_130 = _GEN_796 & _GEN_799 ? counter1[15:0] : counterRegs1_0_2; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_131 = _GEN_796 & _GEN_801 ? counter1[15:0] : counterRegs1_0_3; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_132 = _GEN_796 & _GEN_803 ? counter1[15:0] : counterRegs1_0_4; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_133 = _GEN_796 & _GEN_805 ? counter1[15:0] : counterRegs1_0_5; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_134 = _GEN_796 & _GEN_807 ? counter1[15:0] : counterRegs1_0_6; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_135 = _GEN_796 & _GEN_809 ? counter1[15:0] : counterRegs1_0_7; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_136 = _GEN_810 & _GEN_811 ? counter1[15:0] : counterRegs1_1_0; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_137 = _GEN_810 & _GEN_797 ? counter1[15:0] : counterRegs1_1_1; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_138 = _GEN_810 & _GEN_799 ? counter1[15:0] : counterRegs1_1_2; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_139 = _GEN_810 & _GEN_801 ? counter1[15:0] : counterRegs1_1_3; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_140 = _GEN_810 & _GEN_803 ? counter1[15:0] : counterRegs1_1_4; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_141 = _GEN_810 & _GEN_805 ? counter1[15:0] : counterRegs1_1_5; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_142 = _GEN_810 & _GEN_807 ? counter1[15:0] : counterRegs1_1_6; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_143 = _GEN_810 & _GEN_809 ? counter1[15:0] : counterRegs1_1_7; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_144 = _GEN_826 & _GEN_811 ? counter1[15:0] : counterRegs1_2_0; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_145 = _GEN_826 & _GEN_797 ? counter1[15:0] : counterRegs1_2_1; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_146 = _GEN_826 & _GEN_799 ? counter1[15:0] : counterRegs1_2_2; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_147 = _GEN_826 & _GEN_801 ? counter1[15:0] : counterRegs1_2_3; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_148 = _GEN_826 & _GEN_803 ? counter1[15:0] : counterRegs1_2_4; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_149 = _GEN_826 & _GEN_805 ? counter1[15:0] : counterRegs1_2_5; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_150 = _GEN_826 & _GEN_807 ? counter1[15:0] : counterRegs1_2_6; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_151 = _GEN_826 & _GEN_809 ? counter1[15:0] : counterRegs1_2_7; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_152 = _GEN_842 & _GEN_811 ? counter1[15:0] : counterRegs1_3_0; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_153 = _GEN_842 & _GEN_797 ? counter1[15:0] : counterRegs1_3_1; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_154 = _GEN_842 & _GEN_799 ? counter1[15:0] : counterRegs1_3_2; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_155 = _GEN_842 & _GEN_801 ? counter1[15:0] : counterRegs1_3_3; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_156 = _GEN_842 & _GEN_803 ? counter1[15:0] : counterRegs1_3_4; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_157 = _GEN_842 & _GEN_805 ? counter1[15:0] : counterRegs1_3_5; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_158 = _GEN_842 & _GEN_807 ? counter1[15:0] : counterRegs1_3_6; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_159 = _GEN_842 & _GEN_809 ? counter1[15:0] : counterRegs1_3_7; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_160 = _GEN_858 & _GEN_811 ? counter1[15:0] : counterRegs1_4_0; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_161 = _GEN_858 & _GEN_797 ? counter1[15:0] : counterRegs1_4_1; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_162 = _GEN_858 & _GEN_799 ? counter1[15:0] : counterRegs1_4_2; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_163 = _GEN_858 & _GEN_801 ? counter1[15:0] : counterRegs1_4_3; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_164 = _GEN_858 & _GEN_803 ? counter1[15:0] : counterRegs1_4_4; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_165 = _GEN_858 & _GEN_805 ? counter1[15:0] : counterRegs1_4_5; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_166 = _GEN_858 & _GEN_807 ? counter1[15:0] : counterRegs1_4_6; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_167 = _GEN_858 & _GEN_809 ? counter1[15:0] : counterRegs1_4_7; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_168 = _GEN_874 & _GEN_811 ? counter1[15:0] : counterRegs1_5_0; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_169 = _GEN_874 & _GEN_797 ? counter1[15:0] : counterRegs1_5_1; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_170 = _GEN_874 & _GEN_799 ? counter1[15:0] : counterRegs1_5_2; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_171 = _GEN_874 & _GEN_801 ? counter1[15:0] : counterRegs1_5_3; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_172 = _GEN_874 & _GEN_803 ? counter1[15:0] : counterRegs1_5_4; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_173 = _GEN_874 & _GEN_805 ? counter1[15:0] : counterRegs1_5_5; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_174 = _GEN_874 & _GEN_807 ? counter1[15:0] : counterRegs1_5_6; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_175 = _GEN_874 & _GEN_809 ? counter1[15:0] : counterRegs1_5_7; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_176 = _GEN_890 & _GEN_811 ? counter1[15:0] : counterRegs1_6_0; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_177 = _GEN_890 & _GEN_797 ? counter1[15:0] : counterRegs1_6_1; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_178 = _GEN_890 & _GEN_799 ? counter1[15:0] : counterRegs1_6_2; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_179 = _GEN_890 & _GEN_801 ? counter1[15:0] : counterRegs1_6_3; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_180 = _GEN_890 & _GEN_803 ? counter1[15:0] : counterRegs1_6_4; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_181 = _GEN_890 & _GEN_805 ? counter1[15:0] : counterRegs1_6_5; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_182 = _GEN_890 & _GEN_807 ? counter1[15:0] : counterRegs1_6_6; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_183 = _GEN_890 & _GEN_809 ? counter1[15:0] : counterRegs1_6_7; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_184 = _GEN_906 & _GEN_811 ? counter1[15:0] : counterRegs1_7_0; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_185 = _GEN_906 & _GEN_797 ? counter1[15:0] : counterRegs1_7_1; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_186 = _GEN_906 & _GEN_799 ? counter1[15:0] : counterRegs1_7_2; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_187 = _GEN_906 & _GEN_801 ? counter1[15:0] : counterRegs1_7_3; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_188 = _GEN_906 & _GEN_803 ? counter1[15:0] : counterRegs1_7_4; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_189 = _GEN_906 & _GEN_805 ? counter1[15:0] : counterRegs1_7_5; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_190 = _GEN_906 & _GEN_807 ? counter1[15:0] : counterRegs1_7_6; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [15:0] _GEN_191 = _GEN_906 & _GEN_809 ? counter1[15:0] : counterRegs1_7_7; // @[SourceDestination.scala 55:{28,28} 17:31]
  wire [31:0] _counter1_T_1 = counter1 + 32'h1; // @[SourceDestination.scala 57:32]
  wire [31:0] _GEN_192 = ~_reg_i_T_2 ? _counter1_T_1 : counter1; // @[SourceDestination.scala 56:83 57:20 28:27]
  wire [15:0] _GEN_193 = _GEN_796 & _GEN_811 ? 16'h1 : counterRegs1_0_0; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_194 = _GEN_796 & _GEN_797 ? 16'h1 : counterRegs1_0_1; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_195 = _GEN_796 & _GEN_799 ? 16'h1 : counterRegs1_0_2; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_196 = _GEN_796 & _GEN_801 ? 16'h1 : counterRegs1_0_3; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_197 = _GEN_796 & _GEN_803 ? 16'h1 : counterRegs1_0_4; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_198 = _GEN_796 & _GEN_805 ? 16'h1 : counterRegs1_0_5; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_199 = _GEN_796 & _GEN_807 ? 16'h1 : counterRegs1_0_6; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_200 = _GEN_796 & _GEN_809 ? 16'h1 : counterRegs1_0_7; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_201 = _GEN_810 & _GEN_811 ? 16'h1 : counterRegs1_1_0; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_202 = _GEN_810 & _GEN_797 ? 16'h1 : counterRegs1_1_1; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_203 = _GEN_810 & _GEN_799 ? 16'h1 : counterRegs1_1_2; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_204 = _GEN_810 & _GEN_801 ? 16'h1 : counterRegs1_1_3; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_205 = _GEN_810 & _GEN_803 ? 16'h1 : counterRegs1_1_4; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_206 = _GEN_810 & _GEN_805 ? 16'h1 : counterRegs1_1_5; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_207 = _GEN_810 & _GEN_807 ? 16'h1 : counterRegs1_1_6; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_208 = _GEN_810 & _GEN_809 ? 16'h1 : counterRegs1_1_7; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_209 = _GEN_826 & _GEN_811 ? 16'h1 : counterRegs1_2_0; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_210 = _GEN_826 & _GEN_797 ? 16'h1 : counterRegs1_2_1; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_211 = _GEN_826 & _GEN_799 ? 16'h1 : counterRegs1_2_2; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_212 = _GEN_826 & _GEN_801 ? 16'h1 : counterRegs1_2_3; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_213 = _GEN_826 & _GEN_803 ? 16'h1 : counterRegs1_2_4; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_214 = _GEN_826 & _GEN_805 ? 16'h1 : counterRegs1_2_5; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_215 = _GEN_826 & _GEN_807 ? 16'h1 : counterRegs1_2_6; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_216 = _GEN_826 & _GEN_809 ? 16'h1 : counterRegs1_2_7; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_217 = _GEN_842 & _GEN_811 ? 16'h1 : counterRegs1_3_0; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_218 = _GEN_842 & _GEN_797 ? 16'h1 : counterRegs1_3_1; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_219 = _GEN_842 & _GEN_799 ? 16'h1 : counterRegs1_3_2; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_220 = _GEN_842 & _GEN_801 ? 16'h1 : counterRegs1_3_3; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_221 = _GEN_842 & _GEN_803 ? 16'h1 : counterRegs1_3_4; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_222 = _GEN_842 & _GEN_805 ? 16'h1 : counterRegs1_3_5; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_223 = _GEN_842 & _GEN_807 ? 16'h1 : counterRegs1_3_6; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_224 = _GEN_842 & _GEN_809 ? 16'h1 : counterRegs1_3_7; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_225 = _GEN_858 & _GEN_811 ? 16'h1 : counterRegs1_4_0; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_226 = _GEN_858 & _GEN_797 ? 16'h1 : counterRegs1_4_1; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_227 = _GEN_858 & _GEN_799 ? 16'h1 : counterRegs1_4_2; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_228 = _GEN_858 & _GEN_801 ? 16'h1 : counterRegs1_4_3; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_229 = _GEN_858 & _GEN_803 ? 16'h1 : counterRegs1_4_4; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_230 = _GEN_858 & _GEN_805 ? 16'h1 : counterRegs1_4_5; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_231 = _GEN_858 & _GEN_807 ? 16'h1 : counterRegs1_4_6; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_232 = _GEN_858 & _GEN_809 ? 16'h1 : counterRegs1_4_7; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_233 = _GEN_874 & _GEN_811 ? 16'h1 : counterRegs1_5_0; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_234 = _GEN_874 & _GEN_797 ? 16'h1 : counterRegs1_5_1; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_235 = _GEN_874 & _GEN_799 ? 16'h1 : counterRegs1_5_2; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_236 = _GEN_874 & _GEN_801 ? 16'h1 : counterRegs1_5_3; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_237 = _GEN_874 & _GEN_803 ? 16'h1 : counterRegs1_5_4; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_238 = _GEN_874 & _GEN_805 ? 16'h1 : counterRegs1_5_5; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_239 = _GEN_874 & _GEN_807 ? 16'h1 : counterRegs1_5_6; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_240 = _GEN_874 & _GEN_809 ? 16'h1 : counterRegs1_5_7; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_241 = _GEN_890 & _GEN_811 ? 16'h1 : counterRegs1_6_0; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_242 = _GEN_890 & _GEN_797 ? 16'h1 : counterRegs1_6_1; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_243 = _GEN_890 & _GEN_799 ? 16'h1 : counterRegs1_6_2; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_244 = _GEN_890 & _GEN_801 ? 16'h1 : counterRegs1_6_3; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_245 = _GEN_890 & _GEN_803 ? 16'h1 : counterRegs1_6_4; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_246 = _GEN_890 & _GEN_805 ? 16'h1 : counterRegs1_6_5; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_247 = _GEN_890 & _GEN_807 ? 16'h1 : counterRegs1_6_6; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_248 = _GEN_890 & _GEN_809 ? 16'h1 : counterRegs1_6_7; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_249 = _GEN_906 & _GEN_811 ? 16'h1 : counterRegs1_7_0; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_250 = _GEN_906 & _GEN_797 ? 16'h1 : counterRegs1_7_1; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_251 = _GEN_906 & _GEN_799 ? 16'h1 : counterRegs1_7_2; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_252 = _GEN_906 & _GEN_801 ? 16'h1 : counterRegs1_7_3; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_253 = _GEN_906 & _GEN_803 ? 16'h1 : counterRegs1_7_4; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_254 = _GEN_906 & _GEN_805 ? 16'h1 : counterRegs1_7_5; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_255 = _GEN_906 & _GEN_807 ? 16'h1 : counterRegs1_7_6; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_256 = _GEN_906 & _GEN_809 ? 16'h1 : counterRegs1_7_7; // @[SourceDestination.scala 60:{28,28} 17:31]
  wire [15:0] _GEN_257 = counter1 < 32'h5 ? _GEN_128 : _GEN_193; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_258 = counter1 < 32'h5 ? _GEN_129 : _GEN_194; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_259 = counter1 < 32'h5 ? _GEN_130 : _GEN_195; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_260 = counter1 < 32'h5 ? _GEN_131 : _GEN_196; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_261 = counter1 < 32'h5 ? _GEN_132 : _GEN_197; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_262 = counter1 < 32'h5 ? _GEN_133 : _GEN_198; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_263 = counter1 < 32'h5 ? _GEN_134 : _GEN_199; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_264 = counter1 < 32'h5 ? _GEN_135 : _GEN_200; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_265 = counter1 < 32'h5 ? _GEN_136 : _GEN_201; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_266 = counter1 < 32'h5 ? _GEN_137 : _GEN_202; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_267 = counter1 < 32'h5 ? _GEN_138 : _GEN_203; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_268 = counter1 < 32'h5 ? _GEN_139 : _GEN_204; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_269 = counter1 < 32'h5 ? _GEN_140 : _GEN_205; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_270 = counter1 < 32'h5 ? _GEN_141 : _GEN_206; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_271 = counter1 < 32'h5 ? _GEN_142 : _GEN_207; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_272 = counter1 < 32'h5 ? _GEN_143 : _GEN_208; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_273 = counter1 < 32'h5 ? _GEN_144 : _GEN_209; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_274 = counter1 < 32'h5 ? _GEN_145 : _GEN_210; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_275 = counter1 < 32'h5 ? _GEN_146 : _GEN_211; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_276 = counter1 < 32'h5 ? _GEN_147 : _GEN_212; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_277 = counter1 < 32'h5 ? _GEN_148 : _GEN_213; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_278 = counter1 < 32'h5 ? _GEN_149 : _GEN_214; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_279 = counter1 < 32'h5 ? _GEN_150 : _GEN_215; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_280 = counter1 < 32'h5 ? _GEN_151 : _GEN_216; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_281 = counter1 < 32'h5 ? _GEN_152 : _GEN_217; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_282 = counter1 < 32'h5 ? _GEN_153 : _GEN_218; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_283 = counter1 < 32'h5 ? _GEN_154 : _GEN_219; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_284 = counter1 < 32'h5 ? _GEN_155 : _GEN_220; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_285 = counter1 < 32'h5 ? _GEN_156 : _GEN_221; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_286 = counter1 < 32'h5 ? _GEN_157 : _GEN_222; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_287 = counter1 < 32'h5 ? _GEN_158 : _GEN_223; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_288 = counter1 < 32'h5 ? _GEN_159 : _GEN_224; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_289 = counter1 < 32'h5 ? _GEN_160 : _GEN_225; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_290 = counter1 < 32'h5 ? _GEN_161 : _GEN_226; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_291 = counter1 < 32'h5 ? _GEN_162 : _GEN_227; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_292 = counter1 < 32'h5 ? _GEN_163 : _GEN_228; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_293 = counter1 < 32'h5 ? _GEN_164 : _GEN_229; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_294 = counter1 < 32'h5 ? _GEN_165 : _GEN_230; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_295 = counter1 < 32'h5 ? _GEN_166 : _GEN_231; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_296 = counter1 < 32'h5 ? _GEN_167 : _GEN_232; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_297 = counter1 < 32'h5 ? _GEN_168 : _GEN_233; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_298 = counter1 < 32'h5 ? _GEN_169 : _GEN_234; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_299 = counter1 < 32'h5 ? _GEN_170 : _GEN_235; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_300 = counter1 < 32'h5 ? _GEN_171 : _GEN_236; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_301 = counter1 < 32'h5 ? _GEN_172 : _GEN_237; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_302 = counter1 < 32'h5 ? _GEN_173 : _GEN_238; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_303 = counter1 < 32'h5 ? _GEN_174 : _GEN_239; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_304 = counter1 < 32'h5 ? _GEN_175 : _GEN_240; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_305 = counter1 < 32'h5 ? _GEN_176 : _GEN_241; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_306 = counter1 < 32'h5 ? _GEN_177 : _GEN_242; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_307 = counter1 < 32'h5 ? _GEN_178 : _GEN_243; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_308 = counter1 < 32'h5 ? _GEN_179 : _GEN_244; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_309 = counter1 < 32'h5 ? _GEN_180 : _GEN_245; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_310 = counter1 < 32'h5 ? _GEN_181 : _GEN_246; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_311 = counter1 < 32'h5 ? _GEN_182 : _GEN_247; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_312 = counter1 < 32'h5 ? _GEN_183 : _GEN_248; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_313 = counter1 < 32'h5 ? _GEN_184 : _GEN_249; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_314 = counter1 < 32'h5 ? _GEN_185 : _GEN_250; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_315 = counter1 < 32'h5 ? _GEN_186 : _GEN_251; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_316 = counter1 < 32'h5 ? _GEN_187 : _GEN_252; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_317 = counter1 < 32'h5 ? _GEN_188 : _GEN_253; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_318 = counter1 < 32'h5 ? _GEN_189 : _GEN_254; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_319 = counter1 < 32'h5 ? _GEN_190 : _GEN_255; // @[SourceDestination.scala 54:48]
  wire [15:0] _GEN_320 = counter1 < 32'h5 ? _GEN_191 : _GEN_256; // @[SourceDestination.scala 54:48]
  wire [31:0] _GEN_321 = counter1 < 32'h5 ? _GEN_192 : 32'h2; // @[SourceDestination.scala 54:48 61:18]
  wire [15:0] _GEN_322 = _GEN_796 & _GEN_811 ? 16'h0 : counterRegs1_0_0; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_323 = _GEN_796 & _GEN_797 ? 16'h0 : counterRegs1_0_1; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_324 = _GEN_796 & _GEN_799 ? 16'h0 : counterRegs1_0_2; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_325 = _GEN_796 & _GEN_801 ? 16'h0 : counterRegs1_0_3; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_326 = _GEN_796 & _GEN_803 ? 16'h0 : counterRegs1_0_4; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_327 = _GEN_796 & _GEN_805 ? 16'h0 : counterRegs1_0_5; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_328 = _GEN_796 & _GEN_807 ? 16'h0 : counterRegs1_0_6; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_329 = _GEN_796 & _GEN_809 ? 16'h0 : counterRegs1_0_7; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_330 = _GEN_810 & _GEN_811 ? 16'h0 : counterRegs1_1_0; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_331 = _GEN_810 & _GEN_797 ? 16'h0 : counterRegs1_1_1; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_332 = _GEN_810 & _GEN_799 ? 16'h0 : counterRegs1_1_2; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_333 = _GEN_810 & _GEN_801 ? 16'h0 : counterRegs1_1_3; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_334 = _GEN_810 & _GEN_803 ? 16'h0 : counterRegs1_1_4; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_335 = _GEN_810 & _GEN_805 ? 16'h0 : counterRegs1_1_5; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_336 = _GEN_810 & _GEN_807 ? 16'h0 : counterRegs1_1_6; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_337 = _GEN_810 & _GEN_809 ? 16'h0 : counterRegs1_1_7; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_338 = _GEN_826 & _GEN_811 ? 16'h0 : counterRegs1_2_0; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_339 = _GEN_826 & _GEN_797 ? 16'h0 : counterRegs1_2_1; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_340 = _GEN_826 & _GEN_799 ? 16'h0 : counterRegs1_2_2; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_341 = _GEN_826 & _GEN_801 ? 16'h0 : counterRegs1_2_3; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_342 = _GEN_826 & _GEN_803 ? 16'h0 : counterRegs1_2_4; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_343 = _GEN_826 & _GEN_805 ? 16'h0 : counterRegs1_2_5; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_344 = _GEN_826 & _GEN_807 ? 16'h0 : counterRegs1_2_6; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_345 = _GEN_826 & _GEN_809 ? 16'h0 : counterRegs1_2_7; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_346 = _GEN_842 & _GEN_811 ? 16'h0 : counterRegs1_3_0; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_347 = _GEN_842 & _GEN_797 ? 16'h0 : counterRegs1_3_1; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_348 = _GEN_842 & _GEN_799 ? 16'h0 : counterRegs1_3_2; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_349 = _GEN_842 & _GEN_801 ? 16'h0 : counterRegs1_3_3; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_350 = _GEN_842 & _GEN_803 ? 16'h0 : counterRegs1_3_4; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_351 = _GEN_842 & _GEN_805 ? 16'h0 : counterRegs1_3_5; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_352 = _GEN_842 & _GEN_807 ? 16'h0 : counterRegs1_3_6; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_353 = _GEN_842 & _GEN_809 ? 16'h0 : counterRegs1_3_7; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_354 = _GEN_858 & _GEN_811 ? 16'h0 : counterRegs1_4_0; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_355 = _GEN_858 & _GEN_797 ? 16'h0 : counterRegs1_4_1; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_356 = _GEN_858 & _GEN_799 ? 16'h0 : counterRegs1_4_2; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_357 = _GEN_858 & _GEN_801 ? 16'h0 : counterRegs1_4_3; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_358 = _GEN_858 & _GEN_803 ? 16'h0 : counterRegs1_4_4; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_359 = _GEN_858 & _GEN_805 ? 16'h0 : counterRegs1_4_5; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_360 = _GEN_858 & _GEN_807 ? 16'h0 : counterRegs1_4_6; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_361 = _GEN_858 & _GEN_809 ? 16'h0 : counterRegs1_4_7; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_362 = _GEN_874 & _GEN_811 ? 16'h0 : counterRegs1_5_0; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_363 = _GEN_874 & _GEN_797 ? 16'h0 : counterRegs1_5_1; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_364 = _GEN_874 & _GEN_799 ? 16'h0 : counterRegs1_5_2; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_365 = _GEN_874 & _GEN_801 ? 16'h0 : counterRegs1_5_3; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_366 = _GEN_874 & _GEN_803 ? 16'h0 : counterRegs1_5_4; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_367 = _GEN_874 & _GEN_805 ? 16'h0 : counterRegs1_5_5; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_368 = _GEN_874 & _GEN_807 ? 16'h0 : counterRegs1_5_6; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_369 = _GEN_874 & _GEN_809 ? 16'h0 : counterRegs1_5_7; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_370 = _GEN_890 & _GEN_811 ? 16'h0 : counterRegs1_6_0; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_371 = _GEN_890 & _GEN_797 ? 16'h0 : counterRegs1_6_1; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_372 = _GEN_890 & _GEN_799 ? 16'h0 : counterRegs1_6_2; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_373 = _GEN_890 & _GEN_801 ? 16'h0 : counterRegs1_6_3; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_374 = _GEN_890 & _GEN_803 ? 16'h0 : counterRegs1_6_4; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_375 = _GEN_890 & _GEN_805 ? 16'h0 : counterRegs1_6_5; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_376 = _GEN_890 & _GEN_807 ? 16'h0 : counterRegs1_6_6; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_377 = _GEN_890 & _GEN_809 ? 16'h0 : counterRegs1_6_7; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_378 = _GEN_906 & _GEN_811 ? 16'h0 : counterRegs1_7_0; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_379 = _GEN_906 & _GEN_797 ? 16'h0 : counterRegs1_7_1; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_380 = _GEN_906 & _GEN_799 ? 16'h0 : counterRegs1_7_2; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_381 = _GEN_906 & _GEN_801 ? 16'h0 : counterRegs1_7_3; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_382 = _GEN_906 & _GEN_803 ? 16'h0 : counterRegs1_7_4; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_383 = _GEN_906 & _GEN_805 ? 16'h0 : counterRegs1_7_5; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_384 = _GEN_906 & _GEN_807 ? 16'h0 : counterRegs1_7_6; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_385 = _GEN_906 & _GEN_809 ? 16'h0 : counterRegs1_7_7; // @[SourceDestination.scala 64:{26,26} 17:31]
  wire [15:0] _GEN_386 = _GEN_127 != 16'h0 ? _GEN_257 : _GEN_322; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_387 = _GEN_127 != 16'h0 ? _GEN_258 : _GEN_323; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_388 = _GEN_127 != 16'h0 ? _GEN_259 : _GEN_324; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_389 = _GEN_127 != 16'h0 ? _GEN_260 : _GEN_325; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_390 = _GEN_127 != 16'h0 ? _GEN_261 : _GEN_326; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_391 = _GEN_127 != 16'h0 ? _GEN_262 : _GEN_327; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_392 = _GEN_127 != 16'h0 ? _GEN_263 : _GEN_328; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_393 = _GEN_127 != 16'h0 ? _GEN_264 : _GEN_329; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_394 = _GEN_127 != 16'h0 ? _GEN_265 : _GEN_330; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_395 = _GEN_127 != 16'h0 ? _GEN_266 : _GEN_331; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_396 = _GEN_127 != 16'h0 ? _GEN_267 : _GEN_332; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_397 = _GEN_127 != 16'h0 ? _GEN_268 : _GEN_333; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_398 = _GEN_127 != 16'h0 ? _GEN_269 : _GEN_334; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_399 = _GEN_127 != 16'h0 ? _GEN_270 : _GEN_335; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_400 = _GEN_127 != 16'h0 ? _GEN_271 : _GEN_336; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_401 = _GEN_127 != 16'h0 ? _GEN_272 : _GEN_337; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_402 = _GEN_127 != 16'h0 ? _GEN_273 : _GEN_338; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_403 = _GEN_127 != 16'h0 ? _GEN_274 : _GEN_339; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_404 = _GEN_127 != 16'h0 ? _GEN_275 : _GEN_340; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_405 = _GEN_127 != 16'h0 ? _GEN_276 : _GEN_341; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_406 = _GEN_127 != 16'h0 ? _GEN_277 : _GEN_342; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_407 = _GEN_127 != 16'h0 ? _GEN_278 : _GEN_343; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_408 = _GEN_127 != 16'h0 ? _GEN_279 : _GEN_344; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_409 = _GEN_127 != 16'h0 ? _GEN_280 : _GEN_345; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_410 = _GEN_127 != 16'h0 ? _GEN_281 : _GEN_346; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_411 = _GEN_127 != 16'h0 ? _GEN_282 : _GEN_347; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_412 = _GEN_127 != 16'h0 ? _GEN_283 : _GEN_348; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_413 = _GEN_127 != 16'h0 ? _GEN_284 : _GEN_349; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_414 = _GEN_127 != 16'h0 ? _GEN_285 : _GEN_350; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_415 = _GEN_127 != 16'h0 ? _GEN_286 : _GEN_351; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_416 = _GEN_127 != 16'h0 ? _GEN_287 : _GEN_352; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_417 = _GEN_127 != 16'h0 ? _GEN_288 : _GEN_353; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_418 = _GEN_127 != 16'h0 ? _GEN_289 : _GEN_354; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_419 = _GEN_127 != 16'h0 ? _GEN_290 : _GEN_355; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_420 = _GEN_127 != 16'h0 ? _GEN_291 : _GEN_356; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_421 = _GEN_127 != 16'h0 ? _GEN_292 : _GEN_357; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_422 = _GEN_127 != 16'h0 ? _GEN_293 : _GEN_358; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_423 = _GEN_127 != 16'h0 ? _GEN_294 : _GEN_359; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_424 = _GEN_127 != 16'h0 ? _GEN_295 : _GEN_360; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_425 = _GEN_127 != 16'h0 ? _GEN_296 : _GEN_361; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_426 = _GEN_127 != 16'h0 ? _GEN_297 : _GEN_362; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_427 = _GEN_127 != 16'h0 ? _GEN_298 : _GEN_363; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_428 = _GEN_127 != 16'h0 ? _GEN_299 : _GEN_364; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_429 = _GEN_127 != 16'h0 ? _GEN_300 : _GEN_365; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_430 = _GEN_127 != 16'h0 ? _GEN_301 : _GEN_366; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_431 = _GEN_127 != 16'h0 ? _GEN_302 : _GEN_367; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_432 = _GEN_127 != 16'h0 ? _GEN_303 : _GEN_368; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_433 = _GEN_127 != 16'h0 ? _GEN_304 : _GEN_369; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_434 = _GEN_127 != 16'h0 ? _GEN_305 : _GEN_370; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_435 = _GEN_127 != 16'h0 ? _GEN_306 : _GEN_371; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_436 = _GEN_127 != 16'h0 ? _GEN_307 : _GEN_372; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_437 = _GEN_127 != 16'h0 ? _GEN_308 : _GEN_373; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_438 = _GEN_127 != 16'h0 ? _GEN_309 : _GEN_374; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_439 = _GEN_127 != 16'h0 ? _GEN_310 : _GEN_375; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_440 = _GEN_127 != 16'h0 ? _GEN_311 : _GEN_376; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_441 = _GEN_127 != 16'h0 ? _GEN_312 : _GEN_377; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_442 = _GEN_127 != 16'h0 ? _GEN_313 : _GEN_378; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_443 = _GEN_127 != 16'h0 ? _GEN_314 : _GEN_379; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_444 = _GEN_127 != 16'h0 ? _GEN_315 : _GEN_380; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_445 = _GEN_127 != 16'h0 ? _GEN_316 : _GEN_381; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_446 = _GEN_127 != 16'h0 ? _GEN_317 : _GEN_382; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_447 = _GEN_127 != 16'h0 ? _GEN_318 : _GEN_383; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_448 = _GEN_127 != 16'h0 ? _GEN_319 : _GEN_384; // @[SourceDestination.scala 53:47]
  wire [15:0] _GEN_449 = _GEN_127 != 16'h0 ? _GEN_320 : _GEN_385; // @[SourceDestination.scala 53:47]
  wire [31:0] _GEN_450 = _GEN_127 != 16'h0 ? _GEN_321 : counter1; // @[SourceDestination.scala 28:27 53:47]
  wire [15:0] _GEN_452 = 3'h1 == k[2:0] ? io_Streaming_matrix_1 : io_Streaming_matrix_0; // @[SourceDestination.scala 67:{34,34}]
  wire [15:0] _GEN_453 = 3'h2 == k[2:0] ? io_Streaming_matrix_2 : _GEN_452; // @[SourceDestination.scala 67:{34,34}]
  wire [15:0] _GEN_454 = 3'h3 == k[2:0] ? io_Streaming_matrix_3 : _GEN_453; // @[SourceDestination.scala 67:{34,34}]
  wire [15:0] _GEN_455 = 3'h4 == k[2:0] ? io_Streaming_matrix_4 : _GEN_454; // @[SourceDestination.scala 67:{34,34}]
  wire [15:0] _GEN_456 = 3'h5 == k[2:0] ? io_Streaming_matrix_5 : _GEN_455; // @[SourceDestination.scala 67:{34,34}]
  wire [15:0] _GEN_457 = 3'h6 == k[2:0] ? io_Streaming_matrix_6 : _GEN_456; // @[SourceDestination.scala 67:{34,34}]
  wire [15:0] _GEN_458 = 3'h7 == k[2:0] ? io_Streaming_matrix_7 : _GEN_457; // @[SourceDestination.scala 67:{34,34}]
  wire [15:0] _GEN_459 = 3'h0 == k[2:0] ? counter2[15:0] : counterRegs2_0; // @[SourceDestination.scala 68:{23,23} 18:31]
  wire [15:0] _GEN_460 = 3'h1 == k[2:0] ? counter2[15:0] : counterRegs2_1; // @[SourceDestination.scala 68:{23,23} 18:31]
  wire [15:0] _GEN_461 = 3'h2 == k[2:0] ? counter2[15:0] : counterRegs2_2; // @[SourceDestination.scala 68:{23,23} 18:31]
  wire [15:0] _GEN_462 = 3'h3 == k[2:0] ? counter2[15:0] : counterRegs2_3; // @[SourceDestination.scala 68:{23,23} 18:31]
  wire [15:0] _GEN_463 = 3'h4 == k[2:0] ? counter2[15:0] : counterRegs2_4; // @[SourceDestination.scala 68:{23,23} 18:31]
  wire [15:0] _GEN_464 = 3'h5 == k[2:0] ? counter2[15:0] : counterRegs2_5; // @[SourceDestination.scala 68:{23,23} 18:31]
  wire [15:0] _GEN_465 = 3'h6 == k[2:0] ? counter2[15:0] : counterRegs2_6; // @[SourceDestination.scala 68:{23,23} 18:31]
  wire [15:0] _GEN_466 = 3'h7 == k[2:0] ? counter2[15:0] : counterRegs2_7; // @[SourceDestination.scala 68:{23,23} 18:31]
  wire [31:0] _counter2_T_1 = counter2 + 32'h1; // @[SourceDestination.scala 69:28]
  wire [15:0] _GEN_467 = _GEN_458 != 16'h0 ? _GEN_459 : counterRegs2_0; // @[SourceDestination.scala 18:31 67:43]
  wire [15:0] _GEN_468 = _GEN_458 != 16'h0 ? _GEN_460 : counterRegs2_1; // @[SourceDestination.scala 18:31 67:43]
  wire [15:0] _GEN_469 = _GEN_458 != 16'h0 ? _GEN_461 : counterRegs2_2; // @[SourceDestination.scala 18:31 67:43]
  wire [15:0] _GEN_470 = _GEN_458 != 16'h0 ? _GEN_462 : counterRegs2_3; // @[SourceDestination.scala 18:31 67:43]
  wire [15:0] _GEN_471 = _GEN_458 != 16'h0 ? _GEN_463 : counterRegs2_4; // @[SourceDestination.scala 18:31 67:43]
  wire [15:0] _GEN_472 = _GEN_458 != 16'h0 ? _GEN_464 : counterRegs2_5; // @[SourceDestination.scala 18:31 67:43]
  wire [15:0] _GEN_473 = _GEN_458 != 16'h0 ? _GEN_465 : counterRegs2_6; // @[SourceDestination.scala 18:31 67:43]
  wire [15:0] _GEN_474 = _GEN_458 != 16'h0 ? _GEN_466 : counterRegs2_7; // @[SourceDestination.scala 18:31 67:43]
  wire [31:0] _GEN_475 = _GEN_458 != 16'h0 ? _counter2_T_1 : counter2; // @[SourceDestination.scala 67:43 69:16 29:27]
  wire [31:0] _k_T_1 = k + 32'h1; // @[SourceDestination.scala 77:16]
  wire [31:0] _GEN_477 = k == 32'h7 ? k : _k_T_1; // @[SourceDestination.scala 73:37 74:9]
  wire [31:0] _GEN_478 = k == 32'h7 ? counter2 : _GEN_475; // @[SourceDestination.scala 73:37 75:16]
  wire [31:0] _j_T_1 = j + 32'h1; // @[SourceDestination.scala 81:16]
  wire [31:0] _i_T_1 = i + 32'h1; // @[SourceDestination.scala 87:18]
  wire [31:0] _GEN_479 = i < 32'h7 ? _i_T_1 : i; // @[SourceDestination.scala 86:42 87:13 20:20]
  wire [31:0] _GEN_481 = _reg_i_T_2 ? j : 32'h0; // @[SourceDestination.scala 21:20 82:83 85:11]
  wire [31:0] _GEN_482 = _reg_i_T_2 ? i : _GEN_479; // @[SourceDestination.scala 20:20 82:83]
  wire  _GEN_484 = j < 32'h7 ? 1'h0 : _reg_i_T_2; // @[SourceDestination.scala 49:12 80:40]
  wire  _GEN_564 = ~jValid & _GEN_484; // @[SourceDestination.scala 49:12 79:26]
  wire [31:0] _GEN_724 = io_start ? {{16'd0}, counterRegs1_0_0} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_725 = io_start ? {{16'd0}, counterRegs1_0_1} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_726 = io_start ? {{16'd0}, counterRegs1_0_2} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_727 = io_start ? {{16'd0}, counterRegs1_0_3} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_728 = io_start ? {{16'd0}, counterRegs1_0_4} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_729 = io_start ? {{16'd0}, counterRegs1_0_5} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_730 = io_start ? {{16'd0}, counterRegs1_0_6} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_731 = io_start ? {{16'd0}, counterRegs1_0_7} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_732 = io_start ? {{16'd0}, counterRegs1_1_0} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_733 = io_start ? {{16'd0}, counterRegs1_1_1} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_734 = io_start ? {{16'd0}, counterRegs1_1_2} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_735 = io_start ? {{16'd0}, counterRegs1_1_3} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_736 = io_start ? {{16'd0}, counterRegs1_1_4} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_737 = io_start ? {{16'd0}, counterRegs1_1_5} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_738 = io_start ? {{16'd0}, counterRegs1_1_6} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_739 = io_start ? {{16'd0}, counterRegs1_1_7} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_740 = io_start ? {{16'd0}, counterRegs1_2_0} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_741 = io_start ? {{16'd0}, counterRegs1_2_1} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_742 = io_start ? {{16'd0}, counterRegs1_2_2} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_743 = io_start ? {{16'd0}, counterRegs1_2_3} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_744 = io_start ? {{16'd0}, counterRegs1_2_4} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_745 = io_start ? {{16'd0}, counterRegs1_2_5} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_746 = io_start ? {{16'd0}, counterRegs1_2_6} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_747 = io_start ? {{16'd0}, counterRegs1_2_7} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_748 = io_start ? {{16'd0}, counterRegs1_3_0} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_749 = io_start ? {{16'd0}, counterRegs1_3_1} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_750 = io_start ? {{16'd0}, counterRegs1_3_2} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_751 = io_start ? {{16'd0}, counterRegs1_3_3} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_752 = io_start ? {{16'd0}, counterRegs1_3_4} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_753 = io_start ? {{16'd0}, counterRegs1_3_5} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_754 = io_start ? {{16'd0}, counterRegs1_3_6} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_755 = io_start ? {{16'd0}, counterRegs1_3_7} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_756 = io_start ? {{16'd0}, counterRegs1_4_0} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_757 = io_start ? {{16'd0}, counterRegs1_4_1} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_758 = io_start ? {{16'd0}, counterRegs1_4_2} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_759 = io_start ? {{16'd0}, counterRegs1_4_3} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_760 = io_start ? {{16'd0}, counterRegs1_4_4} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_761 = io_start ? {{16'd0}, counterRegs1_4_5} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_762 = io_start ? {{16'd0}, counterRegs1_4_6} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_763 = io_start ? {{16'd0}, counterRegs1_4_7} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_764 = io_start ? {{16'd0}, counterRegs1_5_0} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_765 = io_start ? {{16'd0}, counterRegs1_5_1} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_766 = io_start ? {{16'd0}, counterRegs1_5_2} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_767 = io_start ? {{16'd0}, counterRegs1_5_3} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_768 = io_start ? {{16'd0}, counterRegs1_5_4} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_769 = io_start ? {{16'd0}, counterRegs1_5_5} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_770 = io_start ? {{16'd0}, counterRegs1_5_6} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_771 = io_start ? {{16'd0}, counterRegs1_5_7} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_772 = io_start ? {{16'd0}, counterRegs1_6_0} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_773 = io_start ? {{16'd0}, counterRegs1_6_1} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_774 = io_start ? {{16'd0}, counterRegs1_6_2} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_775 = io_start ? {{16'd0}, counterRegs1_6_3} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_776 = io_start ? {{16'd0}, counterRegs1_6_4} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_777 = io_start ? {{16'd0}, counterRegs1_6_5} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_778 = io_start ? {{16'd0}, counterRegs1_6_6} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_779 = io_start ? {{16'd0}, counterRegs1_6_7} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_780 = io_start ? {{16'd0}, counterRegs1_7_0} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_781 = io_start ? {{16'd0}, counterRegs1_7_1} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_782 = io_start ? {{16'd0}, counterRegs1_7_2} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_783 = io_start ? {{16'd0}, counterRegs1_7_3} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_784 = io_start ? {{16'd0}, counterRegs1_7_4} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_785 = io_start ? {{16'd0}, counterRegs1_7_5} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_786 = io_start ? {{16'd0}, counterRegs1_7_6} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_787 = io_start ? {{16'd0}, counterRegs1_7_7} : 32'h0; // @[SourceDestination.scala 34:17 114:28 118:26]
  wire [31:0] _GEN_788 = io_start ? {{16'd0}, counterRegs2_0} : 32'h0; // @[SourceDestination.scala 34:17 115:28 119:26]
  wire [31:0] _GEN_789 = io_start ? {{16'd0}, counterRegs2_1} : 32'h0; // @[SourceDestination.scala 34:17 115:28 119:26]
  wire [31:0] _GEN_790 = io_start ? {{16'd0}, counterRegs2_2} : 32'h0; // @[SourceDestination.scala 34:17 115:28 119:26]
  wire [31:0] _GEN_791 = io_start ? {{16'd0}, counterRegs2_3} : 32'h0; // @[SourceDestination.scala 34:17 115:28 119:26]
  wire [31:0] _GEN_792 = io_start ? {{16'd0}, counterRegs2_4} : 32'h0; // @[SourceDestination.scala 34:17 115:28 119:26]
  wire [31:0] _GEN_793 = io_start ? {{16'd0}, counterRegs2_5} : 32'h0; // @[SourceDestination.scala 34:17 115:28 119:26]
  wire [31:0] _GEN_794 = io_start ? {{16'd0}, counterRegs2_6} : 32'h0; // @[SourceDestination.scala 34:17 115:28 119:26]
  wire [31:0] _GEN_795 = io_start ? {{16'd0}, counterRegs2_7} : 32'h0; // @[SourceDestination.scala 34:17 115:28 119:26]
  assign io_counterMatrix1_bits_0_0 = _GEN_724[15:0];
  assign io_counterMatrix1_bits_0_1 = _GEN_725[15:0];
  assign io_counterMatrix1_bits_0_2 = _GEN_726[15:0];
  assign io_counterMatrix1_bits_0_3 = _GEN_727[15:0];
  assign io_counterMatrix1_bits_0_4 = _GEN_728[15:0];
  assign io_counterMatrix1_bits_0_5 = _GEN_729[15:0];
  assign io_counterMatrix1_bits_0_6 = _GEN_730[15:0];
  assign io_counterMatrix1_bits_0_7 = _GEN_731[15:0];
  assign io_counterMatrix1_bits_1_0 = _GEN_732[15:0];
  assign io_counterMatrix1_bits_1_1 = _GEN_733[15:0];
  assign io_counterMatrix1_bits_1_2 = _GEN_734[15:0];
  assign io_counterMatrix1_bits_1_3 = _GEN_735[15:0];
  assign io_counterMatrix1_bits_1_4 = _GEN_736[15:0];
  assign io_counterMatrix1_bits_1_5 = _GEN_737[15:0];
  assign io_counterMatrix1_bits_1_6 = _GEN_738[15:0];
  assign io_counterMatrix1_bits_1_7 = _GEN_739[15:0];
  assign io_counterMatrix1_bits_2_0 = _GEN_740[15:0];
  assign io_counterMatrix1_bits_2_1 = _GEN_741[15:0];
  assign io_counterMatrix1_bits_2_2 = _GEN_742[15:0];
  assign io_counterMatrix1_bits_2_3 = _GEN_743[15:0];
  assign io_counterMatrix1_bits_2_4 = _GEN_744[15:0];
  assign io_counterMatrix1_bits_2_5 = _GEN_745[15:0];
  assign io_counterMatrix1_bits_2_6 = _GEN_746[15:0];
  assign io_counterMatrix1_bits_2_7 = _GEN_747[15:0];
  assign io_counterMatrix1_bits_3_0 = _GEN_748[15:0];
  assign io_counterMatrix1_bits_3_1 = _GEN_749[15:0];
  assign io_counterMatrix1_bits_3_2 = _GEN_750[15:0];
  assign io_counterMatrix1_bits_3_3 = _GEN_751[15:0];
  assign io_counterMatrix1_bits_3_4 = _GEN_752[15:0];
  assign io_counterMatrix1_bits_3_5 = _GEN_753[15:0];
  assign io_counterMatrix1_bits_3_6 = _GEN_754[15:0];
  assign io_counterMatrix1_bits_3_7 = _GEN_755[15:0];
  assign io_counterMatrix1_bits_4_0 = _GEN_756[15:0];
  assign io_counterMatrix1_bits_4_1 = _GEN_757[15:0];
  assign io_counterMatrix1_bits_4_2 = _GEN_758[15:0];
  assign io_counterMatrix1_bits_4_3 = _GEN_759[15:0];
  assign io_counterMatrix1_bits_4_4 = _GEN_760[15:0];
  assign io_counterMatrix1_bits_4_5 = _GEN_761[15:0];
  assign io_counterMatrix1_bits_4_6 = _GEN_762[15:0];
  assign io_counterMatrix1_bits_4_7 = _GEN_763[15:0];
  assign io_counterMatrix1_bits_5_0 = _GEN_764[15:0];
  assign io_counterMatrix1_bits_5_1 = _GEN_765[15:0];
  assign io_counterMatrix1_bits_5_2 = _GEN_766[15:0];
  assign io_counterMatrix1_bits_5_3 = _GEN_767[15:0];
  assign io_counterMatrix1_bits_5_4 = _GEN_768[15:0];
  assign io_counterMatrix1_bits_5_5 = _GEN_769[15:0];
  assign io_counterMatrix1_bits_5_6 = _GEN_770[15:0];
  assign io_counterMatrix1_bits_5_7 = _GEN_771[15:0];
  assign io_counterMatrix1_bits_6_0 = _GEN_772[15:0];
  assign io_counterMatrix1_bits_6_1 = _GEN_773[15:0];
  assign io_counterMatrix1_bits_6_2 = _GEN_774[15:0];
  assign io_counterMatrix1_bits_6_3 = _GEN_775[15:0];
  assign io_counterMatrix1_bits_6_4 = _GEN_776[15:0];
  assign io_counterMatrix1_bits_6_5 = _GEN_777[15:0];
  assign io_counterMatrix1_bits_6_6 = _GEN_778[15:0];
  assign io_counterMatrix1_bits_6_7 = _GEN_779[15:0];
  assign io_counterMatrix1_bits_7_0 = _GEN_780[15:0];
  assign io_counterMatrix1_bits_7_1 = _GEN_781[15:0];
  assign io_counterMatrix1_bits_7_2 = _GEN_782[15:0];
  assign io_counterMatrix1_bits_7_3 = _GEN_783[15:0];
  assign io_counterMatrix1_bits_7_4 = _GEN_784[15:0];
  assign io_counterMatrix1_bits_7_5 = _GEN_785[15:0];
  assign io_counterMatrix1_bits_7_6 = _GEN_786[15:0];
  assign io_counterMatrix1_bits_7_7 = _GEN_787[15:0];
  assign io_counterMatrix2_bits_0 = _GEN_788[15:0];
  assign io_counterMatrix2_bits_1 = _GEN_789[15:0];
  assign io_counterMatrix2_bits_2 = _GEN_790[15:0];
  assign io_counterMatrix2_bits_3 = _GEN_791[15:0];
  assign io_counterMatrix2_bits_4 = _GEN_792[15:0];
  assign io_counterMatrix2_bits_5 = _GEN_793[15:0];
  assign io_counterMatrix2_bits_6 = _GEN_794[15:0];
  assign io_counterMatrix2_bits_7 = _GEN_795[15:0];
  assign io_valid = io_start & (i == 32'h3 & j == 32'h3); // @[SourceDestination.scala 104:14 122:12 34:17]
  always @(posedge clock) begin
    prevStationary_matrix_0_0 <= io_Stationary_matrix_0_0; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_0_1 <= io_Stationary_matrix_0_1; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_0_2 <= io_Stationary_matrix_0_2; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_0_3 <= io_Stationary_matrix_0_3; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_0_4 <= io_Stationary_matrix_0_4; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_0_5 <= io_Stationary_matrix_0_5; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_0_6 <= io_Stationary_matrix_0_6; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_0_7 <= io_Stationary_matrix_0_7; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_1_0 <= io_Stationary_matrix_1_0; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_1_1 <= io_Stationary_matrix_1_1; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_1_2 <= io_Stationary_matrix_1_2; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_1_3 <= io_Stationary_matrix_1_3; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_1_4 <= io_Stationary_matrix_1_4; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_1_5 <= io_Stationary_matrix_1_5; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_1_6 <= io_Stationary_matrix_1_6; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_1_7 <= io_Stationary_matrix_1_7; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_2_0 <= io_Stationary_matrix_2_0; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_2_1 <= io_Stationary_matrix_2_1; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_2_2 <= io_Stationary_matrix_2_2; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_2_3 <= io_Stationary_matrix_2_3; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_2_4 <= io_Stationary_matrix_2_4; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_2_5 <= io_Stationary_matrix_2_5; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_2_6 <= io_Stationary_matrix_2_6; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_2_7 <= io_Stationary_matrix_2_7; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_3_0 <= io_Stationary_matrix_3_0; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_3_1 <= io_Stationary_matrix_3_1; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_3_2 <= io_Stationary_matrix_3_2; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_3_3 <= io_Stationary_matrix_3_3; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_3_4 <= io_Stationary_matrix_3_4; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_3_5 <= io_Stationary_matrix_3_5; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_3_6 <= io_Stationary_matrix_3_6; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_3_7 <= io_Stationary_matrix_3_7; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_4_0 <= io_Stationary_matrix_4_0; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_4_1 <= io_Stationary_matrix_4_1; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_4_2 <= io_Stationary_matrix_4_2; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_4_3 <= io_Stationary_matrix_4_3; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_4_4 <= io_Stationary_matrix_4_4; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_4_5 <= io_Stationary_matrix_4_5; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_4_6 <= io_Stationary_matrix_4_6; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_4_7 <= io_Stationary_matrix_4_7; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_5_0 <= io_Stationary_matrix_5_0; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_5_1 <= io_Stationary_matrix_5_1; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_5_2 <= io_Stationary_matrix_5_2; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_5_3 <= io_Stationary_matrix_5_3; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_5_4 <= io_Stationary_matrix_5_4; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_5_5 <= io_Stationary_matrix_5_5; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_5_6 <= io_Stationary_matrix_5_6; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_5_7 <= io_Stationary_matrix_5_7; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_6_0 <= io_Stationary_matrix_6_0; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_6_1 <= io_Stationary_matrix_6_1; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_6_2 <= io_Stationary_matrix_6_2; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_6_3 <= io_Stationary_matrix_6_3; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_6_4 <= io_Stationary_matrix_6_4; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_6_5 <= io_Stationary_matrix_6_5; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_6_6 <= io_Stationary_matrix_6_6; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_6_7 <= io_Stationary_matrix_6_7; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_7_0 <= io_Stationary_matrix_7_0; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_7_1 <= io_Stationary_matrix_7_1; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_7_2 <= io_Stationary_matrix_7_2; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_7_3 <= io_Stationary_matrix_7_3; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_7_4 <= io_Stationary_matrix_7_4; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_7_5 <= io_Stationary_matrix_7_5; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_7_6 <= io_Stationary_matrix_7_6; // @[SourceDestination.scala 15:40]
    prevStationary_matrix_7_7 <= io_Stationary_matrix_7_7; // @[SourceDestination.scala 15:40]
    if (io_start) begin // @[SourceDestination.scala 34:17]
      if (io_Stationary_matrix_7_7 != prevStationary_matrix_7_7) begin // @[SourceDestination.scala 40:74]
        matricesAreEqual <= 1'h0; // @[SourceDestination.scala 41:28]
      end else if (io_Stationary_matrix_7_6 != prevStationary_matrix_7_6) begin // @[SourceDestination.scala 40:74]
        matricesAreEqual <= 1'h0; // @[SourceDestination.scala 41:28]
      end else if (io_Stationary_matrix_7_5 != prevStationary_matrix_7_5) begin // @[SourceDestination.scala 40:74]
        matricesAreEqual <= 1'h0; // @[SourceDestination.scala 41:28]
      end else begin
        matricesAreEqual <= _GEN_60;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_0_0 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_0_0 <= _GEN_386;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_0_0 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_0_0 <= _GEN_386;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_0_1 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_0_1 <= _GEN_387;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_0_1 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_0_1 <= _GEN_387;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_0_2 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_0_2 <= _GEN_388;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_0_2 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_0_2 <= _GEN_388;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_0_3 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_0_3 <= _GEN_389;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_0_3 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_0_3 <= _GEN_389;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_0_4 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_0_4 <= _GEN_390;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_0_4 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_0_4 <= _GEN_390;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_0_5 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_0_5 <= _GEN_391;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_0_5 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_0_5 <= _GEN_391;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_0_6 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_0_6 <= _GEN_392;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_0_6 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_0_6 <= _GEN_392;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_0_7 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_0_7 <= _GEN_393;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_0_7 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_0_7 <= _GEN_393;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_1_0 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_1_0 <= _GEN_394;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_1_0 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_1_0 <= _GEN_394;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_1_1 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_1_1 <= _GEN_395;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_1_1 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_1_1 <= _GEN_395;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_1_2 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_1_2 <= _GEN_396;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_1_2 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_1_2 <= _GEN_396;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_1_3 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_1_3 <= _GEN_397;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_1_3 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_1_3 <= _GEN_397;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_1_4 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_1_4 <= _GEN_398;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_1_4 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_1_4 <= _GEN_398;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_1_5 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_1_5 <= _GEN_399;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_1_5 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_1_5 <= _GEN_399;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_1_6 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_1_6 <= _GEN_400;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_1_6 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_1_6 <= _GEN_400;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_1_7 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_1_7 <= _GEN_401;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_1_7 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_1_7 <= _GEN_401;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_2_0 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_2_0 <= _GEN_402;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_2_0 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_2_0 <= _GEN_402;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_2_1 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_2_1 <= _GEN_403;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_2_1 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_2_1 <= _GEN_403;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_2_2 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_2_2 <= _GEN_404;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_2_2 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_2_2 <= _GEN_404;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_2_3 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_2_3 <= _GEN_405;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_2_3 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_2_3 <= _GEN_405;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_2_4 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_2_4 <= _GEN_406;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_2_4 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_2_4 <= _GEN_406;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_2_5 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_2_5 <= _GEN_407;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_2_5 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_2_5 <= _GEN_407;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_2_6 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_2_6 <= _GEN_408;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_2_6 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_2_6 <= _GEN_408;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_2_7 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_2_7 <= _GEN_409;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_2_7 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_2_7 <= _GEN_409;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_3_0 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_3_0 <= _GEN_410;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_3_0 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_3_0 <= _GEN_410;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_3_1 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_3_1 <= _GEN_411;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_3_1 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_3_1 <= _GEN_411;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_3_2 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_3_2 <= _GEN_412;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_3_2 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_3_2 <= _GEN_412;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_3_3 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_3_3 <= _GEN_413;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_3_3 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_3_3 <= _GEN_413;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_3_4 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_3_4 <= _GEN_414;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_3_4 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_3_4 <= _GEN_414;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_3_5 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_3_5 <= _GEN_415;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_3_5 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_3_5 <= _GEN_415;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_3_6 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_3_6 <= _GEN_416;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_3_6 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_3_6 <= _GEN_416;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_3_7 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_3_7 <= _GEN_417;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_3_7 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_3_7 <= _GEN_417;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_4_0 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_4_0 <= _GEN_418;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_4_0 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_4_0 <= _GEN_418;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_4_1 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_4_1 <= _GEN_419;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_4_1 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_4_1 <= _GEN_419;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_4_2 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_4_2 <= _GEN_420;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_4_2 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_4_2 <= _GEN_420;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_4_3 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_4_3 <= _GEN_421;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_4_3 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_4_3 <= _GEN_421;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_4_4 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_4_4 <= _GEN_422;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_4_4 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_4_4 <= _GEN_422;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_4_5 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_4_5 <= _GEN_423;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_4_5 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_4_5 <= _GEN_423;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_4_6 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_4_6 <= _GEN_424;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_4_6 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_4_6 <= _GEN_424;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_4_7 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_4_7 <= _GEN_425;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_4_7 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_4_7 <= _GEN_425;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_5_0 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_5_0 <= _GEN_426;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_5_0 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_5_0 <= _GEN_426;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_5_1 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_5_1 <= _GEN_427;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_5_1 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_5_1 <= _GEN_427;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_5_2 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_5_2 <= _GEN_428;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_5_2 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_5_2 <= _GEN_428;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_5_3 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_5_3 <= _GEN_429;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_5_3 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_5_3 <= _GEN_429;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_5_4 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_5_4 <= _GEN_430;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_5_4 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_5_4 <= _GEN_430;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_5_5 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_5_5 <= _GEN_431;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_5_5 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_5_5 <= _GEN_431;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_5_6 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_5_6 <= _GEN_432;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_5_6 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_5_6 <= _GEN_432;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_5_7 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_5_7 <= _GEN_433;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_5_7 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_5_7 <= _GEN_433;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_6_0 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_6_0 <= _GEN_434;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_6_0 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_6_0 <= _GEN_434;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_6_1 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_6_1 <= _GEN_435;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_6_1 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_6_1 <= _GEN_435;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_6_2 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_6_2 <= _GEN_436;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_6_2 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_6_2 <= _GEN_436;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_6_3 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_6_3 <= _GEN_437;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_6_3 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_6_3 <= _GEN_437;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_6_4 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_6_4 <= _GEN_438;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_6_4 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_6_4 <= _GEN_438;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_6_5 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_6_5 <= _GEN_439;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_6_5 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_6_5 <= _GEN_439;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_6_6 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_6_6 <= _GEN_440;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_6_6 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_6_6 <= _GEN_440;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_6_7 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_6_7 <= _GEN_441;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_6_7 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_6_7 <= _GEN_441;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_7_0 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_7_0 <= _GEN_442;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_7_0 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_7_0 <= _GEN_442;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_7_1 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_7_1 <= _GEN_443;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_7_1 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_7_1 <= _GEN_443;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_7_2 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_7_2 <= _GEN_444;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_7_2 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_7_2 <= _GEN_444;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_7_3 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_7_3 <= _GEN_445;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_7_3 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_7_3 <= _GEN_445;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_7_4 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_7_4 <= _GEN_446;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_7_4 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_7_4 <= _GEN_446;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_7_5 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_7_5 <= _GEN_447;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_7_5 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_7_5 <= _GEN_447;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_7_6 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_7_6 <= _GEN_448;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_7_6 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_7_6 <= _GEN_448;
      end
    end
    if (reset) begin // @[SourceDestination.scala 17:31]
      counterRegs1_7_7 <= 16'h0; // @[SourceDestination.scala 17:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs1_7_7 <= _GEN_449;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs1_7_7 <= 16'h0; // @[SourceDestination.scala 98:30]
      end else begin
        counterRegs1_7_7 <= _GEN_449;
      end
    end
    if (reset) begin // @[SourceDestination.scala 18:31]
      counterRegs2_0 <= 16'h0; // @[SourceDestination.scala 18:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs2_0 <= _GEN_467;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs2_0 <= 16'h0; // @[SourceDestination.scala 100:25]
      end else begin
        counterRegs2_0 <= _GEN_467;
      end
    end
    if (reset) begin // @[SourceDestination.scala 18:31]
      counterRegs2_1 <= 16'h0; // @[SourceDestination.scala 18:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs2_1 <= _GEN_468;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs2_1 <= 16'h0; // @[SourceDestination.scala 100:25]
      end else begin
        counterRegs2_1 <= _GEN_468;
      end
    end
    if (reset) begin // @[SourceDestination.scala 18:31]
      counterRegs2_2 <= 16'h0; // @[SourceDestination.scala 18:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs2_2 <= _GEN_469;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs2_2 <= 16'h0; // @[SourceDestination.scala 100:25]
      end else begin
        counterRegs2_2 <= _GEN_469;
      end
    end
    if (reset) begin // @[SourceDestination.scala 18:31]
      counterRegs2_3 <= 16'h0; // @[SourceDestination.scala 18:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs2_3 <= _GEN_470;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs2_3 <= 16'h0; // @[SourceDestination.scala 100:25]
      end else begin
        counterRegs2_3 <= _GEN_470;
      end
    end
    if (reset) begin // @[SourceDestination.scala 18:31]
      counterRegs2_4 <= 16'h0; // @[SourceDestination.scala 18:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs2_4 <= _GEN_471;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs2_4 <= 16'h0; // @[SourceDestination.scala 100:25]
      end else begin
        counterRegs2_4 <= _GEN_471;
      end
    end
    if (reset) begin // @[SourceDestination.scala 18:31]
      counterRegs2_5 <= 16'h0; // @[SourceDestination.scala 18:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs2_5 <= _GEN_472;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs2_5 <= 16'h0; // @[SourceDestination.scala 100:25]
      end else begin
        counterRegs2_5 <= _GEN_472;
      end
    end
    if (reset) begin // @[SourceDestination.scala 18:31]
      counterRegs2_6 <= 16'h0; // @[SourceDestination.scala 18:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs2_6 <= _GEN_473;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs2_6 <= 16'h0; // @[SourceDestination.scala 100:25]
      end else begin
        counterRegs2_6 <= _GEN_473;
      end
    end
    if (reset) begin // @[SourceDestination.scala 18:31]
      counterRegs2_7 <= 16'h0; // @[SourceDestination.scala 18:31]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counterRegs2_7 <= _GEN_474;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counterRegs2_7 <= 16'h0; // @[SourceDestination.scala 100:25]
      end else begin
        counterRegs2_7 <= _GEN_474;
      end
    end
    if (reset) begin // @[SourceDestination.scala 20:20]
      i <= 32'h0; // @[SourceDestination.scala 20:20]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        if (!(j < 32'h7)) begin // @[SourceDestination.scala 80:40]
          i <= _GEN_482;
        end
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        i <= 32'h0; // @[SourceDestination.scala 91:9]
      end
    end
    if (reset) begin // @[SourceDestination.scala 21:20]
      j <= 32'h0; // @[SourceDestination.scala 21:20]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        if (j < 32'h7) begin // @[SourceDestination.scala 80:40]
          j <= _j_T_1; // @[SourceDestination.scala 81:11]
        end else begin
          j <= _GEN_481;
        end
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        j <= 32'h0; // @[SourceDestination.scala 92:9]
      end
    end
    if (io_start) begin // @[SourceDestination.scala 34:17]
      jValid <= _GEN_564;
    end
    if (reset) begin // @[SourceDestination.scala 26:20]
      k <= 32'h0; // @[SourceDestination.scala 26:20]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        k <= _GEN_477;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        k <= 32'h0; // @[SourceDestination.scala 93:9]
      end else begin
        k <= _GEN_477;
      end
    end
    if (reset) begin // @[SourceDestination.scala 28:27]
      counter1 <= 32'h1; // @[SourceDestination.scala 28:27]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counter1 <= _GEN_450;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counter1 <= 32'h1; // @[SourceDestination.scala 94:16]
      end else begin
        counter1 <= _GEN_450;
      end
    end
    if (reset) begin // @[SourceDestination.scala 29:27]
      counter2 <= 32'h1; // @[SourceDestination.scala 29:27]
    end else if (io_start) begin // @[SourceDestination.scala 34:17]
      if (~jValid) begin // @[SourceDestination.scala 79:26]
        counter2 <= _GEN_478;
      end else if (jValid & ~matricesAreEqual) begin // @[SourceDestination.scala 90:64]
        counter2 <= 32'h1; // @[SourceDestination.scala 95:16]
      end else begin
        counter2 <= _GEN_478;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  prevStationary_matrix_0_0 = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  prevStationary_matrix_0_1 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  prevStationary_matrix_0_2 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  prevStationary_matrix_0_3 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  prevStationary_matrix_0_4 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  prevStationary_matrix_0_5 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  prevStationary_matrix_0_6 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  prevStationary_matrix_0_7 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  prevStationary_matrix_1_0 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  prevStationary_matrix_1_1 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  prevStationary_matrix_1_2 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  prevStationary_matrix_1_3 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  prevStationary_matrix_1_4 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  prevStationary_matrix_1_5 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  prevStationary_matrix_1_6 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  prevStationary_matrix_1_7 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  prevStationary_matrix_2_0 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  prevStationary_matrix_2_1 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  prevStationary_matrix_2_2 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  prevStationary_matrix_2_3 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  prevStationary_matrix_2_4 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  prevStationary_matrix_2_5 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  prevStationary_matrix_2_6 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  prevStationary_matrix_2_7 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  prevStationary_matrix_3_0 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  prevStationary_matrix_3_1 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  prevStationary_matrix_3_2 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  prevStationary_matrix_3_3 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  prevStationary_matrix_3_4 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  prevStationary_matrix_3_5 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  prevStationary_matrix_3_6 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  prevStationary_matrix_3_7 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  prevStationary_matrix_4_0 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  prevStationary_matrix_4_1 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  prevStationary_matrix_4_2 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  prevStationary_matrix_4_3 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  prevStationary_matrix_4_4 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  prevStationary_matrix_4_5 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  prevStationary_matrix_4_6 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  prevStationary_matrix_4_7 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  prevStationary_matrix_5_0 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  prevStationary_matrix_5_1 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  prevStationary_matrix_5_2 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  prevStationary_matrix_5_3 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  prevStationary_matrix_5_4 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  prevStationary_matrix_5_5 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  prevStationary_matrix_5_6 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  prevStationary_matrix_5_7 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  prevStationary_matrix_6_0 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  prevStationary_matrix_6_1 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  prevStationary_matrix_6_2 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  prevStationary_matrix_6_3 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  prevStationary_matrix_6_4 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  prevStationary_matrix_6_5 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  prevStationary_matrix_6_6 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  prevStationary_matrix_6_7 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  prevStationary_matrix_7_0 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  prevStationary_matrix_7_1 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  prevStationary_matrix_7_2 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  prevStationary_matrix_7_3 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  prevStationary_matrix_7_4 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  prevStationary_matrix_7_5 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  prevStationary_matrix_7_6 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  prevStationary_matrix_7_7 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  matricesAreEqual = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  counterRegs1_0_0 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  counterRegs1_0_1 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  counterRegs1_0_2 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  counterRegs1_0_3 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  counterRegs1_0_4 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  counterRegs1_0_5 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  counterRegs1_0_6 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  counterRegs1_0_7 = _RAND_72[15:0];
  _RAND_73 = {1{`RANDOM}};
  counterRegs1_1_0 = _RAND_73[15:0];
  _RAND_74 = {1{`RANDOM}};
  counterRegs1_1_1 = _RAND_74[15:0];
  _RAND_75 = {1{`RANDOM}};
  counterRegs1_1_2 = _RAND_75[15:0];
  _RAND_76 = {1{`RANDOM}};
  counterRegs1_1_3 = _RAND_76[15:0];
  _RAND_77 = {1{`RANDOM}};
  counterRegs1_1_4 = _RAND_77[15:0];
  _RAND_78 = {1{`RANDOM}};
  counterRegs1_1_5 = _RAND_78[15:0];
  _RAND_79 = {1{`RANDOM}};
  counterRegs1_1_6 = _RAND_79[15:0];
  _RAND_80 = {1{`RANDOM}};
  counterRegs1_1_7 = _RAND_80[15:0];
  _RAND_81 = {1{`RANDOM}};
  counterRegs1_2_0 = _RAND_81[15:0];
  _RAND_82 = {1{`RANDOM}};
  counterRegs1_2_1 = _RAND_82[15:0];
  _RAND_83 = {1{`RANDOM}};
  counterRegs1_2_2 = _RAND_83[15:0];
  _RAND_84 = {1{`RANDOM}};
  counterRegs1_2_3 = _RAND_84[15:0];
  _RAND_85 = {1{`RANDOM}};
  counterRegs1_2_4 = _RAND_85[15:0];
  _RAND_86 = {1{`RANDOM}};
  counterRegs1_2_5 = _RAND_86[15:0];
  _RAND_87 = {1{`RANDOM}};
  counterRegs1_2_6 = _RAND_87[15:0];
  _RAND_88 = {1{`RANDOM}};
  counterRegs1_2_7 = _RAND_88[15:0];
  _RAND_89 = {1{`RANDOM}};
  counterRegs1_3_0 = _RAND_89[15:0];
  _RAND_90 = {1{`RANDOM}};
  counterRegs1_3_1 = _RAND_90[15:0];
  _RAND_91 = {1{`RANDOM}};
  counterRegs1_3_2 = _RAND_91[15:0];
  _RAND_92 = {1{`RANDOM}};
  counterRegs1_3_3 = _RAND_92[15:0];
  _RAND_93 = {1{`RANDOM}};
  counterRegs1_3_4 = _RAND_93[15:0];
  _RAND_94 = {1{`RANDOM}};
  counterRegs1_3_5 = _RAND_94[15:0];
  _RAND_95 = {1{`RANDOM}};
  counterRegs1_3_6 = _RAND_95[15:0];
  _RAND_96 = {1{`RANDOM}};
  counterRegs1_3_7 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  counterRegs1_4_0 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  counterRegs1_4_1 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  counterRegs1_4_2 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  counterRegs1_4_3 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  counterRegs1_4_4 = _RAND_101[15:0];
  _RAND_102 = {1{`RANDOM}};
  counterRegs1_4_5 = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  counterRegs1_4_6 = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  counterRegs1_4_7 = _RAND_104[15:0];
  _RAND_105 = {1{`RANDOM}};
  counterRegs1_5_0 = _RAND_105[15:0];
  _RAND_106 = {1{`RANDOM}};
  counterRegs1_5_1 = _RAND_106[15:0];
  _RAND_107 = {1{`RANDOM}};
  counterRegs1_5_2 = _RAND_107[15:0];
  _RAND_108 = {1{`RANDOM}};
  counterRegs1_5_3 = _RAND_108[15:0];
  _RAND_109 = {1{`RANDOM}};
  counterRegs1_5_4 = _RAND_109[15:0];
  _RAND_110 = {1{`RANDOM}};
  counterRegs1_5_5 = _RAND_110[15:0];
  _RAND_111 = {1{`RANDOM}};
  counterRegs1_5_6 = _RAND_111[15:0];
  _RAND_112 = {1{`RANDOM}};
  counterRegs1_5_7 = _RAND_112[15:0];
  _RAND_113 = {1{`RANDOM}};
  counterRegs1_6_0 = _RAND_113[15:0];
  _RAND_114 = {1{`RANDOM}};
  counterRegs1_6_1 = _RAND_114[15:0];
  _RAND_115 = {1{`RANDOM}};
  counterRegs1_6_2 = _RAND_115[15:0];
  _RAND_116 = {1{`RANDOM}};
  counterRegs1_6_3 = _RAND_116[15:0];
  _RAND_117 = {1{`RANDOM}};
  counterRegs1_6_4 = _RAND_117[15:0];
  _RAND_118 = {1{`RANDOM}};
  counterRegs1_6_5 = _RAND_118[15:0];
  _RAND_119 = {1{`RANDOM}};
  counterRegs1_6_6 = _RAND_119[15:0];
  _RAND_120 = {1{`RANDOM}};
  counterRegs1_6_7 = _RAND_120[15:0];
  _RAND_121 = {1{`RANDOM}};
  counterRegs1_7_0 = _RAND_121[15:0];
  _RAND_122 = {1{`RANDOM}};
  counterRegs1_7_1 = _RAND_122[15:0];
  _RAND_123 = {1{`RANDOM}};
  counterRegs1_7_2 = _RAND_123[15:0];
  _RAND_124 = {1{`RANDOM}};
  counterRegs1_7_3 = _RAND_124[15:0];
  _RAND_125 = {1{`RANDOM}};
  counterRegs1_7_4 = _RAND_125[15:0];
  _RAND_126 = {1{`RANDOM}};
  counterRegs1_7_5 = _RAND_126[15:0];
  _RAND_127 = {1{`RANDOM}};
  counterRegs1_7_6 = _RAND_127[15:0];
  _RAND_128 = {1{`RANDOM}};
  counterRegs1_7_7 = _RAND_128[15:0];
  _RAND_129 = {1{`RANDOM}};
  counterRegs2_0 = _RAND_129[15:0];
  _RAND_130 = {1{`RANDOM}};
  counterRegs2_1 = _RAND_130[15:0];
  _RAND_131 = {1{`RANDOM}};
  counterRegs2_2 = _RAND_131[15:0];
  _RAND_132 = {1{`RANDOM}};
  counterRegs2_3 = _RAND_132[15:0];
  _RAND_133 = {1{`RANDOM}};
  counterRegs2_4 = _RAND_133[15:0];
  _RAND_134 = {1{`RANDOM}};
  counterRegs2_5 = _RAND_134[15:0];
  _RAND_135 = {1{`RANDOM}};
  counterRegs2_6 = _RAND_135[15:0];
  _RAND_136 = {1{`RANDOM}};
  counterRegs2_7 = _RAND_136[15:0];
  _RAND_137 = {1{`RANDOM}};
  i = _RAND_137[31:0];
  _RAND_138 = {1{`RANDOM}};
  j = _RAND_138[31:0];
  _RAND_139 = {1{`RANDOM}};
  jValid = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  k = _RAND_140[31:0];
  _RAND_141 = {1{`RANDOM}};
  counter1 = _RAND_141[31:0];
  _RAND_142 = {1{`RANDOM}};
  counter2 = _RAND_142[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SingleLoop2(
  input         clock,
  input         reset,
  input  [31:0] io_IDex,
  input  [31:0] io_JDex,
  input         io_valid,
  input  [31:0] io_mat_0_0,
  input  [31:0] io_mat_0_1,
  input  [31:0] io_mat_0_2,
  input  [31:0] io_mat_0_3,
  input  [31:0] io_mat_0_4,
  input  [31:0] io_mat_0_5,
  input  [31:0] io_mat_0_6,
  input  [31:0] io_mat_0_7,
  input  [31:0] io_mat_1_0,
  input  [31:0] io_mat_1_1,
  input  [31:0] io_mat_1_2,
  input  [31:0] io_mat_1_3,
  input  [31:0] io_mat_1_4,
  input  [31:0] io_mat_1_5,
  input  [31:0] io_mat_1_6,
  input  [31:0] io_mat_1_7,
  input  [31:0] io_mat_2_0,
  input  [31:0] io_mat_2_1,
  input  [31:0] io_mat_2_2,
  input  [31:0] io_mat_2_3,
  input  [31:0] io_mat_2_4,
  input  [31:0] io_mat_2_5,
  input  [31:0] io_mat_2_6,
  input  [31:0] io_mat_2_7,
  input  [31:0] io_mat_3_0,
  input  [31:0] io_mat_3_1,
  input  [31:0] io_mat_3_2,
  input  [31:0] io_mat_3_3,
  input  [31:0] io_mat_3_4,
  input  [31:0] io_mat_3_5,
  input  [31:0] io_mat_3_6,
  input  [31:0] io_mat_3_7,
  input  [31:0] io_mat_4_0,
  input  [31:0] io_mat_4_1,
  input  [31:0] io_mat_4_2,
  input  [31:0] io_mat_4_3,
  input  [31:0] io_mat_4_4,
  input  [31:0] io_mat_4_5,
  input  [31:0] io_mat_4_6,
  input  [31:0] io_mat_4_7,
  input  [31:0] io_mat_5_0,
  input  [31:0] io_mat_5_1,
  input  [31:0] io_mat_5_2,
  input  [31:0] io_mat_5_3,
  input  [31:0] io_mat_5_4,
  input  [31:0] io_mat_5_5,
  input  [31:0] io_mat_5_6,
  input  [31:0] io_mat_5_7,
  input  [31:0] io_mat_6_0,
  input  [31:0] io_mat_6_1,
  input  [31:0] io_mat_6_2,
  input  [31:0] io_mat_6_3,
  input  [31:0] io_mat_6_4,
  input  [31:0] io_mat_6_5,
  input  [31:0] io_mat_6_6,
  input  [31:0] io_mat_6_7,
  input  [31:0] io_mat_7_0,
  input  [31:0] io_mat_7_1,
  input  [31:0] io_mat_7_2,
  input  [31:0] io_mat_7_3,
  input  [31:0] io_mat_7_4,
  input  [31:0] io_mat_7_5,
  input  [31:0] io_mat_7_6,
  input  [31:0] io_mat_7_7,
  output [31:0] io_OutMat_0_0,
  output [31:0] io_OutMat_0_1,
  output [31:0] io_OutMat_0_2,
  output [31:0] io_OutMat_0_3,
  output [31:0] io_OutMat_0_4,
  output [31:0] io_OutMat_0_5,
  output [31:0] io_OutMat_0_6,
  output [31:0] io_OutMat_0_7,
  output [31:0] io_OutMat_1_0,
  output [31:0] io_OutMat_1_1,
  output [31:0] io_OutMat_1_2,
  output [31:0] io_OutMat_1_3,
  output [31:0] io_OutMat_1_4,
  output [31:0] io_OutMat_1_5,
  output [31:0] io_OutMat_1_6,
  output [31:0] io_OutMat_1_7,
  output [31:0] io_OutMat_2_0,
  output [31:0] io_OutMat_2_1,
  output [31:0] io_OutMat_2_2,
  output [31:0] io_OutMat_2_3,
  output [31:0] io_OutMat_2_4,
  output [31:0] io_OutMat_2_5,
  output [31:0] io_OutMat_2_6,
  output [31:0] io_OutMat_2_7,
  output [31:0] io_OutMat_3_0,
  output [31:0] io_OutMat_3_1,
  output [31:0] io_OutMat_3_2,
  output [31:0] io_OutMat_3_3,
  output [31:0] io_OutMat_3_4,
  output [31:0] io_OutMat_3_5,
  output [31:0] io_OutMat_3_6,
  output [31:0] io_OutMat_3_7,
  output [31:0] io_OutMat_4_0,
  output [31:0] io_OutMat_4_1,
  output [31:0] io_OutMat_4_2,
  output [31:0] io_OutMat_4_3,
  output [31:0] io_OutMat_4_4,
  output [31:0] io_OutMat_4_5,
  output [31:0] io_OutMat_4_6,
  output [31:0] io_OutMat_4_7,
  output [31:0] io_OutMat_5_0,
  output [31:0] io_OutMat_5_1,
  output [31:0] io_OutMat_5_2,
  output [31:0] io_OutMat_5_3,
  output [31:0] io_OutMat_5_4,
  output [31:0] io_OutMat_5_5,
  output [31:0] io_OutMat_5_6,
  output [31:0] io_OutMat_5_7,
  output [31:0] io_OutMat_6_0,
  output [31:0] io_OutMat_6_1,
  output [31:0] io_OutMat_6_2,
  output [31:0] io_OutMat_6_3,
  output [31:0] io_OutMat_6_4,
  output [31:0] io_OutMat_6_5,
  output [31:0] io_OutMat_6_6,
  output [31:0] io_OutMat_6_7,
  output [31:0] io_OutMat_7_0,
  output [31:0] io_OutMat_7_1,
  output [31:0] io_OutMat_7_2,
  output [31:0] io_OutMat_7_3,
  output [31:0] io_OutMat_7_4,
  output [31:0] io_OutMat_7_5,
  output [31:0] io_OutMat_7_6,
  output [31:0] io_OutMat_7_7,
  output        io_Ovalid,
  output        io_ProcessValid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] b_0_0; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_0_1; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_0_2; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_0_3; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_0_4; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_0_5; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_0_6; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_0_7; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_1_0; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_1_1; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_1_2; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_1_3; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_1_4; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_1_5; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_1_6; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_1_7; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_2_0; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_2_1; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_2_2; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_2_3; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_2_4; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_2_5; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_2_6; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_2_7; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_3_0; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_3_1; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_3_2; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_3_3; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_3_4; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_3_5; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_3_6; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_3_7; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_4_0; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_4_1; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_4_2; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_4_3; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_4_4; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_4_5; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_4_6; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_4_7; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_5_0; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_5_1; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_5_2; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_5_3; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_5_4; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_5_5; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_5_6; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_5_7; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_6_0; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_6_1; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_6_2; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_6_3; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_6_4; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_6_5; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_6_6; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_6_7; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_7_0; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_7_1; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_7_2; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_7_3; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_7_4; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_7_5; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_7_6; // @[SingleLoop2.scala 17:20]
  reg [31:0] b_7_7; // @[SingleLoop2.scala 17:20]
  reg [31:0] j; // @[SingleLoop2.scala 19:16]
  wire [31:0] _GEN_65 = 3'h0 == io_IDex[2:0] & 3'h1 == j[2:0] ? io_mat_0_1 : io_mat_0_0; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_66 = 3'h0 == io_IDex[2:0] & 3'h2 == j[2:0] ? io_mat_0_2 : _GEN_65; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_67 = 3'h0 == io_IDex[2:0] & 3'h3 == j[2:0] ? io_mat_0_3 : _GEN_66; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_68 = 3'h0 == io_IDex[2:0] & 3'h4 == j[2:0] ? io_mat_0_4 : _GEN_67; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_69 = 3'h0 == io_IDex[2:0] & 3'h5 == j[2:0] ? io_mat_0_5 : _GEN_68; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_70 = 3'h0 == io_IDex[2:0] & 3'h6 == j[2:0] ? io_mat_0_6 : _GEN_69; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_71 = 3'h0 == io_IDex[2:0] & 3'h7 == j[2:0] ? io_mat_0_7 : _GEN_70; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_72 = 3'h1 == io_IDex[2:0] & 3'h0 == j[2:0] ? io_mat_1_0 : _GEN_71; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_73 = 3'h1 == io_IDex[2:0] & 3'h1 == j[2:0] ? io_mat_1_1 : _GEN_72; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_74 = 3'h1 == io_IDex[2:0] & 3'h2 == j[2:0] ? io_mat_1_2 : _GEN_73; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_75 = 3'h1 == io_IDex[2:0] & 3'h3 == j[2:0] ? io_mat_1_3 : _GEN_74; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_76 = 3'h1 == io_IDex[2:0] & 3'h4 == j[2:0] ? io_mat_1_4 : _GEN_75; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_77 = 3'h1 == io_IDex[2:0] & 3'h5 == j[2:0] ? io_mat_1_5 : _GEN_76; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_78 = 3'h1 == io_IDex[2:0] & 3'h6 == j[2:0] ? io_mat_1_6 : _GEN_77; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_79 = 3'h1 == io_IDex[2:0] & 3'h7 == j[2:0] ? io_mat_1_7 : _GEN_78; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_80 = 3'h2 == io_IDex[2:0] & 3'h0 == j[2:0] ? io_mat_2_0 : _GEN_79; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_81 = 3'h2 == io_IDex[2:0] & 3'h1 == j[2:0] ? io_mat_2_1 : _GEN_80; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_82 = 3'h2 == io_IDex[2:0] & 3'h2 == j[2:0] ? io_mat_2_2 : _GEN_81; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_83 = 3'h2 == io_IDex[2:0] & 3'h3 == j[2:0] ? io_mat_2_3 : _GEN_82; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_84 = 3'h2 == io_IDex[2:0] & 3'h4 == j[2:0] ? io_mat_2_4 : _GEN_83; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_85 = 3'h2 == io_IDex[2:0] & 3'h5 == j[2:0] ? io_mat_2_5 : _GEN_84; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_86 = 3'h2 == io_IDex[2:0] & 3'h6 == j[2:0] ? io_mat_2_6 : _GEN_85; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_87 = 3'h2 == io_IDex[2:0] & 3'h7 == j[2:0] ? io_mat_2_7 : _GEN_86; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_88 = 3'h3 == io_IDex[2:0] & 3'h0 == j[2:0] ? io_mat_3_0 : _GEN_87; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_89 = 3'h3 == io_IDex[2:0] & 3'h1 == j[2:0] ? io_mat_3_1 : _GEN_88; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_90 = 3'h3 == io_IDex[2:0] & 3'h2 == j[2:0] ? io_mat_3_2 : _GEN_89; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_91 = 3'h3 == io_IDex[2:0] & 3'h3 == j[2:0] ? io_mat_3_3 : _GEN_90; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_92 = 3'h3 == io_IDex[2:0] & 3'h4 == j[2:0] ? io_mat_3_4 : _GEN_91; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_93 = 3'h3 == io_IDex[2:0] & 3'h5 == j[2:0] ? io_mat_3_5 : _GEN_92; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_94 = 3'h3 == io_IDex[2:0] & 3'h6 == j[2:0] ? io_mat_3_6 : _GEN_93; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_95 = 3'h3 == io_IDex[2:0] & 3'h7 == j[2:0] ? io_mat_3_7 : _GEN_94; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_96 = 3'h4 == io_IDex[2:0] & 3'h0 == j[2:0] ? io_mat_4_0 : _GEN_95; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_97 = 3'h4 == io_IDex[2:0] & 3'h1 == j[2:0] ? io_mat_4_1 : _GEN_96; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_98 = 3'h4 == io_IDex[2:0] & 3'h2 == j[2:0] ? io_mat_4_2 : _GEN_97; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_99 = 3'h4 == io_IDex[2:0] & 3'h3 == j[2:0] ? io_mat_4_3 : _GEN_98; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_100 = 3'h4 == io_IDex[2:0] & 3'h4 == j[2:0] ? io_mat_4_4 : _GEN_99; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_101 = 3'h4 == io_IDex[2:0] & 3'h5 == j[2:0] ? io_mat_4_5 : _GEN_100; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_102 = 3'h4 == io_IDex[2:0] & 3'h6 == j[2:0] ? io_mat_4_6 : _GEN_101; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_103 = 3'h4 == io_IDex[2:0] & 3'h7 == j[2:0] ? io_mat_4_7 : _GEN_102; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_104 = 3'h5 == io_IDex[2:0] & 3'h0 == j[2:0] ? io_mat_5_0 : _GEN_103; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_105 = 3'h5 == io_IDex[2:0] & 3'h1 == j[2:0] ? io_mat_5_1 : _GEN_104; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_106 = 3'h5 == io_IDex[2:0] & 3'h2 == j[2:0] ? io_mat_5_2 : _GEN_105; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_107 = 3'h5 == io_IDex[2:0] & 3'h3 == j[2:0] ? io_mat_5_3 : _GEN_106; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_108 = 3'h5 == io_IDex[2:0] & 3'h4 == j[2:0] ? io_mat_5_4 : _GEN_107; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_109 = 3'h5 == io_IDex[2:0] & 3'h5 == j[2:0] ? io_mat_5_5 : _GEN_108; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_110 = 3'h5 == io_IDex[2:0] & 3'h6 == j[2:0] ? io_mat_5_6 : _GEN_109; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_111 = 3'h5 == io_IDex[2:0] & 3'h7 == j[2:0] ? io_mat_5_7 : _GEN_110; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_112 = 3'h6 == io_IDex[2:0] & 3'h0 == j[2:0] ? io_mat_6_0 : _GEN_111; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_113 = 3'h6 == io_IDex[2:0] & 3'h1 == j[2:0] ? io_mat_6_1 : _GEN_112; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_114 = 3'h6 == io_IDex[2:0] & 3'h2 == j[2:0] ? io_mat_6_2 : _GEN_113; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_115 = 3'h6 == io_IDex[2:0] & 3'h3 == j[2:0] ? io_mat_6_3 : _GEN_114; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_116 = 3'h6 == io_IDex[2:0] & 3'h4 == j[2:0] ? io_mat_6_4 : _GEN_115; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_117 = 3'h6 == io_IDex[2:0] & 3'h5 == j[2:0] ? io_mat_6_5 : _GEN_116; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_118 = 3'h6 == io_IDex[2:0] & 3'h6 == j[2:0] ? io_mat_6_6 : _GEN_117; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_119 = 3'h6 == io_IDex[2:0] & 3'h7 == j[2:0] ? io_mat_6_7 : _GEN_118; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_120 = 3'h7 == io_IDex[2:0] & 3'h0 == j[2:0] ? io_mat_7_0 : _GEN_119; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_121 = 3'h7 == io_IDex[2:0] & 3'h1 == j[2:0] ? io_mat_7_1 : _GEN_120; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_122 = 3'h7 == io_IDex[2:0] & 3'h2 == j[2:0] ? io_mat_7_2 : _GEN_121; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_123 = 3'h7 == io_IDex[2:0] & 3'h3 == j[2:0] ? io_mat_7_3 : _GEN_122; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_124 = 3'h7 == io_IDex[2:0] & 3'h4 == j[2:0] ? io_mat_7_4 : _GEN_123; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_125 = 3'h7 == io_IDex[2:0] & 3'h5 == j[2:0] ? io_mat_7_5 : _GEN_124; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_126 = 3'h7 == io_IDex[2:0] & 3'h6 == j[2:0] ? io_mat_7_6 : _GEN_125; // @[SingleLoop2.scala 23:{19,19}]
  wire [31:0] _GEN_127 = 3'h7 == io_IDex[2:0] & 3'h7 == j[2:0] ? io_mat_7_7 : _GEN_126; // @[SingleLoop2.scala 23:{19,19}]
  wire  _T_4 = _GEN_127 == 32'h4; // @[SingleLoop2.scala 26:30]
  wire  _T_5 = j == 32'h7; // @[SingleLoop2.scala 30:18]
  wire  _T_9 = j == 32'h7 & _T_4; // @[SingleLoop2.scala 30:43]
  wire [31:0] _j_T_1 = j + 32'h1; // @[SingleLoop2.scala 40:16]
  assign io_OutMat_0_0 = b_0_0; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_0_1 = b_0_1; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_0_2 = b_0_2; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_0_3 = b_0_3; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_0_4 = b_0_4; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_0_5 = b_0_5; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_0_6 = b_0_6; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_0_7 = b_0_7; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_1_0 = b_1_0; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_1_1 = b_1_1; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_1_2 = b_1_2; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_1_3 = b_1_3; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_1_4 = b_1_4; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_1_5 = b_1_5; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_1_6 = b_1_6; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_1_7 = b_1_7; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_2_0 = b_2_0; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_2_1 = b_2_1; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_2_2 = b_2_2; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_2_3 = b_2_3; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_2_4 = b_2_4; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_2_5 = b_2_5; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_2_6 = b_2_6; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_2_7 = b_2_7; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_3_0 = b_3_0; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_3_1 = b_3_1; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_3_2 = b_3_2; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_3_3 = b_3_3; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_3_4 = b_3_4; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_3_5 = b_3_5; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_3_6 = b_3_6; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_3_7 = b_3_7; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_4_0 = b_4_0; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_4_1 = b_4_1; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_4_2 = b_4_2; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_4_3 = b_4_3; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_4_4 = b_4_4; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_4_5 = b_4_5; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_4_6 = b_4_6; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_4_7 = b_4_7; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_5_0 = b_5_0; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_5_1 = b_5_1; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_5_2 = b_5_2; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_5_3 = b_5_3; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_5_4 = b_5_4; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_5_5 = b_5_5; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_5_6 = b_5_6; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_5_7 = b_5_7; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_6_0 = b_6_0; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_6_1 = b_6_1; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_6_2 = b_6_2; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_6_3 = b_6_3; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_6_4 = b_6_4; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_6_5 = b_6_5; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_6_6 = b_6_6; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_6_7 = b_6_7; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_7_0 = b_7_0; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_7_1 = b_7_1; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_7_2 = b_7_2; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_7_3 = b_7_3; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_7_4 = b_7_4; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_7_5 = b_7_5; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_7_6 = b_7_6; // @[SingleLoop2.scala 18:15]
  assign io_OutMat_7_7 = b_7_7; // @[SingleLoop2.scala 18:15]
  assign io_Ovalid = _GEN_127 == 32'h4 | _T_9; // @[SingleLoop2.scala 26:53 28:19]
  assign io_ProcessValid = j == 32'h7; // @[SingleLoop2.scala 36:35]
  always @(posedge clock) begin
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_0_0 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h0 == io_IDex[2:0] & 3'h0 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_0_0 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_0_0 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_0_1 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h0 == io_IDex[2:0] & 3'h1 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_0_1 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_0_1 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_0_2 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h0 == io_IDex[2:0] & 3'h2 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_0_2 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_0_2 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_0_3 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h0 == io_IDex[2:0] & 3'h3 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_0_3 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_0_3 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_0_4 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h0 == io_IDex[2:0] & 3'h4 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_0_4 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_0_4 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_0_5 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h0 == io_IDex[2:0] & 3'h5 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_0_5 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_0_5 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_0_6 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h0 == io_IDex[2:0] & 3'h6 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_0_6 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_0_6 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_0_7 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h0 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_0_7 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_0_7 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_1_0 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h1 == io_IDex[2:0] & 3'h0 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_1_0 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_1_0 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_1_1 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h1 == io_IDex[2:0] & 3'h1 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_1_1 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_1_1 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_1_2 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h1 == io_IDex[2:0] & 3'h2 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_1_2 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_1_2 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_1_3 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h1 == io_IDex[2:0] & 3'h3 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_1_3 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_1_3 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_1_4 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h1 == io_IDex[2:0] & 3'h4 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_1_4 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_1_4 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_1_5 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h1 == io_IDex[2:0] & 3'h5 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_1_5 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_1_5 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_1_6 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h1 == io_IDex[2:0] & 3'h6 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_1_6 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_1_6 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_1_7 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h1 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_1_7 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_1_7 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_2_0 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h2 == io_IDex[2:0] & 3'h0 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_2_0 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_2_0 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_2_1 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h2 == io_IDex[2:0] & 3'h1 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_2_1 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_2_1 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_2_2 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h2 == io_IDex[2:0] & 3'h2 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_2_2 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_2_2 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_2_3 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h2 == io_IDex[2:0] & 3'h3 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_2_3 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_2_3 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_2_4 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h2 == io_IDex[2:0] & 3'h4 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_2_4 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_2_4 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_2_5 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h2 == io_IDex[2:0] & 3'h5 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_2_5 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_2_5 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_2_6 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h2 == io_IDex[2:0] & 3'h6 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_2_6 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_2_6 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_2_7 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h2 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_2_7 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_2_7 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_3_0 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h3 == io_IDex[2:0] & 3'h0 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_3_0 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_3_0 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_3_1 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h3 == io_IDex[2:0] & 3'h1 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_3_1 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_3_1 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_3_2 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h3 == io_IDex[2:0] & 3'h2 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_3_2 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_3_2 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_3_3 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h3 == io_IDex[2:0] & 3'h3 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_3_3 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_3_3 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_3_4 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h3 == io_IDex[2:0] & 3'h4 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_3_4 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_3_4 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_3_5 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h3 == io_IDex[2:0] & 3'h5 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_3_5 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_3_5 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_3_6 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h3 == io_IDex[2:0] & 3'h6 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_3_6 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_3_6 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_3_7 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h3 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_3_7 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_3_7 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_4_0 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h4 == io_IDex[2:0] & 3'h0 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_4_0 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_4_0 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_4_1 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h4 == io_IDex[2:0] & 3'h1 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_4_1 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_4_1 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_4_2 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h4 == io_IDex[2:0] & 3'h2 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_4_2 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_4_2 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_4_3 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h4 == io_IDex[2:0] & 3'h3 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_4_3 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_4_3 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_4_4 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h4 == io_IDex[2:0] & 3'h4 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_4_4 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_4_4 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_4_5 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h4 == io_IDex[2:0] & 3'h5 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_4_5 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_4_5 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_4_6 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h4 == io_IDex[2:0] & 3'h6 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_4_6 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_4_6 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_4_7 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h4 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_4_7 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_4_7 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_5_0 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h5 == io_IDex[2:0] & 3'h0 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_5_0 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_5_0 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_5_1 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h5 == io_IDex[2:0] & 3'h1 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_5_1 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_5_1 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_5_2 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h5 == io_IDex[2:0] & 3'h2 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_5_2 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_5_2 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_5_3 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h5 == io_IDex[2:0] & 3'h3 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_5_3 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_5_3 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_5_4 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h5 == io_IDex[2:0] & 3'h4 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_5_4 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_5_4 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_5_5 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h5 == io_IDex[2:0] & 3'h5 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_5_5 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_5_5 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_5_6 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h5 == io_IDex[2:0] & 3'h6 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_5_6 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_5_6 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_5_7 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h5 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_5_7 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_5_7 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_6_0 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h6 == io_IDex[2:0] & 3'h0 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_6_0 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_6_0 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_6_1 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h6 == io_IDex[2:0] & 3'h1 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_6_1 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_6_1 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_6_2 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h6 == io_IDex[2:0] & 3'h2 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_6_2 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_6_2 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_6_3 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h6 == io_IDex[2:0] & 3'h3 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_6_3 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_6_3 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_6_4 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h6 == io_IDex[2:0] & 3'h4 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_6_4 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_6_4 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_6_5 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h6 == io_IDex[2:0] & 3'h5 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_6_5 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_6_5 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_6_6 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h6 == io_IDex[2:0] & 3'h6 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_6_6 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_6_6 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_6_7 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h6 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_6_7 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_6_7 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_7_0 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h7 == io_IDex[2:0] & 3'h0 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_7_0 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_7_0 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_7_1 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h7 == io_IDex[2:0] & 3'h1 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_7_1 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_7_1 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_7_2 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h7 == io_IDex[2:0] & 3'h2 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_7_2 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_7_2 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_7_3 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h7 == io_IDex[2:0] & 3'h3 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_7_3 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_7_3 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_7_4 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h7 == io_IDex[2:0] & 3'h4 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_7_4 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_7_4 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_7_5 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h7 == io_IDex[2:0] & 3'h5 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_7_5 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_7_5 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_7_6 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h7 == io_IDex[2:0] & 3'h6 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_7_6 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_7_6 <= _GEN_126;
        end
      end
    end
    if (reset) begin // @[SingleLoop2.scala 17:20]
      b_7_7 <= 32'h0; // @[SingleLoop2.scala 17:20]
    end else if (io_valid) begin // @[SingleLoop2.scala 22:19]
      if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
        if (3'h7 == io_IDex[2:0] & 3'h7 == j[2:0]) begin // @[SingleLoop2.scala 23:19]
          b_7_7 <= io_mat_7_7; // @[SingleLoop2.scala 23:19]
        end else begin
          b_7_7 <= _GEN_126;
        end
      end
    end
    if (io_valid & j < 32'h7) begin // @[SingleLoop2.scala 39:50]
      j <= _j_T_1; // @[SingleLoop2.scala 40:11]
    end else if (!(_T_5)) begin // @[SingleLoop2.scala 41:43]
      if (!(_GEN_127 == 32'h4)) begin // @[SingleLoop2.scala 26:53]
        j <= io_JDex; // @[SingleLoop2.scala 20:7]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  b_0_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  b_0_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  b_0_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  b_0_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  b_0_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  b_0_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  b_0_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  b_0_7 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  b_1_0 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  b_1_1 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  b_1_2 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  b_1_3 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  b_1_4 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  b_1_5 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  b_1_6 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  b_1_7 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  b_2_0 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  b_2_1 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  b_2_2 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  b_2_3 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  b_2_4 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  b_2_5 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  b_2_6 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  b_2_7 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  b_3_0 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  b_3_1 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  b_3_2 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  b_3_3 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  b_3_4 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  b_3_5 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  b_3_6 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  b_3_7 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  b_4_0 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  b_4_1 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  b_4_2 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  b_4_3 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  b_4_4 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  b_4_5 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  b_4_6 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  b_4_7 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  b_5_0 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  b_5_1 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  b_5_2 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  b_5_3 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  b_5_4 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  b_5_5 = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  b_5_6 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  b_5_7 = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  b_6_0 = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  b_6_1 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  b_6_2 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  b_6_3 = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  b_6_4 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  b_6_5 = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  b_6_6 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  b_6_7 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  b_7_0 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  b_7_1 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  b_7_2 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  b_7_3 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  b_7_4 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  b_7_5 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  b_7_6 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  b_7_7 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  j = _RAND_64[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MergeDistribution2(
  input         clock,
  input         reset,
  input  [31:0] io_IDex,
  input  [31:0] io_mat_0_0,
  input  [31:0] io_mat_0_1,
  input  [31:0] io_mat_0_2,
  input  [31:0] io_mat_0_3,
  input  [31:0] io_mat_0_4,
  input  [31:0] io_mat_0_5,
  input  [31:0] io_mat_0_6,
  input  [31:0] io_mat_0_7,
  input  [31:0] io_mat_1_0,
  input  [31:0] io_mat_1_1,
  input  [31:0] io_mat_1_2,
  input  [31:0] io_mat_1_3,
  input  [31:0] io_mat_1_4,
  input  [31:0] io_mat_1_5,
  input  [31:0] io_mat_1_6,
  input  [31:0] io_mat_1_7,
  input  [31:0] io_mat_2_0,
  input  [31:0] io_mat_2_1,
  input  [31:0] io_mat_2_2,
  input  [31:0] io_mat_2_3,
  input  [31:0] io_mat_2_4,
  input  [31:0] io_mat_2_5,
  input  [31:0] io_mat_2_6,
  input  [31:0] io_mat_2_7,
  input  [31:0] io_mat_3_0,
  input  [31:0] io_mat_3_1,
  input  [31:0] io_mat_3_2,
  input  [31:0] io_mat_3_3,
  input  [31:0] io_mat_3_4,
  input  [31:0] io_mat_3_5,
  input  [31:0] io_mat_3_6,
  input  [31:0] io_mat_3_7,
  input  [31:0] io_mat_4_0,
  input  [31:0] io_mat_4_1,
  input  [31:0] io_mat_4_2,
  input  [31:0] io_mat_4_3,
  input  [31:0] io_mat_4_4,
  input  [31:0] io_mat_4_5,
  input  [31:0] io_mat_4_6,
  input  [31:0] io_mat_4_7,
  input  [31:0] io_mat_5_0,
  input  [31:0] io_mat_5_1,
  input  [31:0] io_mat_5_2,
  input  [31:0] io_mat_5_3,
  input  [31:0] io_mat_5_4,
  input  [31:0] io_mat_5_5,
  input  [31:0] io_mat_5_6,
  input  [31:0] io_mat_5_7,
  input  [31:0] io_mat_6_0,
  input  [31:0] io_mat_6_1,
  input  [31:0] io_mat_6_2,
  input  [31:0] io_mat_6_3,
  input  [31:0] io_mat_6_4,
  input  [31:0] io_mat_6_5,
  input  [31:0] io_mat_6_6,
  input  [31:0] io_mat_6_7,
  input  [31:0] io_mat_7_0,
  input  [31:0] io_mat_7_1,
  input  [31:0] io_mat_7_2,
  input  [31:0] io_mat_7_3,
  input  [31:0] io_mat_7_4,
  input  [31:0] io_mat_7_5,
  input  [31:0] io_mat_7_6,
  input  [31:0] io_mat_7_7,
  input         io_i_valid,
  output        io_valid,
  output [31:0] io_Omat_0_0,
  output [31:0] io_Omat_0_1,
  output [31:0] io_Omat_0_2,
  output [31:0] io_Omat_0_3,
  output [31:0] io_Omat_0_4,
  output [31:0] io_Omat_0_5,
  output [31:0] io_Omat_0_6,
  output [31:0] io_Omat_0_7,
  output [31:0] io_Omat_1_0,
  output [31:0] io_Omat_1_1,
  output [31:0] io_Omat_1_2,
  output [31:0] io_Omat_1_3,
  output [31:0] io_Omat_1_4,
  output [31:0] io_Omat_1_5,
  output [31:0] io_Omat_1_6,
  output [31:0] io_Omat_1_7,
  output [31:0] io_Omat_2_0,
  output [31:0] io_Omat_2_1,
  output [31:0] io_Omat_2_2,
  output [31:0] io_Omat_2_3,
  output [31:0] io_Omat_2_4,
  output [31:0] io_Omat_2_5,
  output [31:0] io_Omat_2_6,
  output [31:0] io_Omat_2_7,
  output [31:0] io_Omat_3_0,
  output [31:0] io_Omat_3_1,
  output [31:0] io_Omat_3_2,
  output [31:0] io_Omat_3_3,
  output [31:0] io_Omat_3_4,
  output [31:0] io_Omat_3_5,
  output [31:0] io_Omat_3_6,
  output [31:0] io_Omat_3_7,
  output [31:0] io_Omat_4_0,
  output [31:0] io_Omat_4_1,
  output [31:0] io_Omat_4_2,
  output [31:0] io_Omat_4_3,
  output [31:0] io_Omat_4_4,
  output [31:0] io_Omat_4_5,
  output [31:0] io_Omat_4_6,
  output [31:0] io_Omat_4_7,
  output [31:0] io_Omat_5_0,
  output [31:0] io_Omat_5_1,
  output [31:0] io_Omat_5_2,
  output [31:0] io_Omat_5_3,
  output [31:0] io_Omat_5_4,
  output [31:0] io_Omat_5_5,
  output [31:0] io_Omat_5_6,
  output [31:0] io_Omat_5_7,
  output [31:0] io_Omat_6_0,
  output [31:0] io_Omat_6_1,
  output [31:0] io_Omat_6_2,
  output [31:0] io_Omat_6_3,
  output [31:0] io_Omat_6_4,
  output [31:0] io_Omat_6_5,
  output [31:0] io_Omat_6_6,
  output [31:0] io_Omat_6_7,
  output [31:0] io_Omat_7_0,
  output [31:0] io_Omat_7_1,
  output [31:0] io_Omat_7_2,
  output [31:0] io_Omat_7_3,
  output [31:0] io_Omat_7_4,
  output [31:0] io_Omat_7_5,
  output [31:0] io_Omat_7_6,
  output [31:0] io_Omat_7_7
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] b_0_0; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_0_1; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_0_2; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_0_3; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_0_4; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_0_5; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_0_6; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_0_7; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_1_0; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_1_1; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_1_2; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_1_3; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_1_4; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_1_5; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_1_6; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_1_7; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_2_0; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_2_1; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_2_2; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_2_3; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_2_4; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_2_5; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_2_6; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_2_7; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_3_0; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_3_1; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_3_2; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_3_3; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_3_4; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_3_5; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_3_6; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_3_7; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_4_0; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_4_1; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_4_2; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_4_3; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_4_4; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_4_5; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_4_6; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_4_7; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_5_0; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_5_1; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_5_2; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_5_3; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_5_4; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_5_5; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_5_6; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_5_7; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_6_0; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_6_1; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_6_2; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_6_3; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_6_4; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_6_5; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_6_6; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_6_7; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_7_0; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_7_1; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_7_2; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_7_3; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_7_4; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_7_5; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_7_6; // @[MergeDistribution2.scala 16:18]
  reg [31:0] b_7_7; // @[MergeDistribution2.scala 16:18]
  reg [31:0] i; // @[MergeDistribution2.scala 21:18]
  reg [31:0] j; // @[MergeDistribution2.scala 22:18]
  wire [31:0] _i_T_1 = io_IDex + 32'h1; // @[MergeDistribution2.scala 30:16]
  wire  _GEN_276 = 3'h0 == i[2:0]; // @[MergeDistribution2.scala 34:{27,27}]
  wire  _GEN_277 = 3'h1 == j[2:0]; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_1 = 3'h0 == i[2:0] & 3'h1 == j[2:0] ? io_mat_0_1 : io_mat_0_0; // @[MergeDistribution2.scala 34:{27,27}]
  wire  _GEN_279 = 3'h2 == j[2:0]; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_2 = 3'h0 == i[2:0] & 3'h2 == j[2:0] ? io_mat_0_2 : _GEN_1; // @[MergeDistribution2.scala 34:{27,27}]
  wire  _GEN_281 = 3'h3 == j[2:0]; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_3 = 3'h0 == i[2:0] & 3'h3 == j[2:0] ? io_mat_0_3 : _GEN_2; // @[MergeDistribution2.scala 34:{27,27}]
  wire  _GEN_283 = 3'h4 == j[2:0]; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_4 = 3'h0 == i[2:0] & 3'h4 == j[2:0] ? io_mat_0_4 : _GEN_3; // @[MergeDistribution2.scala 34:{27,27}]
  wire  _GEN_285 = 3'h5 == j[2:0]; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_5 = 3'h0 == i[2:0] & 3'h5 == j[2:0] ? io_mat_0_5 : _GEN_4; // @[MergeDistribution2.scala 34:{27,27}]
  wire  _GEN_287 = 3'h6 == j[2:0]; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_6 = 3'h0 == i[2:0] & 3'h6 == j[2:0] ? io_mat_0_6 : _GEN_5; // @[MergeDistribution2.scala 34:{27,27}]
  wire  _GEN_289 = 3'h7 == j[2:0]; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_7 = 3'h0 == i[2:0] & 3'h7 == j[2:0] ? io_mat_0_7 : _GEN_6; // @[MergeDistribution2.scala 34:{27,27}]
  wire  _GEN_290 = 3'h1 == i[2:0]; // @[MergeDistribution2.scala 34:{27,27}]
  wire  _GEN_291 = 3'h0 == j[2:0]; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_8 = 3'h1 == i[2:0] & 3'h0 == j[2:0] ? io_mat_1_0 : _GEN_7; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_9 = 3'h1 == i[2:0] & 3'h1 == j[2:0] ? io_mat_1_1 : _GEN_8; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_10 = 3'h1 == i[2:0] & 3'h2 == j[2:0] ? io_mat_1_2 : _GEN_9; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_11 = 3'h1 == i[2:0] & 3'h3 == j[2:0] ? io_mat_1_3 : _GEN_10; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_12 = 3'h1 == i[2:0] & 3'h4 == j[2:0] ? io_mat_1_4 : _GEN_11; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_13 = 3'h1 == i[2:0] & 3'h5 == j[2:0] ? io_mat_1_5 : _GEN_12; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_14 = 3'h1 == i[2:0] & 3'h6 == j[2:0] ? io_mat_1_6 : _GEN_13; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_15 = 3'h1 == i[2:0] & 3'h7 == j[2:0] ? io_mat_1_7 : _GEN_14; // @[MergeDistribution2.scala 34:{27,27}]
  wire  _GEN_306 = 3'h2 == i[2:0]; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_16 = 3'h2 == i[2:0] & 3'h0 == j[2:0] ? io_mat_2_0 : _GEN_15; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_17 = 3'h2 == i[2:0] & 3'h1 == j[2:0] ? io_mat_2_1 : _GEN_16; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_18 = 3'h2 == i[2:0] & 3'h2 == j[2:0] ? io_mat_2_2 : _GEN_17; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_19 = 3'h2 == i[2:0] & 3'h3 == j[2:0] ? io_mat_2_3 : _GEN_18; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_20 = 3'h2 == i[2:0] & 3'h4 == j[2:0] ? io_mat_2_4 : _GEN_19; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_21 = 3'h2 == i[2:0] & 3'h5 == j[2:0] ? io_mat_2_5 : _GEN_20; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_22 = 3'h2 == i[2:0] & 3'h6 == j[2:0] ? io_mat_2_6 : _GEN_21; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_23 = 3'h2 == i[2:0] & 3'h7 == j[2:0] ? io_mat_2_7 : _GEN_22; // @[MergeDistribution2.scala 34:{27,27}]
  wire  _GEN_322 = 3'h3 == i[2:0]; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_24 = 3'h3 == i[2:0] & 3'h0 == j[2:0] ? io_mat_3_0 : _GEN_23; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_25 = 3'h3 == i[2:0] & 3'h1 == j[2:0] ? io_mat_3_1 : _GEN_24; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_26 = 3'h3 == i[2:0] & 3'h2 == j[2:0] ? io_mat_3_2 : _GEN_25; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_27 = 3'h3 == i[2:0] & 3'h3 == j[2:0] ? io_mat_3_3 : _GEN_26; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_28 = 3'h3 == i[2:0] & 3'h4 == j[2:0] ? io_mat_3_4 : _GEN_27; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_29 = 3'h3 == i[2:0] & 3'h5 == j[2:0] ? io_mat_3_5 : _GEN_28; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_30 = 3'h3 == i[2:0] & 3'h6 == j[2:0] ? io_mat_3_6 : _GEN_29; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_31 = 3'h3 == i[2:0] & 3'h7 == j[2:0] ? io_mat_3_7 : _GEN_30; // @[MergeDistribution2.scala 34:{27,27}]
  wire  _GEN_338 = 3'h4 == i[2:0]; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_32 = 3'h4 == i[2:0] & 3'h0 == j[2:0] ? io_mat_4_0 : _GEN_31; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_33 = 3'h4 == i[2:0] & 3'h1 == j[2:0] ? io_mat_4_1 : _GEN_32; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_34 = 3'h4 == i[2:0] & 3'h2 == j[2:0] ? io_mat_4_2 : _GEN_33; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_35 = 3'h4 == i[2:0] & 3'h3 == j[2:0] ? io_mat_4_3 : _GEN_34; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_36 = 3'h4 == i[2:0] & 3'h4 == j[2:0] ? io_mat_4_4 : _GEN_35; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_37 = 3'h4 == i[2:0] & 3'h5 == j[2:0] ? io_mat_4_5 : _GEN_36; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_38 = 3'h4 == i[2:0] & 3'h6 == j[2:0] ? io_mat_4_6 : _GEN_37; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_39 = 3'h4 == i[2:0] & 3'h7 == j[2:0] ? io_mat_4_7 : _GEN_38; // @[MergeDistribution2.scala 34:{27,27}]
  wire  _GEN_354 = 3'h5 == i[2:0]; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_40 = 3'h5 == i[2:0] & 3'h0 == j[2:0] ? io_mat_5_0 : _GEN_39; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_41 = 3'h5 == i[2:0] & 3'h1 == j[2:0] ? io_mat_5_1 : _GEN_40; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_42 = 3'h5 == i[2:0] & 3'h2 == j[2:0] ? io_mat_5_2 : _GEN_41; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_43 = 3'h5 == i[2:0] & 3'h3 == j[2:0] ? io_mat_5_3 : _GEN_42; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_44 = 3'h5 == i[2:0] & 3'h4 == j[2:0] ? io_mat_5_4 : _GEN_43; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_45 = 3'h5 == i[2:0] & 3'h5 == j[2:0] ? io_mat_5_5 : _GEN_44; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_46 = 3'h5 == i[2:0] & 3'h6 == j[2:0] ? io_mat_5_6 : _GEN_45; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_47 = 3'h5 == i[2:0] & 3'h7 == j[2:0] ? io_mat_5_7 : _GEN_46; // @[MergeDistribution2.scala 34:{27,27}]
  wire  _GEN_370 = 3'h6 == i[2:0]; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_48 = 3'h6 == i[2:0] & 3'h0 == j[2:0] ? io_mat_6_0 : _GEN_47; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_49 = 3'h6 == i[2:0] & 3'h1 == j[2:0] ? io_mat_6_1 : _GEN_48; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_50 = 3'h6 == i[2:0] & 3'h2 == j[2:0] ? io_mat_6_2 : _GEN_49; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_51 = 3'h6 == i[2:0] & 3'h3 == j[2:0] ? io_mat_6_3 : _GEN_50; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_52 = 3'h6 == i[2:0] & 3'h4 == j[2:0] ? io_mat_6_4 : _GEN_51; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_53 = 3'h6 == i[2:0] & 3'h5 == j[2:0] ? io_mat_6_5 : _GEN_52; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_54 = 3'h6 == i[2:0] & 3'h6 == j[2:0] ? io_mat_6_6 : _GEN_53; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_55 = 3'h6 == i[2:0] & 3'h7 == j[2:0] ? io_mat_6_7 : _GEN_54; // @[MergeDistribution2.scala 34:{27,27}]
  wire  _GEN_386 = 3'h7 == i[2:0]; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_56 = 3'h7 == i[2:0] & 3'h0 == j[2:0] ? io_mat_7_0 : _GEN_55; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_57 = 3'h7 == i[2:0] & 3'h1 == j[2:0] ? io_mat_7_1 : _GEN_56; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_58 = 3'h7 == i[2:0] & 3'h2 == j[2:0] ? io_mat_7_2 : _GEN_57; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_59 = 3'h7 == i[2:0] & 3'h3 == j[2:0] ? io_mat_7_3 : _GEN_58; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_60 = 3'h7 == i[2:0] & 3'h4 == j[2:0] ? io_mat_7_4 : _GEN_59; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_61 = 3'h7 == i[2:0] & 3'h5 == j[2:0] ? io_mat_7_5 : _GEN_60; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_62 = 3'h7 == i[2:0] & 3'h6 == j[2:0] ? io_mat_7_6 : _GEN_61; // @[MergeDistribution2.scala 34:{27,27}]
  wire [31:0] _GEN_63 = 3'h7 == i[2:0] & 3'h7 == j[2:0] ? io_mat_7_7 : _GEN_62; // @[MergeDistribution2.scala 34:{27,27}]
  wire  _T_7 = i < 32'h7; // @[MergeDistribution2.scala 39:16]
  wire  _T_8 = j == 32'h7; // @[MergeDistribution2.scala 39:46]
  wire [31:0] _i_T_3 = i + 32'h1; // @[MergeDistribution2.scala 40:14]
  wire  _T_10 = i == 32'h7; // @[MergeDistribution2.scala 44:17]
  wire  _T_11 = j < 32'h7; // @[MergeDistribution2.scala 44:51]
  wire [31:0] _j_T_1 = j + 32'h1; // @[MergeDistribution2.scala 47:12]
  wire  _T_15 = _T_10 & _T_8; // @[MergeDistribution2.scala 50:45]
  wire [31:0] _GEN_64 = _T_7 & _T_11 ? _j_T_1 : j; // @[MergeDistribution2.scala 22:18 55:74 56:9]
  wire [31:0] _GEN_68 = _T_10 & _T_8 ? j : _GEN_64; // @[MergeDistribution2.scala 50:80 54:9]
  wire [31:0] _GEN_70 = i == 32'h7 & j < 32'h7 ? _j_T_1 : _GEN_68; // @[MergeDistribution2.scala 44:77 47:7]
  wire  _GEN_71 = i == 32'h7 & j < 32'h7 ? 1'h0 : _T_15; // @[MergeDistribution2.scala 44:77 48:14]
  wire [31:0] _GEN_72 = i < 32'h7 & j == 32'h7 ? _i_T_3 : i; // @[MergeDistribution2.scala 39:74 40:9]
  wire [31:0] _GEN_73 = i < 32'h7 & j == 32'h7 ? 32'h0 : _GEN_70; // @[MergeDistribution2.scala 39:74 41:9]
  wire  _GEN_74 = i < 32'h7 & j == 32'h7 ? 1'h0 : _GEN_71; // @[MergeDistribution2.scala 39:74 42:16]
  wire  _GEN_77 = _GEN_63 == 32'h4 | _GEN_74; // @[MergeDistribution2.scala 34:36 37:16]
  wire  _GEN_80 = io_i_valid & i == 32'h0 & j == 32'h0 ? 1'h0 : _GEN_77; // @[MergeDistribution2.scala 29:47 32:14]
  assign io_valid = io_i_valid & _GEN_80; // @[MergeDistribution2.scala 26:20 62:14]
  assign io_Omat_0_0 = b_0_0; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_0_1 = b_0_1; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_0_2 = b_0_2; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_0_3 = b_0_3; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_0_4 = b_0_4; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_0_5 = b_0_5; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_0_6 = b_0_6; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_0_7 = b_0_7; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_1_0 = b_1_0; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_1_1 = b_1_1; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_1_2 = b_1_2; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_1_3 = b_1_3; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_1_4 = b_1_4; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_1_5 = b_1_5; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_1_6 = b_1_6; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_1_7 = b_1_7; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_2_0 = b_2_0; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_2_1 = b_2_1; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_2_2 = b_2_2; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_2_3 = b_2_3; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_2_4 = b_2_4; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_2_5 = b_2_5; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_2_6 = b_2_6; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_2_7 = b_2_7; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_3_0 = b_3_0; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_3_1 = b_3_1; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_3_2 = b_3_2; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_3_3 = b_3_3; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_3_4 = b_3_4; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_3_5 = b_3_5; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_3_6 = b_3_6; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_3_7 = b_3_7; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_4_0 = b_4_0; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_4_1 = b_4_1; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_4_2 = b_4_2; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_4_3 = b_4_3; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_4_4 = b_4_4; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_4_5 = b_4_5; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_4_6 = b_4_6; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_4_7 = b_4_7; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_5_0 = b_5_0; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_5_1 = b_5_1; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_5_2 = b_5_2; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_5_3 = b_5_3; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_5_4 = b_5_4; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_5_5 = b_5_5; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_5_6 = b_5_6; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_5_7 = b_5_7; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_6_0 = b_6_0; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_6_1 = b_6_1; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_6_2 = b_6_2; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_6_3 = b_6_3; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_6_4 = b_6_4; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_6_5 = b_6_5; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_6_6 = b_6_6; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_6_7 = b_6_7; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_7_0 = b_7_0; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_7_1 = b_7_1; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_7_2 = b_7_2; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_7_3 = b_7_3; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_7_4 = b_7_4; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_7_5 = b_7_5; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_7_6 = b_7_6; // @[MergeDistribution2.scala 17:11]
  assign io_Omat_7_7 = b_7_7; // @[MergeDistribution2.scala 17:11]
  always @(posedge clock) begin
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_0_0 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_276 & _GEN_291) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_0_0 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_0_0 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_0_1 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_276 & _GEN_277) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_0_1 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_0_1 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_0_2 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_276 & _GEN_279) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_0_2 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_0_2 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_0_3 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_276 & _GEN_281) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_0_3 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_0_3 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_0_4 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_276 & _GEN_283) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_0_4 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_0_4 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_0_5 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_276 & _GEN_285) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_0_5 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_0_5 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_0_6 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_276 & _GEN_287) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_0_6 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_0_6 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_0_7 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_276 & _GEN_289) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_0_7 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_0_7 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_1_0 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_290 & _GEN_291) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_1_0 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_1_0 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_1_1 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_290 & _GEN_277) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_1_1 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_1_1 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_1_2 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_290 & _GEN_279) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_1_2 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_1_2 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_1_3 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_290 & _GEN_281) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_1_3 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_1_3 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_1_4 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_290 & _GEN_283) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_1_4 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_1_4 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_1_5 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_290 & _GEN_285) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_1_5 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_1_5 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_1_6 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_290 & _GEN_287) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_1_6 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_1_6 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_1_7 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_290 & _GEN_289) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_1_7 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_1_7 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_2_0 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_306 & _GEN_291) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_2_0 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_2_0 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_2_1 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_306 & _GEN_277) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_2_1 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_2_1 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_2_2 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_306 & _GEN_279) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_2_2 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_2_2 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_2_3 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_306 & _GEN_281) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_2_3 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_2_3 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_2_4 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_306 & _GEN_283) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_2_4 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_2_4 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_2_5 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_306 & _GEN_285) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_2_5 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_2_5 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_2_6 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_306 & _GEN_287) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_2_6 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_2_6 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_2_7 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_306 & _GEN_289) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_2_7 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_2_7 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_3_0 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_322 & _GEN_291) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_3_0 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_3_0 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_3_1 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_322 & _GEN_277) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_3_1 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_3_1 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_3_2 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_322 & _GEN_279) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_3_2 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_3_2 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_3_3 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_322 & _GEN_281) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_3_3 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_3_3 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_3_4 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_322 & _GEN_283) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_3_4 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_3_4 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_3_5 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_322 & _GEN_285) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_3_5 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_3_5 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_3_6 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_322 & _GEN_287) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_3_6 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_3_6 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_3_7 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_322 & _GEN_289) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_3_7 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_3_7 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_4_0 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_338 & _GEN_291) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_4_0 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_4_0 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_4_1 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_338 & _GEN_277) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_4_1 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_4_1 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_4_2 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_338 & _GEN_279) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_4_2 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_4_2 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_4_3 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_338 & _GEN_281) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_4_3 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_4_3 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_4_4 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_338 & _GEN_283) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_4_4 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_4_4 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_4_5 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_338 & _GEN_285) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_4_5 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_4_5 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_4_6 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_338 & _GEN_287) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_4_6 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_4_6 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_4_7 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_338 & _GEN_289) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_4_7 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_4_7 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_5_0 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_354 & _GEN_291) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_5_0 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_5_0 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_5_1 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_354 & _GEN_277) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_5_1 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_5_1 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_5_2 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_354 & _GEN_279) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_5_2 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_5_2 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_5_3 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_354 & _GEN_281) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_5_3 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_5_3 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_5_4 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_354 & _GEN_283) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_5_4 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_5_4 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_5_5 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_354 & _GEN_285) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_5_5 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_5_5 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_5_6 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_354 & _GEN_287) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_5_6 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_5_6 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_5_7 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_354 & _GEN_289) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_5_7 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_5_7 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_6_0 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_370 & _GEN_291) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_6_0 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_6_0 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_6_1 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_370 & _GEN_277) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_6_1 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_6_1 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_6_2 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_370 & _GEN_279) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_6_2 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_6_2 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_6_3 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_370 & _GEN_281) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_6_3 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_6_3 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_6_4 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_370 & _GEN_283) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_6_4 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_6_4 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_6_5 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_370 & _GEN_285) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_6_5 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_6_5 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_6_6 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_370 & _GEN_287) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_6_6 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_6_6 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_6_7 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_370 & _GEN_289) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_6_7 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_6_7 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_7_0 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_386 & _GEN_291) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_7_0 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_7_0 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_7_1 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_386 & _GEN_277) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_7_1 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_7_1 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_7_2 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_386 & _GEN_279) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_7_2 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_7_2 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_7_3 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_386 & _GEN_281) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_7_3 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_7_3 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_7_4 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_386 & _GEN_283) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_7_4 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_7_4 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_7_5 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_386 & _GEN_285) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_7_5 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_7_5 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_7_6 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_386 & _GEN_287) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_7_6 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_7_6 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 16:18]
      b_7_7 <= 32'h0; // @[MergeDistribution2.scala 16:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (_GEN_386 & _GEN_289) begin // @[MergeDistribution2.scala 60:13]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[MergeDistribution2.scala 34:27]
          b_7_7 <= io_mat_7_7; // @[MergeDistribution2.scala 34:27]
        end else begin
          b_7_7 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 21:18]
      i <= 32'h0; // @[MergeDistribution2.scala 21:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (io_i_valid & i == 32'h0 & j == 32'h0) begin // @[MergeDistribution2.scala 29:47]
        i <= _i_T_1; // @[MergeDistribution2.scala 30:5]
      end else if (!(_GEN_63 == 32'h4)) begin // @[MergeDistribution2.scala 34:36]
        i <= _GEN_72;
      end
    end
    if (reset) begin // @[MergeDistribution2.scala 22:18]
      j <= 32'h0; // @[MergeDistribution2.scala 22:18]
    end else if (io_i_valid) begin // @[MergeDistribution2.scala 26:20]
      if (io_i_valid & i == 32'h0 & j == 32'h0) begin // @[MergeDistribution2.scala 29:47]
        j <= 32'h0; // @[MergeDistribution2.scala 31:7]
      end else if (!(_GEN_63 == 32'h4)) begin // @[MergeDistribution2.scala 34:36]
        j <= _GEN_73;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  b_0_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  b_0_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  b_0_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  b_0_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  b_0_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  b_0_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  b_0_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  b_0_7 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  b_1_0 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  b_1_1 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  b_1_2 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  b_1_3 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  b_1_4 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  b_1_5 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  b_1_6 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  b_1_7 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  b_2_0 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  b_2_1 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  b_2_2 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  b_2_3 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  b_2_4 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  b_2_5 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  b_2_6 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  b_2_7 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  b_3_0 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  b_3_1 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  b_3_2 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  b_3_3 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  b_3_4 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  b_3_5 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  b_3_6 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  b_3_7 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  b_4_0 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  b_4_1 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  b_4_2 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  b_4_3 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  b_4_4 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  b_4_5 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  b_4_6 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  b_4_7 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  b_5_0 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  b_5_1 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  b_5_2 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  b_5_3 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  b_5_4 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  b_5_5 = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  b_5_6 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  b_5_7 = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  b_6_0 = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  b_6_1 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  b_6_2 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  b_6_3 = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  b_6_4 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  b_6_5 = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  b_6_6 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  b_6_7 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  b_7_0 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  b_7_1 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  b_7_2 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  b_7_3 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  b_7_4 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  b_7_5 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  b_7_6 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  b_7_7 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  i = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  j = _RAND_65[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FinalMerge(
  input         clock,
  input         reset,
  input  [31:0] io_IDex,
  input  [31:0] io_PreMat_0_0,
  input  [31:0] io_PreMat_0_1,
  input  [31:0] io_PreMat_0_2,
  input  [31:0] io_PreMat_0_3,
  input  [31:0] io_PreMat_0_4,
  input  [31:0] io_PreMat_0_5,
  input  [31:0] io_PreMat_0_6,
  input  [31:0] io_PreMat_0_7,
  input  [31:0] io_PreMat_1_0,
  input  [31:0] io_PreMat_1_1,
  input  [31:0] io_PreMat_1_2,
  input  [31:0] io_PreMat_1_3,
  input  [31:0] io_PreMat_1_4,
  input  [31:0] io_PreMat_1_5,
  input  [31:0] io_PreMat_1_6,
  input  [31:0] io_PreMat_1_7,
  input  [31:0] io_PreMat_2_0,
  input  [31:0] io_PreMat_2_1,
  input  [31:0] io_PreMat_2_2,
  input  [31:0] io_PreMat_2_3,
  input  [31:0] io_PreMat_2_4,
  input  [31:0] io_PreMat_2_5,
  input  [31:0] io_PreMat_2_6,
  input  [31:0] io_PreMat_2_7,
  input  [31:0] io_PreMat_3_0,
  input  [31:0] io_PreMat_3_1,
  input  [31:0] io_PreMat_3_2,
  input  [31:0] io_PreMat_3_3,
  input  [31:0] io_PreMat_3_4,
  input  [31:0] io_PreMat_3_5,
  input  [31:0] io_PreMat_3_6,
  input  [31:0] io_PreMat_3_7,
  input  [31:0] io_PreMat_4_0,
  input  [31:0] io_PreMat_4_1,
  input  [31:0] io_PreMat_4_2,
  input  [31:0] io_PreMat_4_3,
  input  [31:0] io_PreMat_4_4,
  input  [31:0] io_PreMat_4_5,
  input  [31:0] io_PreMat_4_6,
  input  [31:0] io_PreMat_4_7,
  input  [31:0] io_PreMat_5_0,
  input  [31:0] io_PreMat_5_1,
  input  [31:0] io_PreMat_5_2,
  input  [31:0] io_PreMat_5_3,
  input  [31:0] io_PreMat_5_4,
  input  [31:0] io_PreMat_5_5,
  input  [31:0] io_PreMat_5_6,
  input  [31:0] io_PreMat_5_7,
  input  [31:0] io_PreMat_6_0,
  input  [31:0] io_PreMat_6_1,
  input  [31:0] io_PreMat_6_2,
  input  [31:0] io_PreMat_6_3,
  input  [31:0] io_PreMat_6_4,
  input  [31:0] io_PreMat_6_5,
  input  [31:0] io_PreMat_6_6,
  input  [31:0] io_PreMat_6_7,
  input  [31:0] io_PreMat_7_0,
  input  [31:0] io_PreMat_7_1,
  input  [31:0] io_PreMat_7_2,
  input  [31:0] io_PreMat_7_3,
  input  [31:0] io_PreMat_7_4,
  input  [31:0] io_PreMat_7_5,
  input  [31:0] io_PreMat_7_6,
  input  [31:0] io_PreMat_7_7,
  input  [31:0] io_lastMat_0_0,
  input  [31:0] io_lastMat_0_1,
  input  [31:0] io_lastMat_0_2,
  input  [31:0] io_lastMat_0_3,
  input  [31:0] io_lastMat_0_4,
  input  [31:0] io_lastMat_0_5,
  input  [31:0] io_lastMat_0_6,
  input  [31:0] io_lastMat_0_7,
  input  [31:0] io_lastMat_1_0,
  input  [31:0] io_lastMat_1_1,
  input  [31:0] io_lastMat_1_2,
  input  [31:0] io_lastMat_1_3,
  input  [31:0] io_lastMat_1_4,
  input  [31:0] io_lastMat_1_5,
  input  [31:0] io_lastMat_1_6,
  input  [31:0] io_lastMat_1_7,
  input  [31:0] io_lastMat_2_0,
  input  [31:0] io_lastMat_2_1,
  input  [31:0] io_lastMat_2_2,
  input  [31:0] io_lastMat_2_3,
  input  [31:0] io_lastMat_2_4,
  input  [31:0] io_lastMat_2_5,
  input  [31:0] io_lastMat_2_6,
  input  [31:0] io_lastMat_2_7,
  input  [31:0] io_lastMat_3_0,
  input  [31:0] io_lastMat_3_1,
  input  [31:0] io_lastMat_3_2,
  input  [31:0] io_lastMat_3_3,
  input  [31:0] io_lastMat_3_4,
  input  [31:0] io_lastMat_3_5,
  input  [31:0] io_lastMat_3_6,
  input  [31:0] io_lastMat_3_7,
  input  [31:0] io_lastMat_4_0,
  input  [31:0] io_lastMat_4_1,
  input  [31:0] io_lastMat_4_2,
  input  [31:0] io_lastMat_4_3,
  input  [31:0] io_lastMat_4_4,
  input  [31:0] io_lastMat_4_5,
  input  [31:0] io_lastMat_4_6,
  input  [31:0] io_lastMat_4_7,
  input  [31:0] io_lastMat_5_0,
  input  [31:0] io_lastMat_5_1,
  input  [31:0] io_lastMat_5_2,
  input  [31:0] io_lastMat_5_3,
  input  [31:0] io_lastMat_5_4,
  input  [31:0] io_lastMat_5_5,
  input  [31:0] io_lastMat_5_6,
  input  [31:0] io_lastMat_5_7,
  input  [31:0] io_lastMat_6_0,
  input  [31:0] io_lastMat_6_1,
  input  [31:0] io_lastMat_6_2,
  input  [31:0] io_lastMat_6_3,
  input  [31:0] io_lastMat_6_4,
  input  [31:0] io_lastMat_6_5,
  input  [31:0] io_lastMat_6_6,
  input  [31:0] io_lastMat_6_7,
  input  [31:0] io_lastMat_7_0,
  input  [31:0] io_lastMat_7_1,
  input  [31:0] io_lastMat_7_2,
  input  [31:0] io_lastMat_7_3,
  input  [31:0] io_lastMat_7_4,
  input  [31:0] io_lastMat_7_5,
  input  [31:0] io_lastMat_7_6,
  input  [31:0] io_lastMat_7_7,
  input         io_valid,
  output        io_Ovalid,
  output [31:0] io_omat_0_0,
  output [31:0] io_omat_0_1,
  output [31:0] io_omat_0_2,
  output [31:0] io_omat_0_3,
  output [31:0] io_omat_0_4,
  output [31:0] io_omat_0_5,
  output [31:0] io_omat_0_6,
  output [31:0] io_omat_0_7,
  output [31:0] io_omat_1_0,
  output [31:0] io_omat_1_1,
  output [31:0] io_omat_1_2,
  output [31:0] io_omat_1_3,
  output [31:0] io_omat_1_4,
  output [31:0] io_omat_1_5,
  output [31:0] io_omat_1_6,
  output [31:0] io_omat_1_7,
  output [31:0] io_omat_2_0,
  output [31:0] io_omat_2_1,
  output [31:0] io_omat_2_2,
  output [31:0] io_omat_2_3,
  output [31:0] io_omat_2_4,
  output [31:0] io_omat_2_5,
  output [31:0] io_omat_2_6,
  output [31:0] io_omat_2_7,
  output [31:0] io_omat_3_0,
  output [31:0] io_omat_3_1,
  output [31:0] io_omat_3_2,
  output [31:0] io_omat_3_3,
  output [31:0] io_omat_3_4,
  output [31:0] io_omat_3_5,
  output [31:0] io_omat_3_6,
  output [31:0] io_omat_3_7,
  output [31:0] io_omat_4_0,
  output [31:0] io_omat_4_1,
  output [31:0] io_omat_4_2,
  output [31:0] io_omat_4_3,
  output [31:0] io_omat_4_4,
  output [31:0] io_omat_4_5,
  output [31:0] io_omat_4_6,
  output [31:0] io_omat_4_7,
  output [31:0] io_omat_5_0,
  output [31:0] io_omat_5_1,
  output [31:0] io_omat_5_2,
  output [31:0] io_omat_5_3,
  output [31:0] io_omat_5_4,
  output [31:0] io_omat_5_5,
  output [31:0] io_omat_5_6,
  output [31:0] io_omat_5_7,
  output [31:0] io_omat_6_0,
  output [31:0] io_omat_6_1,
  output [31:0] io_omat_6_2,
  output [31:0] io_omat_6_3,
  output [31:0] io_omat_6_4,
  output [31:0] io_omat_6_5,
  output [31:0] io_omat_6_6,
  output [31:0] io_omat_6_7,
  output [31:0] io_omat_7_0,
  output [31:0] io_omat_7_1,
  output [31:0] io_omat_7_2,
  output [31:0] io_omat_7_3,
  output [31:0] io_omat_7_4,
  output [31:0] io_omat_7_5,
  output [31:0] io_omat_7_6,
  output [31:0] io_omat_7_7
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] mat_0_0; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_0_1; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_0_2; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_0_3; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_0_4; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_0_5; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_0_6; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_0_7; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_1_0; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_1_1; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_1_2; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_1_3; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_1_4; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_1_5; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_1_6; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_1_7; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_2_0; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_2_1; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_2_2; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_2_3; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_2_4; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_2_5; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_2_6; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_2_7; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_3_0; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_3_1; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_3_2; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_3_3; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_3_4; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_3_5; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_3_6; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_3_7; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_4_0; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_4_1; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_4_2; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_4_3; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_4_4; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_4_5; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_4_6; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_4_7; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_5_0; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_5_1; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_5_2; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_5_3; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_5_4; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_5_5; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_5_6; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_5_7; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_6_0; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_6_1; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_6_2; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_6_3; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_6_4; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_6_5; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_6_6; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_6_7; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_7_0; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_7_1; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_7_2; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_7_3; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_7_4; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_7_5; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_7_6; // @[FinalMerge.scala 16:22]
  reg [31:0] mat_7_7; // @[FinalMerge.scala 16:22]
  reg [31:0] i; // @[FinalMerge.scala 20:20]
  reg [31:0] j; // @[FinalMerge.scala 21:20]
  wire [31:0] _GEN_9 = 3'h1 == io_IDex[2:0] ? io_PreMat_1_0 : io_PreMat_0_0; // @[FinalMerge.scala 25:{25,25}]
  wire [31:0] _GEN_10 = 3'h2 == io_IDex[2:0] ? io_PreMat_2_0 : _GEN_9; // @[FinalMerge.scala 25:{25,25}]
  wire [31:0] _GEN_11 = 3'h3 == io_IDex[2:0] ? io_PreMat_3_0 : _GEN_10; // @[FinalMerge.scala 25:{25,25}]
  wire [31:0] _GEN_12 = 3'h4 == io_IDex[2:0] ? io_PreMat_4_0 : _GEN_11; // @[FinalMerge.scala 25:{25,25}]
  wire [31:0] _GEN_13 = 3'h5 == io_IDex[2:0] ? io_PreMat_5_0 : _GEN_12; // @[FinalMerge.scala 25:{25,25}]
  wire [31:0] _GEN_14 = 3'h6 == io_IDex[2:0] ? io_PreMat_6_0 : _GEN_13; // @[FinalMerge.scala 25:{25,25}]
  wire [31:0] _GEN_15 = 3'h7 == io_IDex[2:0] ? io_PreMat_7_0 : _GEN_14; // @[FinalMerge.scala 25:{25,25}]
  wire [31:0] _GEN_0 = 3'h0 == io_IDex[2:0] ? _GEN_15 : mat_0_0; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_1 = 3'h1 == io_IDex[2:0] ? _GEN_15 : mat_1_0; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_2 = 3'h2 == io_IDex[2:0] ? _GEN_15 : mat_2_0; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_3 = 3'h3 == io_IDex[2:0] ? _GEN_15 : mat_3_0; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_4 = 3'h4 == io_IDex[2:0] ? _GEN_15 : mat_4_0; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_5 = 3'h5 == io_IDex[2:0] ? _GEN_15 : mat_5_0; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_6 = 3'h6 == io_IDex[2:0] ? _GEN_15 : mat_6_0; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_7 = 3'h7 == io_IDex[2:0] ? _GEN_15 : mat_7_0; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_25 = 3'h1 == io_IDex[2:0] ? io_PreMat_1_1 : io_PreMat_0_1; // @[FinalMerge.scala 25:{25,25}]
  wire [31:0] _GEN_26 = 3'h2 == io_IDex[2:0] ? io_PreMat_2_1 : _GEN_25; // @[FinalMerge.scala 25:{25,25}]
  wire [31:0] _GEN_27 = 3'h3 == io_IDex[2:0] ? io_PreMat_3_1 : _GEN_26; // @[FinalMerge.scala 25:{25,25}]
  wire [31:0] _GEN_28 = 3'h4 == io_IDex[2:0] ? io_PreMat_4_1 : _GEN_27; // @[FinalMerge.scala 25:{25,25}]
  wire [31:0] _GEN_29 = 3'h5 == io_IDex[2:0] ? io_PreMat_5_1 : _GEN_28; // @[FinalMerge.scala 25:{25,25}]
  wire [31:0] _GEN_30 = 3'h6 == io_IDex[2:0] ? io_PreMat_6_1 : _GEN_29; // @[FinalMerge.scala 25:{25,25}]
  wire [31:0] _GEN_31 = 3'h7 == io_IDex[2:0] ? io_PreMat_7_1 : _GEN_30; // @[FinalMerge.scala 25:{25,25}]
  wire [31:0] _GEN_16 = 3'h0 == io_IDex[2:0] ? _GEN_31 : mat_0_1; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_17 = 3'h1 == io_IDex[2:0] ? _GEN_31 : mat_1_1; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_18 = 3'h2 == io_IDex[2:0] ? _GEN_31 : mat_2_1; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_19 = 3'h3 == io_IDex[2:0] ? _GEN_31 : mat_3_1; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_20 = 3'h4 == io_IDex[2:0] ? _GEN_31 : mat_4_1; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_21 = 3'h5 == io_IDex[2:0] ? _GEN_31 : mat_5_1; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_22 = 3'h6 == io_IDex[2:0] ? _GEN_31 : mat_6_1; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_23 = 3'h7 == io_IDex[2:0] ? _GEN_31 : mat_7_1; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_41 = 3'h1 == io_IDex[2:0] ? io_PreMat_1_2 : io_PreMat_0_2; // @[FinalMerge.scala 25:{25,25}]
  wire [31:0] _GEN_42 = 3'h2 == io_IDex[2:0] ? io_PreMat_2_2 : _GEN_41; // @[FinalMerge.scala 25:{25,25}]
  wire [31:0] _GEN_43 = 3'h3 == io_IDex[2:0] ? io_PreMat_3_2 : _GEN_42; // @[FinalMerge.scala 25:{25,25}]
  wire [31:0] _GEN_44 = 3'h4 == io_IDex[2:0] ? io_PreMat_4_2 : _GEN_43; // @[FinalMerge.scala 25:{25,25}]
  wire [31:0] _GEN_45 = 3'h5 == io_IDex[2:0] ? io_PreMat_5_2 : _GEN_44; // @[FinalMerge.scala 25:{25,25}]
  wire [31:0] _GEN_46 = 3'h6 == io_IDex[2:0] ? io_PreMat_6_2 : _GEN_45; // @[FinalMerge.scala 25:{25,25}]
  wire [31:0] _GEN_47 = 3'h7 == io_IDex[2:0] ? io_PreMat_7_2 : _GEN_46; // @[FinalMerge.scala 25:{25,25}]
  wire [31:0] _GEN_32 = 3'h0 == io_IDex[2:0] ? _GEN_47 : mat_0_2; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_33 = 3'h1 == io_IDex[2:0] ? _GEN_47 : mat_1_2; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_34 = 3'h2 == io_IDex[2:0] ? _GEN_47 : mat_2_2; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_35 = 3'h3 == io_IDex[2:0] ? _GEN_47 : mat_3_2; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_36 = 3'h4 == io_IDex[2:0] ? _GEN_47 : mat_4_2; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_37 = 3'h5 == io_IDex[2:0] ? _GEN_47 : mat_5_2; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_38 = 3'h6 == io_IDex[2:0] ? _GEN_47 : mat_6_2; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_39 = 3'h7 == io_IDex[2:0] ? _GEN_47 : mat_7_2; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_57 = 3'h1 == io_IDex[2:0] ? io_PreMat_1_3 : io_PreMat_0_3; // @[FinalMerge.scala 25:{25,25}]
  wire [31:0] _GEN_58 = 3'h2 == io_IDex[2:0] ? io_PreMat_2_3 : _GEN_57; // @[FinalMerge.scala 25:{25,25}]
  wire [31:0] _GEN_59 = 3'h3 == io_IDex[2:0] ? io_PreMat_3_3 : _GEN_58; // @[FinalMerge.scala 25:{25,25}]
  wire [31:0] _GEN_60 = 3'h4 == io_IDex[2:0] ? io_PreMat_4_3 : _GEN_59; // @[FinalMerge.scala 25:{25,25}]
  wire [31:0] _GEN_61 = 3'h5 == io_IDex[2:0] ? io_PreMat_5_3 : _GEN_60; // @[FinalMerge.scala 25:{25,25}]
  wire [31:0] _GEN_62 = 3'h6 == io_IDex[2:0] ? io_PreMat_6_3 : _GEN_61; // @[FinalMerge.scala 25:{25,25}]
  wire [31:0] _GEN_63 = 3'h7 == io_IDex[2:0] ? io_PreMat_7_3 : _GEN_62; // @[FinalMerge.scala 25:{25,25}]
  wire [31:0] _GEN_48 = 3'h0 == io_IDex[2:0] ? _GEN_63 : mat_0_3; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_49 = 3'h1 == io_IDex[2:0] ? _GEN_63 : mat_1_3; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_50 = 3'h2 == io_IDex[2:0] ? _GEN_63 : mat_2_3; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_51 = 3'h3 == io_IDex[2:0] ? _GEN_63 : mat_3_3; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_52 = 3'h4 == io_IDex[2:0] ? _GEN_63 : mat_4_3; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_53 = 3'h5 == io_IDex[2:0] ? _GEN_63 : mat_5_3; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_54 = 3'h6 == io_IDex[2:0] ? _GEN_63 : mat_6_3; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_55 = 3'h7 == io_IDex[2:0] ? _GEN_63 : mat_7_3; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_73 = 3'h1 == io_IDex[2:0] ? io_PreMat_1_4 : io_PreMat_0_4; // @[FinalMerge.scala 25:{25,25}]
  wire [31:0] _GEN_74 = 3'h2 == io_IDex[2:0] ? io_PreMat_2_4 : _GEN_73; // @[FinalMerge.scala 25:{25,25}]
  wire [31:0] _GEN_75 = 3'h3 == io_IDex[2:0] ? io_PreMat_3_4 : _GEN_74; // @[FinalMerge.scala 25:{25,25}]
  wire [31:0] _GEN_76 = 3'h4 == io_IDex[2:0] ? io_PreMat_4_4 : _GEN_75; // @[FinalMerge.scala 25:{25,25}]
  wire [31:0] _GEN_77 = 3'h5 == io_IDex[2:0] ? io_PreMat_5_4 : _GEN_76; // @[FinalMerge.scala 25:{25,25}]
  wire [31:0] _GEN_78 = 3'h6 == io_IDex[2:0] ? io_PreMat_6_4 : _GEN_77; // @[FinalMerge.scala 25:{25,25}]
  wire [31:0] _GEN_79 = 3'h7 == io_IDex[2:0] ? io_PreMat_7_4 : _GEN_78; // @[FinalMerge.scala 25:{25,25}]
  wire [31:0] _GEN_64 = 3'h0 == io_IDex[2:0] ? _GEN_79 : mat_0_4; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_65 = 3'h1 == io_IDex[2:0] ? _GEN_79 : mat_1_4; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_66 = 3'h2 == io_IDex[2:0] ? _GEN_79 : mat_2_4; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_67 = 3'h3 == io_IDex[2:0] ? _GEN_79 : mat_3_4; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_68 = 3'h4 == io_IDex[2:0] ? _GEN_79 : mat_4_4; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_69 = 3'h5 == io_IDex[2:0] ? _GEN_79 : mat_5_4; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_70 = 3'h6 == io_IDex[2:0] ? _GEN_79 : mat_6_4; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_71 = 3'h7 == io_IDex[2:0] ? _GEN_79 : mat_7_4; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_89 = 3'h1 == io_IDex[2:0] ? io_PreMat_1_5 : io_PreMat_0_5; // @[FinalMerge.scala 25:{25,25}]
  wire [31:0] _GEN_90 = 3'h2 == io_IDex[2:0] ? io_PreMat_2_5 : _GEN_89; // @[FinalMerge.scala 25:{25,25}]
  wire [31:0] _GEN_91 = 3'h3 == io_IDex[2:0] ? io_PreMat_3_5 : _GEN_90; // @[FinalMerge.scala 25:{25,25}]
  wire [31:0] _GEN_92 = 3'h4 == io_IDex[2:0] ? io_PreMat_4_5 : _GEN_91; // @[FinalMerge.scala 25:{25,25}]
  wire [31:0] _GEN_93 = 3'h5 == io_IDex[2:0] ? io_PreMat_5_5 : _GEN_92; // @[FinalMerge.scala 25:{25,25}]
  wire [31:0] _GEN_94 = 3'h6 == io_IDex[2:0] ? io_PreMat_6_5 : _GEN_93; // @[FinalMerge.scala 25:{25,25}]
  wire [31:0] _GEN_95 = 3'h7 == io_IDex[2:0] ? io_PreMat_7_5 : _GEN_94; // @[FinalMerge.scala 25:{25,25}]
  wire [31:0] _GEN_80 = 3'h0 == io_IDex[2:0] ? _GEN_95 : mat_0_5; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_81 = 3'h1 == io_IDex[2:0] ? _GEN_95 : mat_1_5; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_82 = 3'h2 == io_IDex[2:0] ? _GEN_95 : mat_2_5; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_83 = 3'h3 == io_IDex[2:0] ? _GEN_95 : mat_3_5; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_84 = 3'h4 == io_IDex[2:0] ? _GEN_95 : mat_4_5; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_85 = 3'h5 == io_IDex[2:0] ? _GEN_95 : mat_5_5; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_86 = 3'h6 == io_IDex[2:0] ? _GEN_95 : mat_6_5; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_87 = 3'h7 == io_IDex[2:0] ? _GEN_95 : mat_7_5; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_105 = 3'h1 == io_IDex[2:0] ? io_PreMat_1_6 : io_PreMat_0_6; // @[FinalMerge.scala 25:{25,25}]
  wire [31:0] _GEN_106 = 3'h2 == io_IDex[2:0] ? io_PreMat_2_6 : _GEN_105; // @[FinalMerge.scala 25:{25,25}]
  wire [31:0] _GEN_107 = 3'h3 == io_IDex[2:0] ? io_PreMat_3_6 : _GEN_106; // @[FinalMerge.scala 25:{25,25}]
  wire [31:0] _GEN_108 = 3'h4 == io_IDex[2:0] ? io_PreMat_4_6 : _GEN_107; // @[FinalMerge.scala 25:{25,25}]
  wire [31:0] _GEN_109 = 3'h5 == io_IDex[2:0] ? io_PreMat_5_6 : _GEN_108; // @[FinalMerge.scala 25:{25,25}]
  wire [31:0] _GEN_110 = 3'h6 == io_IDex[2:0] ? io_PreMat_6_6 : _GEN_109; // @[FinalMerge.scala 25:{25,25}]
  wire [31:0] _GEN_111 = 3'h7 == io_IDex[2:0] ? io_PreMat_7_6 : _GEN_110; // @[FinalMerge.scala 25:{25,25}]
  wire [31:0] _GEN_96 = 3'h0 == io_IDex[2:0] ? _GEN_111 : mat_0_6; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_97 = 3'h1 == io_IDex[2:0] ? _GEN_111 : mat_1_6; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_98 = 3'h2 == io_IDex[2:0] ? _GEN_111 : mat_2_6; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_99 = 3'h3 == io_IDex[2:0] ? _GEN_111 : mat_3_6; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_100 = 3'h4 == io_IDex[2:0] ? _GEN_111 : mat_4_6; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_101 = 3'h5 == io_IDex[2:0] ? _GEN_111 : mat_5_6; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_102 = 3'h6 == io_IDex[2:0] ? _GEN_111 : mat_6_6; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_103 = 3'h7 == io_IDex[2:0] ? _GEN_111 : mat_7_6; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_121 = 3'h1 == io_IDex[2:0] ? io_PreMat_1_7 : io_PreMat_0_7; // @[FinalMerge.scala 25:{25,25}]
  wire [31:0] _GEN_122 = 3'h2 == io_IDex[2:0] ? io_PreMat_2_7 : _GEN_121; // @[FinalMerge.scala 25:{25,25}]
  wire [31:0] _GEN_123 = 3'h3 == io_IDex[2:0] ? io_PreMat_3_7 : _GEN_122; // @[FinalMerge.scala 25:{25,25}]
  wire [31:0] _GEN_124 = 3'h4 == io_IDex[2:0] ? io_PreMat_4_7 : _GEN_123; // @[FinalMerge.scala 25:{25,25}]
  wire [31:0] _GEN_125 = 3'h5 == io_IDex[2:0] ? io_PreMat_5_7 : _GEN_124; // @[FinalMerge.scala 25:{25,25}]
  wire [31:0] _GEN_126 = 3'h6 == io_IDex[2:0] ? io_PreMat_6_7 : _GEN_125; // @[FinalMerge.scala 25:{25,25}]
  wire [31:0] _GEN_127 = 3'h7 == io_IDex[2:0] ? io_PreMat_7_7 : _GEN_126; // @[FinalMerge.scala 25:{25,25}]
  wire [31:0] _GEN_112 = 3'h0 == io_IDex[2:0] ? _GEN_127 : mat_0_7; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_113 = 3'h1 == io_IDex[2:0] ? _GEN_127 : mat_1_7; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_114 = 3'h2 == io_IDex[2:0] ? _GEN_127 : mat_2_7; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_115 = 3'h3 == io_IDex[2:0] ? _GEN_127 : mat_3_7; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_116 = 3'h4 == io_IDex[2:0] ? _GEN_127 : mat_4_7; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_117 = 3'h5 == io_IDex[2:0] ? _GEN_127 : mat_5_7; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_118 = 3'h6 == io_IDex[2:0] ? _GEN_127 : mat_6_7; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _GEN_119 = 3'h7 == io_IDex[2:0] ? _GEN_127 : mat_7_7; // @[FinalMerge.scala 16:22 25:{25,25}]
  wire [31:0] _i_T_1 = io_IDex + 32'h1; // @[FinalMerge.scala 30:16]
  wire  _GEN_403 = 3'h0 == i[2:0]; // @[FinalMerge.scala 33:{31,31}]
  wire  _GEN_404 = 3'h1 == j[2:0]; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_129 = 3'h0 == i[2:0] & 3'h1 == j[2:0] ? io_lastMat_0_1 : io_lastMat_0_0; // @[FinalMerge.scala 33:{31,31}]
  wire  _GEN_406 = 3'h2 == j[2:0]; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_130 = 3'h0 == i[2:0] & 3'h2 == j[2:0] ? io_lastMat_0_2 : _GEN_129; // @[FinalMerge.scala 33:{31,31}]
  wire  _GEN_408 = 3'h3 == j[2:0]; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_131 = 3'h0 == i[2:0] & 3'h3 == j[2:0] ? io_lastMat_0_3 : _GEN_130; // @[FinalMerge.scala 33:{31,31}]
  wire  _GEN_410 = 3'h4 == j[2:0]; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_132 = 3'h0 == i[2:0] & 3'h4 == j[2:0] ? io_lastMat_0_4 : _GEN_131; // @[FinalMerge.scala 33:{31,31}]
  wire  _GEN_412 = 3'h5 == j[2:0]; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_133 = 3'h0 == i[2:0] & 3'h5 == j[2:0] ? io_lastMat_0_5 : _GEN_132; // @[FinalMerge.scala 33:{31,31}]
  wire  _GEN_414 = 3'h6 == j[2:0]; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_134 = 3'h0 == i[2:0] & 3'h6 == j[2:0] ? io_lastMat_0_6 : _GEN_133; // @[FinalMerge.scala 33:{31,31}]
  wire  _GEN_416 = 3'h7 == j[2:0]; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_135 = 3'h0 == i[2:0] & 3'h7 == j[2:0] ? io_lastMat_0_7 : _GEN_134; // @[FinalMerge.scala 33:{31,31}]
  wire  _GEN_417 = 3'h1 == i[2:0]; // @[FinalMerge.scala 33:{31,31}]
  wire  _GEN_418 = 3'h0 == j[2:0]; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_136 = 3'h1 == i[2:0] & 3'h0 == j[2:0] ? io_lastMat_1_0 : _GEN_135; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_137 = 3'h1 == i[2:0] & 3'h1 == j[2:0] ? io_lastMat_1_1 : _GEN_136; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_138 = 3'h1 == i[2:0] & 3'h2 == j[2:0] ? io_lastMat_1_2 : _GEN_137; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_139 = 3'h1 == i[2:0] & 3'h3 == j[2:0] ? io_lastMat_1_3 : _GEN_138; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_140 = 3'h1 == i[2:0] & 3'h4 == j[2:0] ? io_lastMat_1_4 : _GEN_139; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_141 = 3'h1 == i[2:0] & 3'h5 == j[2:0] ? io_lastMat_1_5 : _GEN_140; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_142 = 3'h1 == i[2:0] & 3'h6 == j[2:0] ? io_lastMat_1_6 : _GEN_141; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_143 = 3'h1 == i[2:0] & 3'h7 == j[2:0] ? io_lastMat_1_7 : _GEN_142; // @[FinalMerge.scala 33:{31,31}]
  wire  _GEN_433 = 3'h2 == i[2:0]; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_144 = 3'h2 == i[2:0] & 3'h0 == j[2:0] ? io_lastMat_2_0 : _GEN_143; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_145 = 3'h2 == i[2:0] & 3'h1 == j[2:0] ? io_lastMat_2_1 : _GEN_144; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_146 = 3'h2 == i[2:0] & 3'h2 == j[2:0] ? io_lastMat_2_2 : _GEN_145; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_147 = 3'h2 == i[2:0] & 3'h3 == j[2:0] ? io_lastMat_2_3 : _GEN_146; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_148 = 3'h2 == i[2:0] & 3'h4 == j[2:0] ? io_lastMat_2_4 : _GEN_147; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_149 = 3'h2 == i[2:0] & 3'h5 == j[2:0] ? io_lastMat_2_5 : _GEN_148; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_150 = 3'h2 == i[2:0] & 3'h6 == j[2:0] ? io_lastMat_2_6 : _GEN_149; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_151 = 3'h2 == i[2:0] & 3'h7 == j[2:0] ? io_lastMat_2_7 : _GEN_150; // @[FinalMerge.scala 33:{31,31}]
  wire  _GEN_449 = 3'h3 == i[2:0]; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_152 = 3'h3 == i[2:0] & 3'h0 == j[2:0] ? io_lastMat_3_0 : _GEN_151; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_153 = 3'h3 == i[2:0] & 3'h1 == j[2:0] ? io_lastMat_3_1 : _GEN_152; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_154 = 3'h3 == i[2:0] & 3'h2 == j[2:0] ? io_lastMat_3_2 : _GEN_153; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_155 = 3'h3 == i[2:0] & 3'h3 == j[2:0] ? io_lastMat_3_3 : _GEN_154; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_156 = 3'h3 == i[2:0] & 3'h4 == j[2:0] ? io_lastMat_3_4 : _GEN_155; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_157 = 3'h3 == i[2:0] & 3'h5 == j[2:0] ? io_lastMat_3_5 : _GEN_156; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_158 = 3'h3 == i[2:0] & 3'h6 == j[2:0] ? io_lastMat_3_6 : _GEN_157; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_159 = 3'h3 == i[2:0] & 3'h7 == j[2:0] ? io_lastMat_3_7 : _GEN_158; // @[FinalMerge.scala 33:{31,31}]
  wire  _GEN_465 = 3'h4 == i[2:0]; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_160 = 3'h4 == i[2:0] & 3'h0 == j[2:0] ? io_lastMat_4_0 : _GEN_159; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_161 = 3'h4 == i[2:0] & 3'h1 == j[2:0] ? io_lastMat_4_1 : _GEN_160; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_162 = 3'h4 == i[2:0] & 3'h2 == j[2:0] ? io_lastMat_4_2 : _GEN_161; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_163 = 3'h4 == i[2:0] & 3'h3 == j[2:0] ? io_lastMat_4_3 : _GEN_162; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_164 = 3'h4 == i[2:0] & 3'h4 == j[2:0] ? io_lastMat_4_4 : _GEN_163; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_165 = 3'h4 == i[2:0] & 3'h5 == j[2:0] ? io_lastMat_4_5 : _GEN_164; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_166 = 3'h4 == i[2:0] & 3'h6 == j[2:0] ? io_lastMat_4_6 : _GEN_165; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_167 = 3'h4 == i[2:0] & 3'h7 == j[2:0] ? io_lastMat_4_7 : _GEN_166; // @[FinalMerge.scala 33:{31,31}]
  wire  _GEN_481 = 3'h5 == i[2:0]; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_168 = 3'h5 == i[2:0] & 3'h0 == j[2:0] ? io_lastMat_5_0 : _GEN_167; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_169 = 3'h5 == i[2:0] & 3'h1 == j[2:0] ? io_lastMat_5_1 : _GEN_168; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_170 = 3'h5 == i[2:0] & 3'h2 == j[2:0] ? io_lastMat_5_2 : _GEN_169; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_171 = 3'h5 == i[2:0] & 3'h3 == j[2:0] ? io_lastMat_5_3 : _GEN_170; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_172 = 3'h5 == i[2:0] & 3'h4 == j[2:0] ? io_lastMat_5_4 : _GEN_171; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_173 = 3'h5 == i[2:0] & 3'h5 == j[2:0] ? io_lastMat_5_5 : _GEN_172; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_174 = 3'h5 == i[2:0] & 3'h6 == j[2:0] ? io_lastMat_5_6 : _GEN_173; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_175 = 3'h5 == i[2:0] & 3'h7 == j[2:0] ? io_lastMat_5_7 : _GEN_174; // @[FinalMerge.scala 33:{31,31}]
  wire  _GEN_497 = 3'h6 == i[2:0]; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_176 = 3'h6 == i[2:0] & 3'h0 == j[2:0] ? io_lastMat_6_0 : _GEN_175; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_177 = 3'h6 == i[2:0] & 3'h1 == j[2:0] ? io_lastMat_6_1 : _GEN_176; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_178 = 3'h6 == i[2:0] & 3'h2 == j[2:0] ? io_lastMat_6_2 : _GEN_177; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_179 = 3'h6 == i[2:0] & 3'h3 == j[2:0] ? io_lastMat_6_3 : _GEN_178; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_180 = 3'h6 == i[2:0] & 3'h4 == j[2:0] ? io_lastMat_6_4 : _GEN_179; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_181 = 3'h6 == i[2:0] & 3'h5 == j[2:0] ? io_lastMat_6_5 : _GEN_180; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_182 = 3'h6 == i[2:0] & 3'h6 == j[2:0] ? io_lastMat_6_6 : _GEN_181; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_183 = 3'h6 == i[2:0] & 3'h7 == j[2:0] ? io_lastMat_6_7 : _GEN_182; // @[FinalMerge.scala 33:{31,31}]
  wire  _GEN_513 = 3'h7 == i[2:0]; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_184 = 3'h7 == i[2:0] & 3'h0 == j[2:0] ? io_lastMat_7_0 : _GEN_183; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_185 = 3'h7 == i[2:0] & 3'h1 == j[2:0] ? io_lastMat_7_1 : _GEN_184; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_186 = 3'h7 == i[2:0] & 3'h2 == j[2:0] ? io_lastMat_7_2 : _GEN_185; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_187 = 3'h7 == i[2:0] & 3'h3 == j[2:0] ? io_lastMat_7_3 : _GEN_186; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_188 = 3'h7 == i[2:0] & 3'h4 == j[2:0] ? io_lastMat_7_4 : _GEN_187; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_189 = 3'h7 == i[2:0] & 3'h5 == j[2:0] ? io_lastMat_7_5 : _GEN_188; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_190 = 3'h7 == i[2:0] & 3'h6 == j[2:0] ? io_lastMat_7_6 : _GEN_189; // @[FinalMerge.scala 33:{31,31}]
  wire [31:0] _GEN_191 = 3'h7 == i[2:0] & 3'h7 == j[2:0] ? io_lastMat_7_7 : _GEN_190; // @[FinalMerge.scala 33:{31,31}]
  wire  _T_14 = i < 32'h7; // @[FinalMerge.scala 38:16]
  wire  _T_15 = j == 32'h7; // @[FinalMerge.scala 38:46]
  wire [31:0] _i_T_3 = i + 32'h1; // @[FinalMerge.scala 39:14]
  wire  _T_17 = i == 32'h7; // @[FinalMerge.scala 42:17]
  wire  _T_18 = j < 32'h7; // @[FinalMerge.scala 42:51]
  wire [31:0] _j_T_1 = j + 32'h1; // @[FinalMerge.scala 45:12]
  wire  _T_22 = _T_17 & _T_15; // @[FinalMerge.scala 47:45]
  wire [31:0] _GEN_192 = _T_14 & _T_18 ? _j_T_1 : j; // @[FinalMerge.scala 21:20 52:74 53:9]
  wire [31:0] _GEN_195 = _T_17 & _T_15 ? j : _GEN_192; // @[FinalMerge.scala 47:80 51:9]
  wire [31:0] _GEN_197 = i == 32'h7 & j < 32'h7 ? _j_T_1 : _GEN_195; // @[FinalMerge.scala 42:77 45:7]
  wire  _GEN_198 = i == 32'h7 & j < 32'h7 ? 1'h0 : _T_22; // @[FinalMerge.scala 18:15 42:77]
  wire [31:0] _GEN_199 = i < 32'h7 & j == 32'h7 ? _i_T_3 : i; // @[FinalMerge.scala 38:74 39:9]
  wire [31:0] _GEN_200 = i < 32'h7 & j == 32'h7 ? 32'h0 : _GEN_197; // @[FinalMerge.scala 38:74 40:9]
  wire  _GEN_201 = i < 32'h7 & j == 32'h7 ? 1'h0 : _GEN_198; // @[FinalMerge.scala 18:15 38:74]
  wire  _GEN_204 = _GEN_191 == 32'h4 | _GEN_201; // @[FinalMerge.scala 33:40 36:17]
  wire  _GEN_207 = i == 32'h0 & j == 32'h0 ? 1'h0 : _GEN_204; // @[FinalMerge.scala 18:15 29:37]
  assign io_Ovalid = io_valid & _GEN_207; // @[FinalMerge.scala 18:15 28:16]
  assign io_omat_0_0 = mat_0_0; // @[FinalMerge.scala 17:13]
  assign io_omat_0_1 = mat_0_1; // @[FinalMerge.scala 17:13]
  assign io_omat_0_2 = mat_0_2; // @[FinalMerge.scala 17:13]
  assign io_omat_0_3 = mat_0_3; // @[FinalMerge.scala 17:13]
  assign io_omat_0_4 = mat_0_4; // @[FinalMerge.scala 17:13]
  assign io_omat_0_5 = mat_0_5; // @[FinalMerge.scala 17:13]
  assign io_omat_0_6 = mat_0_6; // @[FinalMerge.scala 17:13]
  assign io_omat_0_7 = mat_0_7; // @[FinalMerge.scala 17:13]
  assign io_omat_1_0 = mat_1_0; // @[FinalMerge.scala 17:13]
  assign io_omat_1_1 = mat_1_1; // @[FinalMerge.scala 17:13]
  assign io_omat_1_2 = mat_1_2; // @[FinalMerge.scala 17:13]
  assign io_omat_1_3 = mat_1_3; // @[FinalMerge.scala 17:13]
  assign io_omat_1_4 = mat_1_4; // @[FinalMerge.scala 17:13]
  assign io_omat_1_5 = mat_1_5; // @[FinalMerge.scala 17:13]
  assign io_omat_1_6 = mat_1_6; // @[FinalMerge.scala 17:13]
  assign io_omat_1_7 = mat_1_7; // @[FinalMerge.scala 17:13]
  assign io_omat_2_0 = mat_2_0; // @[FinalMerge.scala 17:13]
  assign io_omat_2_1 = mat_2_1; // @[FinalMerge.scala 17:13]
  assign io_omat_2_2 = mat_2_2; // @[FinalMerge.scala 17:13]
  assign io_omat_2_3 = mat_2_3; // @[FinalMerge.scala 17:13]
  assign io_omat_2_4 = mat_2_4; // @[FinalMerge.scala 17:13]
  assign io_omat_2_5 = mat_2_5; // @[FinalMerge.scala 17:13]
  assign io_omat_2_6 = mat_2_6; // @[FinalMerge.scala 17:13]
  assign io_omat_2_7 = mat_2_7; // @[FinalMerge.scala 17:13]
  assign io_omat_3_0 = mat_3_0; // @[FinalMerge.scala 17:13]
  assign io_omat_3_1 = mat_3_1; // @[FinalMerge.scala 17:13]
  assign io_omat_3_2 = mat_3_2; // @[FinalMerge.scala 17:13]
  assign io_omat_3_3 = mat_3_3; // @[FinalMerge.scala 17:13]
  assign io_omat_3_4 = mat_3_4; // @[FinalMerge.scala 17:13]
  assign io_omat_3_5 = mat_3_5; // @[FinalMerge.scala 17:13]
  assign io_omat_3_6 = mat_3_6; // @[FinalMerge.scala 17:13]
  assign io_omat_3_7 = mat_3_7; // @[FinalMerge.scala 17:13]
  assign io_omat_4_0 = mat_4_0; // @[FinalMerge.scala 17:13]
  assign io_omat_4_1 = mat_4_1; // @[FinalMerge.scala 17:13]
  assign io_omat_4_2 = mat_4_2; // @[FinalMerge.scala 17:13]
  assign io_omat_4_3 = mat_4_3; // @[FinalMerge.scala 17:13]
  assign io_omat_4_4 = mat_4_4; // @[FinalMerge.scala 17:13]
  assign io_omat_4_5 = mat_4_5; // @[FinalMerge.scala 17:13]
  assign io_omat_4_6 = mat_4_6; // @[FinalMerge.scala 17:13]
  assign io_omat_4_7 = mat_4_7; // @[FinalMerge.scala 17:13]
  assign io_omat_5_0 = mat_5_0; // @[FinalMerge.scala 17:13]
  assign io_omat_5_1 = mat_5_1; // @[FinalMerge.scala 17:13]
  assign io_omat_5_2 = mat_5_2; // @[FinalMerge.scala 17:13]
  assign io_omat_5_3 = mat_5_3; // @[FinalMerge.scala 17:13]
  assign io_omat_5_4 = mat_5_4; // @[FinalMerge.scala 17:13]
  assign io_omat_5_5 = mat_5_5; // @[FinalMerge.scala 17:13]
  assign io_omat_5_6 = mat_5_6; // @[FinalMerge.scala 17:13]
  assign io_omat_5_7 = mat_5_7; // @[FinalMerge.scala 17:13]
  assign io_omat_6_0 = mat_6_0; // @[FinalMerge.scala 17:13]
  assign io_omat_6_1 = mat_6_1; // @[FinalMerge.scala 17:13]
  assign io_omat_6_2 = mat_6_2; // @[FinalMerge.scala 17:13]
  assign io_omat_6_3 = mat_6_3; // @[FinalMerge.scala 17:13]
  assign io_omat_6_4 = mat_6_4; // @[FinalMerge.scala 17:13]
  assign io_omat_6_5 = mat_6_5; // @[FinalMerge.scala 17:13]
  assign io_omat_6_6 = mat_6_6; // @[FinalMerge.scala 17:13]
  assign io_omat_6_7 = mat_6_7; // @[FinalMerge.scala 17:13]
  assign io_omat_7_0 = mat_7_0; // @[FinalMerge.scala 17:13]
  assign io_omat_7_1 = mat_7_1; // @[FinalMerge.scala 17:13]
  assign io_omat_7_2 = mat_7_2; // @[FinalMerge.scala 17:13]
  assign io_omat_7_3 = mat_7_3; // @[FinalMerge.scala 17:13]
  assign io_omat_7_4 = mat_7_4; // @[FinalMerge.scala 17:13]
  assign io_omat_7_5 = mat_7_5; // @[FinalMerge.scala 17:13]
  assign io_omat_7_6 = mat_7_6; // @[FinalMerge.scala 17:13]
  assign io_omat_7_7 = mat_7_7; // @[FinalMerge.scala 17:13]
  always @(posedge clock) begin
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_0_0 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_403 & _GEN_418) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_0_0 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_0_0 <= _GEN_190;
        end
      end else begin
        mat_0_0 <= _GEN_0;
      end
    end else begin
      mat_0_0 <= _GEN_0;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_0_1 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_403 & _GEN_404) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_0_1 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_0_1 <= _GEN_190;
        end
      end else begin
        mat_0_1 <= _GEN_16;
      end
    end else begin
      mat_0_1 <= _GEN_16;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_0_2 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_403 & _GEN_406) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_0_2 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_0_2 <= _GEN_190;
        end
      end else begin
        mat_0_2 <= _GEN_32;
      end
    end else begin
      mat_0_2 <= _GEN_32;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_0_3 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_403 & _GEN_408) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_0_3 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_0_3 <= _GEN_190;
        end
      end else begin
        mat_0_3 <= _GEN_48;
      end
    end else begin
      mat_0_3 <= _GEN_48;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_0_4 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_403 & _GEN_410) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_0_4 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_0_4 <= _GEN_190;
        end
      end else begin
        mat_0_4 <= _GEN_64;
      end
    end else begin
      mat_0_4 <= _GEN_64;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_0_5 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_403 & _GEN_412) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_0_5 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_0_5 <= _GEN_190;
        end
      end else begin
        mat_0_5 <= _GEN_80;
      end
    end else begin
      mat_0_5 <= _GEN_80;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_0_6 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_403 & _GEN_414) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_0_6 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_0_6 <= _GEN_190;
        end
      end else begin
        mat_0_6 <= _GEN_96;
      end
    end else begin
      mat_0_6 <= _GEN_96;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_0_7 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_403 & _GEN_416) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_0_7 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_0_7 <= _GEN_190;
        end
      end else begin
        mat_0_7 <= _GEN_112;
      end
    end else begin
      mat_0_7 <= _GEN_112;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_1_0 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_417 & _GEN_418) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_1_0 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_1_0 <= _GEN_190;
        end
      end else begin
        mat_1_0 <= _GEN_1;
      end
    end else begin
      mat_1_0 <= _GEN_1;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_1_1 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_417 & _GEN_404) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_1_1 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_1_1 <= _GEN_190;
        end
      end else begin
        mat_1_1 <= _GEN_17;
      end
    end else begin
      mat_1_1 <= _GEN_17;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_1_2 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_417 & _GEN_406) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_1_2 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_1_2 <= _GEN_190;
        end
      end else begin
        mat_1_2 <= _GEN_33;
      end
    end else begin
      mat_1_2 <= _GEN_33;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_1_3 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_417 & _GEN_408) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_1_3 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_1_3 <= _GEN_190;
        end
      end else begin
        mat_1_3 <= _GEN_49;
      end
    end else begin
      mat_1_3 <= _GEN_49;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_1_4 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_417 & _GEN_410) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_1_4 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_1_4 <= _GEN_190;
        end
      end else begin
        mat_1_4 <= _GEN_65;
      end
    end else begin
      mat_1_4 <= _GEN_65;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_1_5 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_417 & _GEN_412) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_1_5 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_1_5 <= _GEN_190;
        end
      end else begin
        mat_1_5 <= _GEN_81;
      end
    end else begin
      mat_1_5 <= _GEN_81;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_1_6 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_417 & _GEN_414) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_1_6 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_1_6 <= _GEN_190;
        end
      end else begin
        mat_1_6 <= _GEN_97;
      end
    end else begin
      mat_1_6 <= _GEN_97;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_1_7 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_417 & _GEN_416) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_1_7 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_1_7 <= _GEN_190;
        end
      end else begin
        mat_1_7 <= _GEN_113;
      end
    end else begin
      mat_1_7 <= _GEN_113;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_2_0 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_433 & _GEN_418) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_2_0 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_2_0 <= _GEN_190;
        end
      end else begin
        mat_2_0 <= _GEN_2;
      end
    end else begin
      mat_2_0 <= _GEN_2;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_2_1 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_433 & _GEN_404) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_2_1 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_2_1 <= _GEN_190;
        end
      end else begin
        mat_2_1 <= _GEN_18;
      end
    end else begin
      mat_2_1 <= _GEN_18;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_2_2 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_433 & _GEN_406) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_2_2 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_2_2 <= _GEN_190;
        end
      end else begin
        mat_2_2 <= _GEN_34;
      end
    end else begin
      mat_2_2 <= _GEN_34;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_2_3 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_433 & _GEN_408) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_2_3 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_2_3 <= _GEN_190;
        end
      end else begin
        mat_2_3 <= _GEN_50;
      end
    end else begin
      mat_2_3 <= _GEN_50;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_2_4 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_433 & _GEN_410) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_2_4 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_2_4 <= _GEN_190;
        end
      end else begin
        mat_2_4 <= _GEN_66;
      end
    end else begin
      mat_2_4 <= _GEN_66;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_2_5 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_433 & _GEN_412) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_2_5 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_2_5 <= _GEN_190;
        end
      end else begin
        mat_2_5 <= _GEN_82;
      end
    end else begin
      mat_2_5 <= _GEN_82;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_2_6 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_433 & _GEN_414) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_2_6 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_2_6 <= _GEN_190;
        end
      end else begin
        mat_2_6 <= _GEN_98;
      end
    end else begin
      mat_2_6 <= _GEN_98;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_2_7 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_433 & _GEN_416) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_2_7 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_2_7 <= _GEN_190;
        end
      end else begin
        mat_2_7 <= _GEN_114;
      end
    end else begin
      mat_2_7 <= _GEN_114;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_3_0 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_449 & _GEN_418) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_3_0 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_3_0 <= _GEN_190;
        end
      end else begin
        mat_3_0 <= _GEN_3;
      end
    end else begin
      mat_3_0 <= _GEN_3;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_3_1 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_449 & _GEN_404) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_3_1 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_3_1 <= _GEN_190;
        end
      end else begin
        mat_3_1 <= _GEN_19;
      end
    end else begin
      mat_3_1 <= _GEN_19;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_3_2 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_449 & _GEN_406) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_3_2 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_3_2 <= _GEN_190;
        end
      end else begin
        mat_3_2 <= _GEN_35;
      end
    end else begin
      mat_3_2 <= _GEN_35;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_3_3 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_449 & _GEN_408) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_3_3 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_3_3 <= _GEN_190;
        end
      end else begin
        mat_3_3 <= _GEN_51;
      end
    end else begin
      mat_3_3 <= _GEN_51;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_3_4 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_449 & _GEN_410) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_3_4 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_3_4 <= _GEN_190;
        end
      end else begin
        mat_3_4 <= _GEN_67;
      end
    end else begin
      mat_3_4 <= _GEN_67;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_3_5 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_449 & _GEN_412) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_3_5 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_3_5 <= _GEN_190;
        end
      end else begin
        mat_3_5 <= _GEN_83;
      end
    end else begin
      mat_3_5 <= _GEN_83;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_3_6 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_449 & _GEN_414) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_3_6 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_3_6 <= _GEN_190;
        end
      end else begin
        mat_3_6 <= _GEN_99;
      end
    end else begin
      mat_3_6 <= _GEN_99;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_3_7 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_449 & _GEN_416) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_3_7 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_3_7 <= _GEN_190;
        end
      end else begin
        mat_3_7 <= _GEN_115;
      end
    end else begin
      mat_3_7 <= _GEN_115;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_4_0 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_465 & _GEN_418) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_4_0 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_4_0 <= _GEN_190;
        end
      end else begin
        mat_4_0 <= _GEN_4;
      end
    end else begin
      mat_4_0 <= _GEN_4;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_4_1 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_465 & _GEN_404) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_4_1 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_4_1 <= _GEN_190;
        end
      end else begin
        mat_4_1 <= _GEN_20;
      end
    end else begin
      mat_4_1 <= _GEN_20;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_4_2 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_465 & _GEN_406) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_4_2 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_4_2 <= _GEN_190;
        end
      end else begin
        mat_4_2 <= _GEN_36;
      end
    end else begin
      mat_4_2 <= _GEN_36;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_4_3 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_465 & _GEN_408) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_4_3 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_4_3 <= _GEN_190;
        end
      end else begin
        mat_4_3 <= _GEN_52;
      end
    end else begin
      mat_4_3 <= _GEN_52;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_4_4 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_465 & _GEN_410) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_4_4 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_4_4 <= _GEN_190;
        end
      end else begin
        mat_4_4 <= _GEN_68;
      end
    end else begin
      mat_4_4 <= _GEN_68;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_4_5 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_465 & _GEN_412) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_4_5 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_4_5 <= _GEN_190;
        end
      end else begin
        mat_4_5 <= _GEN_84;
      end
    end else begin
      mat_4_5 <= _GEN_84;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_4_6 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_465 & _GEN_414) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_4_6 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_4_6 <= _GEN_190;
        end
      end else begin
        mat_4_6 <= _GEN_100;
      end
    end else begin
      mat_4_6 <= _GEN_100;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_4_7 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_465 & _GEN_416) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_4_7 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_4_7 <= _GEN_190;
        end
      end else begin
        mat_4_7 <= _GEN_116;
      end
    end else begin
      mat_4_7 <= _GEN_116;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_5_0 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_481 & _GEN_418) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_5_0 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_5_0 <= _GEN_190;
        end
      end else begin
        mat_5_0 <= _GEN_5;
      end
    end else begin
      mat_5_0 <= _GEN_5;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_5_1 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_481 & _GEN_404) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_5_1 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_5_1 <= _GEN_190;
        end
      end else begin
        mat_5_1 <= _GEN_21;
      end
    end else begin
      mat_5_1 <= _GEN_21;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_5_2 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_481 & _GEN_406) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_5_2 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_5_2 <= _GEN_190;
        end
      end else begin
        mat_5_2 <= _GEN_37;
      end
    end else begin
      mat_5_2 <= _GEN_37;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_5_3 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_481 & _GEN_408) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_5_3 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_5_3 <= _GEN_190;
        end
      end else begin
        mat_5_3 <= _GEN_53;
      end
    end else begin
      mat_5_3 <= _GEN_53;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_5_4 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_481 & _GEN_410) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_5_4 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_5_4 <= _GEN_190;
        end
      end else begin
        mat_5_4 <= _GEN_69;
      end
    end else begin
      mat_5_4 <= _GEN_69;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_5_5 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_481 & _GEN_412) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_5_5 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_5_5 <= _GEN_190;
        end
      end else begin
        mat_5_5 <= _GEN_85;
      end
    end else begin
      mat_5_5 <= _GEN_85;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_5_6 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_481 & _GEN_414) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_5_6 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_5_6 <= _GEN_190;
        end
      end else begin
        mat_5_6 <= _GEN_101;
      end
    end else begin
      mat_5_6 <= _GEN_101;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_5_7 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_481 & _GEN_416) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_5_7 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_5_7 <= _GEN_190;
        end
      end else begin
        mat_5_7 <= _GEN_117;
      end
    end else begin
      mat_5_7 <= _GEN_117;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_6_0 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_497 & _GEN_418) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_6_0 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_6_0 <= _GEN_190;
        end
      end else begin
        mat_6_0 <= _GEN_6;
      end
    end else begin
      mat_6_0 <= _GEN_6;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_6_1 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_497 & _GEN_404) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_6_1 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_6_1 <= _GEN_190;
        end
      end else begin
        mat_6_1 <= _GEN_22;
      end
    end else begin
      mat_6_1 <= _GEN_22;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_6_2 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_497 & _GEN_406) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_6_2 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_6_2 <= _GEN_190;
        end
      end else begin
        mat_6_2 <= _GEN_38;
      end
    end else begin
      mat_6_2 <= _GEN_38;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_6_3 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_497 & _GEN_408) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_6_3 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_6_3 <= _GEN_190;
        end
      end else begin
        mat_6_3 <= _GEN_54;
      end
    end else begin
      mat_6_3 <= _GEN_54;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_6_4 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_497 & _GEN_410) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_6_4 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_6_4 <= _GEN_190;
        end
      end else begin
        mat_6_4 <= _GEN_70;
      end
    end else begin
      mat_6_4 <= _GEN_70;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_6_5 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_497 & _GEN_412) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_6_5 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_6_5 <= _GEN_190;
        end
      end else begin
        mat_6_5 <= _GEN_86;
      end
    end else begin
      mat_6_5 <= _GEN_86;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_6_6 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_497 & _GEN_414) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_6_6 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_6_6 <= _GEN_190;
        end
      end else begin
        mat_6_6 <= _GEN_102;
      end
    end else begin
      mat_6_6 <= _GEN_102;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_6_7 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_497 & _GEN_416) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_6_7 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_6_7 <= _GEN_190;
        end
      end else begin
        mat_6_7 <= _GEN_118;
      end
    end else begin
      mat_6_7 <= _GEN_118;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_7_0 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_513 & _GEN_418) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_7_0 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_7_0 <= _GEN_190;
        end
      end else begin
        mat_7_0 <= _GEN_7;
      end
    end else begin
      mat_7_0 <= _GEN_7;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_7_1 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_513 & _GEN_404) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_7_1 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_7_1 <= _GEN_190;
        end
      end else begin
        mat_7_1 <= _GEN_23;
      end
    end else begin
      mat_7_1 <= _GEN_23;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_7_2 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_513 & _GEN_406) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_7_2 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_7_2 <= _GEN_190;
        end
      end else begin
        mat_7_2 <= _GEN_39;
      end
    end else begin
      mat_7_2 <= _GEN_39;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_7_3 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_513 & _GEN_408) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_7_3 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_7_3 <= _GEN_190;
        end
      end else begin
        mat_7_3 <= _GEN_55;
      end
    end else begin
      mat_7_3 <= _GEN_55;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_7_4 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_513 & _GEN_410) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_7_4 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_7_4 <= _GEN_190;
        end
      end else begin
        mat_7_4 <= _GEN_71;
      end
    end else begin
      mat_7_4 <= _GEN_71;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_7_5 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_513 & _GEN_412) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_7_5 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_7_5 <= _GEN_190;
        end
      end else begin
        mat_7_5 <= _GEN_87;
      end
    end else begin
      mat_7_5 <= _GEN_87;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_7_6 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_513 & _GEN_414) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_7_6 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_7_6 <= _GEN_190;
        end
      end else begin
        mat_7_6 <= _GEN_103;
      end
    end else begin
      mat_7_6 <= _GEN_103;
    end
    if (reset) begin // @[FinalMerge.scala 16:22]
      mat_7_7 <= 32'h0; // @[FinalMerge.scala 16:22]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (_GEN_513 & _GEN_416) begin // @[FinalMerge.scala 56:15]
        if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[FinalMerge.scala 33:31]
          mat_7_7 <= io_lastMat_7_7; // @[FinalMerge.scala 33:31]
        end else begin
          mat_7_7 <= _GEN_190;
        end
      end else begin
        mat_7_7 <= _GEN_119;
      end
    end else begin
      mat_7_7 <= _GEN_119;
    end
    if (reset) begin // @[FinalMerge.scala 20:20]
      i <= 32'h0; // @[FinalMerge.scala 20:20]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (i == 32'h0 & j == 32'h0) begin // @[FinalMerge.scala 29:37]
        i <= _i_T_1; // @[FinalMerge.scala 30:5]
      end else if (!(_GEN_191 == 32'h4)) begin // @[FinalMerge.scala 33:40]
        i <= _GEN_199;
      end
    end
    if (reset) begin // @[FinalMerge.scala 21:20]
      j <= 32'h0; // @[FinalMerge.scala 21:20]
    end else if (io_valid) begin // @[FinalMerge.scala 28:16]
      if (i == 32'h0 & j == 32'h0) begin // @[FinalMerge.scala 29:37]
        j <= 32'h0; // @[FinalMerge.scala 31:7]
      end else if (!(_GEN_191 == 32'h4)) begin // @[FinalMerge.scala 33:40]
        j <= _GEN_200;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  mat_0_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  mat_0_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  mat_0_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  mat_0_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  mat_0_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  mat_0_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  mat_0_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  mat_0_7 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  mat_1_0 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  mat_1_1 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  mat_1_2 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  mat_1_3 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  mat_1_4 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  mat_1_5 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  mat_1_6 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  mat_1_7 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  mat_2_0 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  mat_2_1 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  mat_2_2 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  mat_2_3 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  mat_2_4 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  mat_2_5 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  mat_2_6 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  mat_2_7 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  mat_3_0 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  mat_3_1 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  mat_3_2 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  mat_3_3 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  mat_3_4 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  mat_3_5 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  mat_3_6 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  mat_3_7 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  mat_4_0 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  mat_4_1 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  mat_4_2 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  mat_4_3 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  mat_4_4 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  mat_4_5 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  mat_4_6 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  mat_4_7 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  mat_5_0 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  mat_5_1 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  mat_5_2 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  mat_5_3 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  mat_5_4 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  mat_5_5 = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  mat_5_6 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  mat_5_7 = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  mat_6_0 = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  mat_6_1 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  mat_6_2 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  mat_6_3 = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  mat_6_4 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  mat_6_5 = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  mat_6_6 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  mat_6_7 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  mat_7_0 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  mat_7_1 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  mat_7_2 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  mat_7_3 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  mat_7_4 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  mat_7_5 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  mat_7_6 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  mat_7_7 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  i = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  j = _RAND_65[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Distribution2(
  input         clock,
  input         reset,
  input  [31:0] io_matrix_0_0,
  input  [31:0] io_matrix_0_1,
  input  [31:0] io_matrix_0_2,
  input  [31:0] io_matrix_0_3,
  input  [31:0] io_matrix_0_4,
  input  [31:0] io_matrix_0_5,
  input  [31:0] io_matrix_0_6,
  input  [31:0] io_matrix_0_7,
  input  [31:0] io_matrix_1_0,
  input  [31:0] io_matrix_1_1,
  input  [31:0] io_matrix_1_2,
  input  [31:0] io_matrix_1_3,
  input  [31:0] io_matrix_1_4,
  input  [31:0] io_matrix_1_5,
  input  [31:0] io_matrix_1_6,
  input  [31:0] io_matrix_1_7,
  input  [31:0] io_matrix_2_0,
  input  [31:0] io_matrix_2_1,
  input  [31:0] io_matrix_2_2,
  input  [31:0] io_matrix_2_3,
  input  [31:0] io_matrix_2_4,
  input  [31:0] io_matrix_2_5,
  input  [31:0] io_matrix_2_6,
  input  [31:0] io_matrix_2_7,
  input  [31:0] io_matrix_3_0,
  input  [31:0] io_matrix_3_1,
  input  [31:0] io_matrix_3_2,
  input  [31:0] io_matrix_3_3,
  input  [31:0] io_matrix_3_4,
  input  [31:0] io_matrix_3_5,
  input  [31:0] io_matrix_3_6,
  input  [31:0] io_matrix_3_7,
  input  [31:0] io_matrix_4_0,
  input  [31:0] io_matrix_4_1,
  input  [31:0] io_matrix_4_2,
  input  [31:0] io_matrix_4_3,
  input  [31:0] io_matrix_4_4,
  input  [31:0] io_matrix_4_5,
  input  [31:0] io_matrix_4_6,
  input  [31:0] io_matrix_4_7,
  input  [31:0] io_matrix_5_0,
  input  [31:0] io_matrix_5_1,
  input  [31:0] io_matrix_5_2,
  input  [31:0] io_matrix_5_3,
  input  [31:0] io_matrix_5_4,
  input  [31:0] io_matrix_5_5,
  input  [31:0] io_matrix_5_6,
  input  [31:0] io_matrix_5_7,
  input  [31:0] io_matrix_6_0,
  input  [31:0] io_matrix_6_1,
  input  [31:0] io_matrix_6_2,
  input  [31:0] io_matrix_6_3,
  input  [31:0] io_matrix_6_4,
  input  [31:0] io_matrix_6_5,
  input  [31:0] io_matrix_6_6,
  input  [31:0] io_matrix_6_7,
  input  [31:0] io_matrix_7_0,
  input  [31:0] io_matrix_7_1,
  input  [31:0] io_matrix_7_2,
  input  [31:0] io_matrix_7_3,
  input  [31:0] io_matrix_7_4,
  input  [31:0] io_matrix_7_5,
  input  [31:0] io_matrix_7_6,
  input  [31:0] io_matrix_7_7,
  input  [31:0] io_s,
  output [31:0] io_out_0_0,
  output [31:0] io_out_0_1,
  output [31:0] io_out_0_2,
  output [31:0] io_out_0_3,
  output [31:0] io_out_0_4,
  output [31:0] io_out_0_5,
  output [31:0] io_out_0_6,
  output [31:0] io_out_0_7,
  output [31:0] io_out_1_0,
  output [31:0] io_out_1_1,
  output [31:0] io_out_1_2,
  output [31:0] io_out_1_3,
  output [31:0] io_out_1_4,
  output [31:0] io_out_1_5,
  output [31:0] io_out_1_6,
  output [31:0] io_out_1_7,
  output [31:0] io_out_2_0,
  output [31:0] io_out_2_1,
  output [31:0] io_out_2_2,
  output [31:0] io_out_2_3,
  output [31:0] io_out_2_4,
  output [31:0] io_out_2_5,
  output [31:0] io_out_2_6,
  output [31:0] io_out_2_7,
  output [31:0] io_out_3_0,
  output [31:0] io_out_3_1,
  output [31:0] io_out_3_2,
  output [31:0] io_out_3_3,
  output [31:0] io_out_3_4,
  output [31:0] io_out_3_5,
  output [31:0] io_out_3_6,
  output [31:0] io_out_3_7,
  output [31:0] io_out_4_0,
  output [31:0] io_out_4_1,
  output [31:0] io_out_4_2,
  output [31:0] io_out_4_3,
  output [31:0] io_out_4_4,
  output [31:0] io_out_4_5,
  output [31:0] io_out_4_6,
  output [31:0] io_out_4_7,
  output [31:0] io_out_5_0,
  output [31:0] io_out_5_1,
  output [31:0] io_out_5_2,
  output [31:0] io_out_5_3,
  output [31:0] io_out_5_4,
  output [31:0] io_out_5_5,
  output [31:0] io_out_5_6,
  output [31:0] io_out_5_7,
  output [31:0] io_out_6_0,
  output [31:0] io_out_6_1,
  output [31:0] io_out_6_2,
  output [31:0] io_out_6_3,
  output [31:0] io_out_6_4,
  output [31:0] io_out_6_5,
  output [31:0] io_out_6_6,
  output [31:0] io_out_6_7,
  output [31:0] io_out_7_0,
  output [31:0] io_out_7_1,
  output [31:0] io_out_7_2,
  output [31:0] io_out_7_3,
  output [31:0] io_out_7_4,
  output [31:0] io_out_7_5,
  output [31:0] io_out_7_6,
  output [31:0] io_out_7_7,
  output        io_ProcessValid,
  input         io_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
`endif // RANDOMIZE_REG_INIT
  wire  part2_clock; // @[Distribution2.scala 75:23]
  wire  part2_reset; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_IDex; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_JDex; // @[Distribution2.scala 75:23]
  wire  part2_io_valid; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_0_0; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_0_1; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_0_2; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_0_3; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_0_4; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_0_5; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_0_6; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_0_7; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_1_0; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_1_1; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_1_2; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_1_3; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_1_4; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_1_5; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_1_6; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_1_7; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_2_0; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_2_1; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_2_2; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_2_3; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_2_4; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_2_5; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_2_6; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_2_7; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_3_0; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_3_1; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_3_2; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_3_3; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_3_4; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_3_5; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_3_6; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_3_7; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_4_0; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_4_1; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_4_2; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_4_3; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_4_4; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_4_5; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_4_6; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_4_7; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_5_0; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_5_1; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_5_2; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_5_3; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_5_4; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_5_5; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_5_6; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_5_7; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_6_0; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_6_1; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_6_2; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_6_3; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_6_4; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_6_5; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_6_6; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_6_7; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_7_0; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_7_1; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_7_2; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_7_3; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_7_4; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_7_5; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_7_6; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_mat_7_7; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_0_0; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_0_1; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_0_2; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_0_3; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_0_4; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_0_5; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_0_6; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_0_7; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_1_0; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_1_1; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_1_2; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_1_3; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_1_4; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_1_5; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_1_6; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_1_7; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_2_0; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_2_1; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_2_2; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_2_3; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_2_4; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_2_5; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_2_6; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_2_7; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_3_0; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_3_1; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_3_2; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_3_3; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_3_4; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_3_5; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_3_6; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_3_7; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_4_0; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_4_1; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_4_2; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_4_3; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_4_4; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_4_5; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_4_6; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_4_7; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_5_0; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_5_1; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_5_2; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_5_3; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_5_4; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_5_5; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_5_6; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_5_7; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_6_0; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_6_1; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_6_2; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_6_3; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_6_4; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_6_5; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_6_6; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_6_7; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_7_0; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_7_1; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_7_2; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_7_3; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_7_4; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_7_5; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_7_6; // @[Distribution2.scala 75:23]
  wire [31:0] part2_io_OutMat_7_7; // @[Distribution2.scala 75:23]
  wire  part2_io_Ovalid; // @[Distribution2.scala 75:23]
  wire  part2_io_ProcessValid; // @[Distribution2.scala 75:23]
  wire  part3_clock; // @[Distribution2.scala 90:23]
  wire  part3_reset; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_IDex; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_0_0; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_0_1; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_0_2; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_0_3; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_0_4; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_0_5; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_0_6; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_0_7; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_1_0; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_1_1; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_1_2; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_1_3; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_1_4; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_1_5; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_1_6; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_1_7; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_2_0; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_2_1; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_2_2; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_2_3; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_2_4; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_2_5; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_2_6; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_2_7; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_3_0; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_3_1; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_3_2; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_3_3; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_3_4; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_3_5; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_3_6; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_3_7; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_4_0; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_4_1; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_4_2; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_4_3; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_4_4; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_4_5; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_4_6; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_4_7; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_5_0; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_5_1; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_5_2; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_5_3; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_5_4; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_5_5; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_5_6; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_5_7; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_6_0; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_6_1; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_6_2; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_6_3; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_6_4; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_6_5; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_6_6; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_6_7; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_7_0; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_7_1; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_7_2; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_7_3; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_7_4; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_7_5; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_7_6; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_mat_7_7; // @[Distribution2.scala 90:23]
  wire  part3_io_i_valid; // @[Distribution2.scala 90:23]
  wire  part3_io_valid; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_0_0; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_0_1; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_0_2; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_0_3; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_0_4; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_0_5; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_0_6; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_0_7; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_1_0; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_1_1; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_1_2; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_1_3; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_1_4; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_1_5; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_1_6; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_1_7; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_2_0; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_2_1; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_2_2; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_2_3; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_2_4; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_2_5; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_2_6; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_2_7; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_3_0; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_3_1; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_3_2; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_3_3; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_3_4; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_3_5; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_3_6; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_3_7; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_4_0; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_4_1; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_4_2; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_4_3; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_4_4; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_4_5; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_4_6; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_4_7; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_5_0; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_5_1; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_5_2; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_5_3; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_5_4; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_5_5; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_5_6; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_5_7; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_6_0; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_6_1; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_6_2; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_6_3; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_6_4; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_6_5; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_6_6; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_6_7; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_7_0; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_7_1; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_7_2; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_7_3; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_7_4; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_7_5; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_7_6; // @[Distribution2.scala 90:23]
  wire [31:0] part3_io_Omat_7_7; // @[Distribution2.scala 90:23]
  wire  Final_clock; // @[Distribution2.scala 114:31]
  wire  Final_reset; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_IDex; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_0_0; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_0_1; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_0_2; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_0_3; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_0_4; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_0_5; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_0_6; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_0_7; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_1_0; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_1_1; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_1_2; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_1_3; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_1_4; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_1_5; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_1_6; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_1_7; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_2_0; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_2_1; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_2_2; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_2_3; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_2_4; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_2_5; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_2_6; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_2_7; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_3_0; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_3_1; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_3_2; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_3_3; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_3_4; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_3_5; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_3_6; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_3_7; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_4_0; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_4_1; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_4_2; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_4_3; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_4_4; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_4_5; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_4_6; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_4_7; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_5_0; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_5_1; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_5_2; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_5_3; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_5_4; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_5_5; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_5_6; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_5_7; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_6_0; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_6_1; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_6_2; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_6_3; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_6_4; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_6_5; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_6_6; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_6_7; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_7_0; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_7_1; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_7_2; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_7_3; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_7_4; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_7_5; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_7_6; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_PreMat_7_7; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_0_0; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_0_1; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_0_2; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_0_3; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_0_4; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_0_5; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_0_6; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_0_7; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_1_0; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_1_1; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_1_2; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_1_3; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_1_4; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_1_5; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_1_6; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_1_7; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_2_0; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_2_1; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_2_2; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_2_3; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_2_4; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_2_5; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_2_6; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_2_7; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_3_0; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_3_1; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_3_2; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_3_3; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_3_4; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_3_5; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_3_6; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_3_7; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_4_0; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_4_1; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_4_2; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_4_3; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_4_4; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_4_5; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_4_6; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_4_7; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_5_0; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_5_1; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_5_2; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_5_3; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_5_4; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_5_5; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_5_6; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_5_7; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_6_0; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_6_1; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_6_2; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_6_3; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_6_4; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_6_5; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_6_6; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_6_7; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_7_0; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_7_1; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_7_2; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_7_3; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_7_4; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_7_5; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_7_6; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_lastMat_7_7; // @[Distribution2.scala 114:31]
  wire  Final_io_valid; // @[Distribution2.scala 114:31]
  wire  Final_io_Ovalid; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_0_0; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_0_1; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_0_2; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_0_3; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_0_4; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_0_5; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_0_6; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_0_7; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_1_0; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_1_1; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_1_2; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_1_3; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_1_4; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_1_5; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_1_6; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_1_7; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_2_0; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_2_1; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_2_2; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_2_3; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_2_4; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_2_5; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_2_6; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_2_7; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_3_0; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_3_1; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_3_2; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_3_3; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_3_4; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_3_5; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_3_6; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_3_7; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_4_0; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_4_1; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_4_2; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_4_3; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_4_4; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_4_5; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_4_6; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_4_7; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_5_0; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_5_1; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_5_2; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_5_3; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_5_4; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_5_5; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_5_6; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_5_7; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_6_0; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_6_1; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_6_2; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_6_3; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_6_4; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_6_5; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_6_6; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_6_7; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_7_0; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_7_1; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_7_2; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_7_3; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_7_4; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_7_5; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_7_6; // @[Distribution2.scala 114:31]
  wire [31:0] Final_io_omat_7_7; // @[Distribution2.scala 114:31]
  reg [31:0] i; // @[Distribution2.scala 22:20]
  reg [31:0] j; // @[Distribution2.scala 23:20]
  reg [31:0] count; // @[Distribution2.scala 24:24]
  reg [31:0] Idex_0; // @[Distribution2.scala 25:23]
  reg [31:0] Idex_1; // @[Distribution2.scala 25:23]
  reg [31:0] Idex_2; // @[Distribution2.scala 25:23]
  reg [31:0] Idex_3; // @[Distribution2.scala 25:23]
  reg [31:0] Idex_4; // @[Distribution2.scala 25:23]
  reg [31:0] Idex_5; // @[Distribution2.scala 25:23]
  reg [31:0] Idex_6; // @[Distribution2.scala 25:23]
  reg [31:0] Idex_7; // @[Distribution2.scala 25:23]
  reg [31:0] Idex_8; // @[Distribution2.scala 25:23]
  reg [31:0] Idex_9; // @[Distribution2.scala 25:23]
  reg [31:0] Idex_10; // @[Distribution2.scala 25:23]
  reg [31:0] Idex_11; // @[Distribution2.scala 25:23]
  reg [31:0] Idex_12; // @[Distribution2.scala 25:23]
  reg [31:0] Idex_13; // @[Distribution2.scala 25:23]
  reg [31:0] Idex_14; // @[Distribution2.scala 25:23]
  reg [31:0] Idex_15; // @[Distribution2.scala 25:23]
  reg [31:0] Jdex_0; // @[Distribution2.scala 26:23]
  reg [31:0] Jdex_1; // @[Distribution2.scala 26:23]
  reg [31:0] Jdex_2; // @[Distribution2.scala 26:23]
  reg [31:0] Jdex_3; // @[Distribution2.scala 26:23]
  reg [31:0] Jdex_4; // @[Distribution2.scala 26:23]
  reg [31:0] Jdex_5; // @[Distribution2.scala 26:23]
  reg [31:0] Jdex_6; // @[Distribution2.scala 26:23]
  reg [31:0] Jdex_7; // @[Distribution2.scala 26:23]
  reg [31:0] Jdex_8; // @[Distribution2.scala 26:23]
  reg [31:0] Jdex_9; // @[Distribution2.scala 26:23]
  reg [31:0] Jdex_10; // @[Distribution2.scala 26:23]
  reg [31:0] Jdex_11; // @[Distribution2.scala 26:23]
  reg [31:0] Jdex_12; // @[Distribution2.scala 26:23]
  reg [31:0] Jdex_13; // @[Distribution2.scala 26:23]
  reg [31:0] Jdex_14; // @[Distribution2.scala 26:23]
  reg [31:0] Jdex_15; // @[Distribution2.scala 26:23]
  wire [31:0] _GEN_1 = 3'h0 == i[2:0] & 3'h1 == j[2:0] ? io_matrix_0_1 : io_matrix_0_0; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_2 = 3'h0 == i[2:0] & 3'h2 == j[2:0] ? io_matrix_0_2 : _GEN_1; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_3 = 3'h0 == i[2:0] & 3'h3 == j[2:0] ? io_matrix_0_3 : _GEN_2; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_4 = 3'h0 == i[2:0] & 3'h4 == j[2:0] ? io_matrix_0_4 : _GEN_3; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_5 = 3'h0 == i[2:0] & 3'h5 == j[2:0] ? io_matrix_0_5 : _GEN_4; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_6 = 3'h0 == i[2:0] & 3'h6 == j[2:0] ? io_matrix_0_6 : _GEN_5; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_7 = 3'h0 == i[2:0] & 3'h7 == j[2:0] ? io_matrix_0_7 : _GEN_6; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_8 = 3'h1 == i[2:0] & 3'h0 == j[2:0] ? io_matrix_1_0 : _GEN_7; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_9 = 3'h1 == i[2:0] & 3'h1 == j[2:0] ? io_matrix_1_1 : _GEN_8; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_10 = 3'h1 == i[2:0] & 3'h2 == j[2:0] ? io_matrix_1_2 : _GEN_9; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_11 = 3'h1 == i[2:0] & 3'h3 == j[2:0] ? io_matrix_1_3 : _GEN_10; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_12 = 3'h1 == i[2:0] & 3'h4 == j[2:0] ? io_matrix_1_4 : _GEN_11; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_13 = 3'h1 == i[2:0] & 3'h5 == j[2:0] ? io_matrix_1_5 : _GEN_12; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_14 = 3'h1 == i[2:0] & 3'h6 == j[2:0] ? io_matrix_1_6 : _GEN_13; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_15 = 3'h1 == i[2:0] & 3'h7 == j[2:0] ? io_matrix_1_7 : _GEN_14; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_16 = 3'h2 == i[2:0] & 3'h0 == j[2:0] ? io_matrix_2_0 : _GEN_15; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_17 = 3'h2 == i[2:0] & 3'h1 == j[2:0] ? io_matrix_2_1 : _GEN_16; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_18 = 3'h2 == i[2:0] & 3'h2 == j[2:0] ? io_matrix_2_2 : _GEN_17; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_19 = 3'h2 == i[2:0] & 3'h3 == j[2:0] ? io_matrix_2_3 : _GEN_18; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_20 = 3'h2 == i[2:0] & 3'h4 == j[2:0] ? io_matrix_2_4 : _GEN_19; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_21 = 3'h2 == i[2:0] & 3'h5 == j[2:0] ? io_matrix_2_5 : _GEN_20; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_22 = 3'h2 == i[2:0] & 3'h6 == j[2:0] ? io_matrix_2_6 : _GEN_21; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_23 = 3'h2 == i[2:0] & 3'h7 == j[2:0] ? io_matrix_2_7 : _GEN_22; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_24 = 3'h3 == i[2:0] & 3'h0 == j[2:0] ? io_matrix_3_0 : _GEN_23; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_25 = 3'h3 == i[2:0] & 3'h1 == j[2:0] ? io_matrix_3_1 : _GEN_24; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_26 = 3'h3 == i[2:0] & 3'h2 == j[2:0] ? io_matrix_3_2 : _GEN_25; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_27 = 3'h3 == i[2:0] & 3'h3 == j[2:0] ? io_matrix_3_3 : _GEN_26; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_28 = 3'h3 == i[2:0] & 3'h4 == j[2:0] ? io_matrix_3_4 : _GEN_27; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_29 = 3'h3 == i[2:0] & 3'h5 == j[2:0] ? io_matrix_3_5 : _GEN_28; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_30 = 3'h3 == i[2:0] & 3'h6 == j[2:0] ? io_matrix_3_6 : _GEN_29; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_31 = 3'h3 == i[2:0] & 3'h7 == j[2:0] ? io_matrix_3_7 : _GEN_30; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_32 = 3'h4 == i[2:0] & 3'h0 == j[2:0] ? io_matrix_4_0 : _GEN_31; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_33 = 3'h4 == i[2:0] & 3'h1 == j[2:0] ? io_matrix_4_1 : _GEN_32; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_34 = 3'h4 == i[2:0] & 3'h2 == j[2:0] ? io_matrix_4_2 : _GEN_33; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_35 = 3'h4 == i[2:0] & 3'h3 == j[2:0] ? io_matrix_4_3 : _GEN_34; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_36 = 3'h4 == i[2:0] & 3'h4 == j[2:0] ? io_matrix_4_4 : _GEN_35; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_37 = 3'h4 == i[2:0] & 3'h5 == j[2:0] ? io_matrix_4_5 : _GEN_36; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_38 = 3'h4 == i[2:0] & 3'h6 == j[2:0] ? io_matrix_4_6 : _GEN_37; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_39 = 3'h4 == i[2:0] & 3'h7 == j[2:0] ? io_matrix_4_7 : _GEN_38; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_40 = 3'h5 == i[2:0] & 3'h0 == j[2:0] ? io_matrix_5_0 : _GEN_39; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_41 = 3'h5 == i[2:0] & 3'h1 == j[2:0] ? io_matrix_5_1 : _GEN_40; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_42 = 3'h5 == i[2:0] & 3'h2 == j[2:0] ? io_matrix_5_2 : _GEN_41; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_43 = 3'h5 == i[2:0] & 3'h3 == j[2:0] ? io_matrix_5_3 : _GEN_42; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_44 = 3'h5 == i[2:0] & 3'h4 == j[2:0] ? io_matrix_5_4 : _GEN_43; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_45 = 3'h5 == i[2:0] & 3'h5 == j[2:0] ? io_matrix_5_5 : _GEN_44; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_46 = 3'h5 == i[2:0] & 3'h6 == j[2:0] ? io_matrix_5_6 : _GEN_45; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_47 = 3'h5 == i[2:0] & 3'h7 == j[2:0] ? io_matrix_5_7 : _GEN_46; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_48 = 3'h6 == i[2:0] & 3'h0 == j[2:0] ? io_matrix_6_0 : _GEN_47; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_49 = 3'h6 == i[2:0] & 3'h1 == j[2:0] ? io_matrix_6_1 : _GEN_48; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_50 = 3'h6 == i[2:0] & 3'h2 == j[2:0] ? io_matrix_6_2 : _GEN_49; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_51 = 3'h6 == i[2:0] & 3'h3 == j[2:0] ? io_matrix_6_3 : _GEN_50; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_52 = 3'h6 == i[2:0] & 3'h4 == j[2:0] ? io_matrix_6_4 : _GEN_51; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_53 = 3'h6 == i[2:0] & 3'h5 == j[2:0] ? io_matrix_6_5 : _GEN_52; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_54 = 3'h6 == i[2:0] & 3'h6 == j[2:0] ? io_matrix_6_6 : _GEN_53; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_55 = 3'h6 == i[2:0] & 3'h7 == j[2:0] ? io_matrix_6_7 : _GEN_54; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_56 = 3'h7 == i[2:0] & 3'h0 == j[2:0] ? io_matrix_7_0 : _GEN_55; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_57 = 3'h7 == i[2:0] & 3'h1 == j[2:0] ? io_matrix_7_1 : _GEN_56; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_58 = 3'h7 == i[2:0] & 3'h2 == j[2:0] ? io_matrix_7_2 : _GEN_57; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_59 = 3'h7 == i[2:0] & 3'h3 == j[2:0] ? io_matrix_7_3 : _GEN_58; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_60 = 3'h7 == i[2:0] & 3'h4 == j[2:0] ? io_matrix_7_4 : _GEN_59; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_61 = 3'h7 == i[2:0] & 3'h5 == j[2:0] ? io_matrix_7_5 : _GEN_60; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_62 = 3'h7 == i[2:0] & 3'h6 == j[2:0] ? io_matrix_7_6 : _GEN_61; // @[Distribution2.scala 49:{27,27}]
  wire [31:0] _GEN_63 = 3'h7 == i[2:0] & 3'h7 == j[2:0] ? io_matrix_7_7 : _GEN_62; // @[Distribution2.scala 49:{27,27}]
  wire  _T_2 = _GEN_63 == 32'h1; // @[Distribution2.scala 49:27]
  wire [31:0] _count_T_1 = count + 32'h1; // @[Distribution2.scala 62:24]
  wire [31:0] _GEN_129 = 4'h0 == count[3:0] ? i : Idex_0; // @[Distribution2.scala 63:{21,21} 25:23]
  wire [31:0] _GEN_130 = 4'h1 == count[3:0] ? i : Idex_1; // @[Distribution2.scala 63:{21,21} 25:23]
  wire [31:0] _GEN_131 = 4'h2 == count[3:0] ? i : Idex_2; // @[Distribution2.scala 63:{21,21} 25:23]
  wire [31:0] _GEN_132 = 4'h3 == count[3:0] ? i : Idex_3; // @[Distribution2.scala 63:{21,21} 25:23]
  wire [31:0] _GEN_133 = 4'h4 == count[3:0] ? i : Idex_4; // @[Distribution2.scala 63:{21,21} 25:23]
  wire [31:0] _GEN_134 = 4'h5 == count[3:0] ? i : Idex_5; // @[Distribution2.scala 63:{21,21} 25:23]
  wire [31:0] _GEN_135 = 4'h6 == count[3:0] ? i : Idex_6; // @[Distribution2.scala 63:{21,21} 25:23]
  wire [31:0] _GEN_136 = 4'h7 == count[3:0] ? i : Idex_7; // @[Distribution2.scala 63:{21,21} 25:23]
  wire [31:0] _GEN_137 = 4'h8 == count[3:0] ? i : Idex_8; // @[Distribution2.scala 63:{21,21} 25:23]
  wire [31:0] _GEN_138 = 4'h9 == count[3:0] ? i : Idex_9; // @[Distribution2.scala 63:{21,21} 25:23]
  wire [31:0] _GEN_139 = 4'ha == count[3:0] ? i : Idex_10; // @[Distribution2.scala 63:{21,21} 25:23]
  wire [31:0] _GEN_140 = 4'hb == count[3:0] ? i : Idex_11; // @[Distribution2.scala 63:{21,21} 25:23]
  wire [31:0] _GEN_141 = 4'hc == count[3:0] ? i : Idex_12; // @[Distribution2.scala 63:{21,21} 25:23]
  wire [31:0] _GEN_142 = 4'hd == count[3:0] ? i : Idex_13; // @[Distribution2.scala 63:{21,21} 25:23]
  wire [31:0] _GEN_143 = 4'he == count[3:0] ? i : Idex_14; // @[Distribution2.scala 63:{21,21} 25:23]
  wire [31:0] _GEN_144 = 4'hf == count[3:0] ? i : Idex_15; // @[Distribution2.scala 63:{21,21} 25:23]
  wire [31:0] _GEN_145 = 4'h0 == count[3:0] ? j : Jdex_0; // @[Distribution2.scala 64:{21,21} 26:23]
  wire [31:0] _GEN_146 = 4'h1 == count[3:0] ? j : Jdex_1; // @[Distribution2.scala 64:{21,21} 26:23]
  wire [31:0] _GEN_147 = 4'h2 == count[3:0] ? j : Jdex_2; // @[Distribution2.scala 64:{21,21} 26:23]
  wire [31:0] _GEN_148 = 4'h3 == count[3:0] ? j : Jdex_3; // @[Distribution2.scala 64:{21,21} 26:23]
  wire [31:0] _GEN_149 = 4'h4 == count[3:0] ? j : Jdex_4; // @[Distribution2.scala 64:{21,21} 26:23]
  wire [31:0] _GEN_150 = 4'h5 == count[3:0] ? j : Jdex_5; // @[Distribution2.scala 64:{21,21} 26:23]
  wire [31:0] _GEN_151 = 4'h6 == count[3:0] ? j : Jdex_6; // @[Distribution2.scala 64:{21,21} 26:23]
  wire [31:0] _GEN_152 = 4'h7 == count[3:0] ? j : Jdex_7; // @[Distribution2.scala 64:{21,21} 26:23]
  wire [31:0] _GEN_153 = 4'h8 == count[3:0] ? j : Jdex_8; // @[Distribution2.scala 64:{21,21} 26:23]
  wire [31:0] _GEN_154 = 4'h9 == count[3:0] ? j : Jdex_9; // @[Distribution2.scala 64:{21,21} 26:23]
  wire [31:0] _GEN_155 = 4'ha == count[3:0] ? j : Jdex_10; // @[Distribution2.scala 64:{21,21} 26:23]
  wire [31:0] _GEN_156 = 4'hb == count[3:0] ? j : Jdex_11; // @[Distribution2.scala 64:{21,21} 26:23]
  wire [31:0] _GEN_157 = 4'hc == count[3:0] ? j : Jdex_12; // @[Distribution2.scala 64:{21,21} 26:23]
  wire [31:0] _GEN_158 = 4'hd == count[3:0] ? j : Jdex_13; // @[Distribution2.scala 64:{21,21} 26:23]
  wire [31:0] _GEN_159 = 4'he == count[3:0] ? j : Jdex_14; // @[Distribution2.scala 64:{21,21} 26:23]
  wire [31:0] _GEN_160 = 4'hf == count[3:0] ? j : Jdex_15; // @[Distribution2.scala 64:{21,21} 26:23]
  wire  _T_15 = i == 32'h7; // @[Distribution2.scala 65:48]
  wire  _T_17 = j == 32'h7; // @[Distribution2.scala 65:80]
  wire  _complete_T_2 = _T_15 & _T_17; // @[Distribution2.scala 78:55]
  reg  complete; // @[Distribution2.scala 78:27]
  wire [31:0] _GEN_356 = 4'h1 == io_s[3:0] ? Idex_1 : Idex_0; // @[Distribution2.scala 83:{23,23}]
  wire [31:0] _GEN_357 = 4'h2 == io_s[3:0] ? Idex_2 : _GEN_356; // @[Distribution2.scala 83:{23,23}]
  wire [31:0] _GEN_358 = 4'h3 == io_s[3:0] ? Idex_3 : _GEN_357; // @[Distribution2.scala 83:{23,23}]
  wire [31:0] _GEN_359 = 4'h4 == io_s[3:0] ? Idex_4 : _GEN_358; // @[Distribution2.scala 83:{23,23}]
  wire [31:0] _GEN_360 = 4'h5 == io_s[3:0] ? Idex_5 : _GEN_359; // @[Distribution2.scala 83:{23,23}]
  wire [31:0] _GEN_361 = 4'h6 == io_s[3:0] ? Idex_6 : _GEN_360; // @[Distribution2.scala 83:{23,23}]
  wire [31:0] _GEN_362 = 4'h7 == io_s[3:0] ? Idex_7 : _GEN_361; // @[Distribution2.scala 83:{23,23}]
  wire [31:0] _GEN_363 = 4'h8 == io_s[3:0] ? Idex_8 : _GEN_362; // @[Distribution2.scala 83:{23,23}]
  wire [31:0] _GEN_364 = 4'h9 == io_s[3:0] ? Idex_9 : _GEN_363; // @[Distribution2.scala 83:{23,23}]
  wire [31:0] _GEN_365 = 4'ha == io_s[3:0] ? Idex_10 : _GEN_364; // @[Distribution2.scala 83:{23,23}]
  wire [31:0] _GEN_366 = 4'hb == io_s[3:0] ? Idex_11 : _GEN_365; // @[Distribution2.scala 83:{23,23}]
  wire [31:0] _GEN_367 = 4'hc == io_s[3:0] ? Idex_12 : _GEN_366; // @[Distribution2.scala 83:{23,23}]
  wire [31:0] _GEN_368 = 4'hd == io_s[3:0] ? Idex_13 : _GEN_367; // @[Distribution2.scala 83:{23,23}]
  wire [31:0] _GEN_369 = 4'he == io_s[3:0] ? Idex_14 : _GEN_368; // @[Distribution2.scala 83:{23,23}]
  wire [31:0] _GEN_370 = 4'hf == io_s[3:0] ? Idex_15 : _GEN_369; // @[Distribution2.scala 83:{23,23}]
  wire [31:0] _GEN_372 = 4'h1 == io_s[3:0] ? Jdex_1 : Jdex_0; // @[Distribution2.scala 84:{23,23}]
  wire [31:0] _GEN_373 = 4'h2 == io_s[3:0] ? Jdex_2 : _GEN_372; // @[Distribution2.scala 84:{23,23}]
  wire [31:0] _GEN_374 = 4'h3 == io_s[3:0] ? Jdex_3 : _GEN_373; // @[Distribution2.scala 84:{23,23}]
  wire [31:0] _GEN_375 = 4'h4 == io_s[3:0] ? Jdex_4 : _GEN_374; // @[Distribution2.scala 84:{23,23}]
  wire [31:0] _GEN_376 = 4'h5 == io_s[3:0] ? Jdex_5 : _GEN_375; // @[Distribution2.scala 84:{23,23}]
  wire [31:0] _GEN_377 = 4'h6 == io_s[3:0] ? Jdex_6 : _GEN_376; // @[Distribution2.scala 84:{23,23}]
  wire [31:0] _GEN_378 = 4'h7 == io_s[3:0] ? Jdex_7 : _GEN_377; // @[Distribution2.scala 84:{23,23}]
  wire [31:0] _GEN_379 = 4'h8 == io_s[3:0] ? Jdex_8 : _GEN_378; // @[Distribution2.scala 84:{23,23}]
  wire [31:0] _GEN_380 = 4'h9 == io_s[3:0] ? Jdex_9 : _GEN_379; // @[Distribution2.scala 84:{23,23}]
  wire [31:0] _GEN_381 = 4'ha == io_s[3:0] ? Jdex_10 : _GEN_380; // @[Distribution2.scala 84:{23,23}]
  wire [31:0] _GEN_382 = 4'hb == io_s[3:0] ? Jdex_11 : _GEN_381; // @[Distribution2.scala 84:{23,23}]
  wire [31:0] _GEN_383 = 4'hc == io_s[3:0] ? Jdex_12 : _GEN_382; // @[Distribution2.scala 84:{23,23}]
  wire [31:0] _GEN_384 = 4'hd == io_s[3:0] ? Jdex_13 : _GEN_383; // @[Distribution2.scala 84:{23,23}]
  wire [31:0] _GEN_385 = 4'he == io_s[3:0] ? Jdex_14 : _GEN_384; // @[Distribution2.scala 84:{23,23}]
  wire [31:0] _GEN_386 = 4'hf == io_s[3:0] ? Jdex_15 : _GEN_385; // @[Distribution2.scala 84:{23,23}]
  wire [31:0] _T_25 = count - 32'h1; // @[Distribution2.scala 107:84]
  wire  _GEN_453 = part3_io_valid ? Final_io_Ovalid : part2_io_ProcessValid; // @[Distribution2.scala 112:35 127:29 192:29]
  wire [31:0] _GEN_454 = part3_io_valid ? Final_io_omat_0_0 : part2_io_OutMat_0_0; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_455 = part3_io_valid ? Final_io_omat_0_1 : part2_io_OutMat_0_1; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_456 = part3_io_valid ? Final_io_omat_0_2 : part2_io_OutMat_0_2; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_457 = part3_io_valid ? Final_io_omat_0_3 : part2_io_OutMat_0_3; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_458 = part3_io_valid ? Final_io_omat_0_4 : part2_io_OutMat_0_4; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_459 = part3_io_valid ? Final_io_omat_0_5 : part2_io_OutMat_0_5; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_460 = part3_io_valid ? Final_io_omat_0_6 : part2_io_OutMat_0_6; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_461 = part3_io_valid ? Final_io_omat_0_7 : part2_io_OutMat_0_7; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_462 = part3_io_valid ? Final_io_omat_1_0 : part2_io_OutMat_1_0; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_463 = part3_io_valid ? Final_io_omat_1_1 : part2_io_OutMat_1_1; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_464 = part3_io_valid ? Final_io_omat_1_2 : part2_io_OutMat_1_2; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_465 = part3_io_valid ? Final_io_omat_1_3 : part2_io_OutMat_1_3; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_466 = part3_io_valid ? Final_io_omat_1_4 : part2_io_OutMat_1_4; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_467 = part3_io_valid ? Final_io_omat_1_5 : part2_io_OutMat_1_5; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_468 = part3_io_valid ? Final_io_omat_1_6 : part2_io_OutMat_1_6; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_469 = part3_io_valid ? Final_io_omat_1_7 : part2_io_OutMat_1_7; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_470 = part3_io_valid ? Final_io_omat_2_0 : part2_io_OutMat_2_0; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_471 = part3_io_valid ? Final_io_omat_2_1 : part2_io_OutMat_2_1; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_472 = part3_io_valid ? Final_io_omat_2_2 : part2_io_OutMat_2_2; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_473 = part3_io_valid ? Final_io_omat_2_3 : part2_io_OutMat_2_3; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_474 = part3_io_valid ? Final_io_omat_2_4 : part2_io_OutMat_2_4; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_475 = part3_io_valid ? Final_io_omat_2_5 : part2_io_OutMat_2_5; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_476 = part3_io_valid ? Final_io_omat_2_6 : part2_io_OutMat_2_6; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_477 = part3_io_valid ? Final_io_omat_2_7 : part2_io_OutMat_2_7; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_478 = part3_io_valid ? Final_io_omat_3_0 : part2_io_OutMat_3_0; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_479 = part3_io_valid ? Final_io_omat_3_1 : part2_io_OutMat_3_1; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_480 = part3_io_valid ? Final_io_omat_3_2 : part2_io_OutMat_3_2; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_481 = part3_io_valid ? Final_io_omat_3_3 : part2_io_OutMat_3_3; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_482 = part3_io_valid ? Final_io_omat_3_4 : part2_io_OutMat_3_4; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_483 = part3_io_valid ? Final_io_omat_3_5 : part2_io_OutMat_3_5; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_484 = part3_io_valid ? Final_io_omat_3_6 : part2_io_OutMat_3_6; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_485 = part3_io_valid ? Final_io_omat_3_7 : part2_io_OutMat_3_7; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_486 = part3_io_valid ? Final_io_omat_4_0 : part2_io_OutMat_4_0; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_487 = part3_io_valid ? Final_io_omat_4_1 : part2_io_OutMat_4_1; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_488 = part3_io_valid ? Final_io_omat_4_2 : part2_io_OutMat_4_2; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_489 = part3_io_valid ? Final_io_omat_4_3 : part2_io_OutMat_4_3; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_490 = part3_io_valid ? Final_io_omat_4_4 : part2_io_OutMat_4_4; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_491 = part3_io_valid ? Final_io_omat_4_5 : part2_io_OutMat_4_5; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_492 = part3_io_valid ? Final_io_omat_4_6 : part2_io_OutMat_4_6; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_493 = part3_io_valid ? Final_io_omat_4_7 : part2_io_OutMat_4_7; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_494 = part3_io_valid ? Final_io_omat_5_0 : part2_io_OutMat_5_0; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_495 = part3_io_valid ? Final_io_omat_5_1 : part2_io_OutMat_5_1; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_496 = part3_io_valid ? Final_io_omat_5_2 : part2_io_OutMat_5_2; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_497 = part3_io_valid ? Final_io_omat_5_3 : part2_io_OutMat_5_3; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_498 = part3_io_valid ? Final_io_omat_5_4 : part2_io_OutMat_5_4; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_499 = part3_io_valid ? Final_io_omat_5_5 : part2_io_OutMat_5_5; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_500 = part3_io_valid ? Final_io_omat_5_6 : part2_io_OutMat_5_6; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_501 = part3_io_valid ? Final_io_omat_5_7 : part2_io_OutMat_5_7; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_502 = part3_io_valid ? Final_io_omat_6_0 : part2_io_OutMat_6_0; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_503 = part3_io_valid ? Final_io_omat_6_1 : part2_io_OutMat_6_1; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_504 = part3_io_valid ? Final_io_omat_6_2 : part2_io_OutMat_6_2; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_505 = part3_io_valid ? Final_io_omat_6_3 : part2_io_OutMat_6_3; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_506 = part3_io_valid ? Final_io_omat_6_4 : part2_io_OutMat_6_4; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_507 = part3_io_valid ? Final_io_omat_6_5 : part2_io_OutMat_6_5; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_508 = part3_io_valid ? Final_io_omat_6_6 : part2_io_OutMat_6_6; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_509 = part3_io_valid ? Final_io_omat_6_7 : part2_io_OutMat_6_7; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_510 = part3_io_valid ? Final_io_omat_7_0 : part2_io_OutMat_7_0; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_511 = part3_io_valid ? Final_io_omat_7_1 : part2_io_OutMat_7_1; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_512 = part3_io_valid ? Final_io_omat_7_2 : part2_io_OutMat_7_2; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_513 = part3_io_valid ? Final_io_omat_7_3 : part2_io_OutMat_7_3; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_514 = part3_io_valid ? Final_io_omat_7_4 : part2_io_OutMat_7_4; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_515 = part3_io_valid ? Final_io_omat_7_5 : part2_io_OutMat_7_5; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_516 = part3_io_valid ? Final_io_omat_7_6 : part2_io_OutMat_7_6; // @[Distribution2.scala 112:35 128:20 193:20]
  wire [31:0] _GEN_517 = part3_io_valid ? Final_io_omat_7_7 : part2_io_OutMat_7_7; // @[Distribution2.scala 112:35 128:20 193:20]
  wire  _GEN_518 = part2_io_Ovalid & io_valid ? part2_io_ProcessValid : _GEN_453; // @[Distribution2.scala 109:42 110:29]
  wire [31:0] _GEN_519 = part2_io_Ovalid & io_valid ? part2_io_OutMat_0_0 : _GEN_454; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_520 = part2_io_Ovalid & io_valid ? part2_io_OutMat_0_1 : _GEN_455; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_521 = part2_io_Ovalid & io_valid ? part2_io_OutMat_0_2 : _GEN_456; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_522 = part2_io_Ovalid & io_valid ? part2_io_OutMat_0_3 : _GEN_457; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_523 = part2_io_Ovalid & io_valid ? part2_io_OutMat_0_4 : _GEN_458; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_524 = part2_io_Ovalid & io_valid ? part2_io_OutMat_0_5 : _GEN_459; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_525 = part2_io_Ovalid & io_valid ? part2_io_OutMat_0_6 : _GEN_460; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_526 = part2_io_Ovalid & io_valid ? part2_io_OutMat_0_7 : _GEN_461; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_527 = part2_io_Ovalid & io_valid ? part2_io_OutMat_1_0 : _GEN_462; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_528 = part2_io_Ovalid & io_valid ? part2_io_OutMat_1_1 : _GEN_463; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_529 = part2_io_Ovalid & io_valid ? part2_io_OutMat_1_2 : _GEN_464; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_530 = part2_io_Ovalid & io_valid ? part2_io_OutMat_1_3 : _GEN_465; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_531 = part2_io_Ovalid & io_valid ? part2_io_OutMat_1_4 : _GEN_466; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_532 = part2_io_Ovalid & io_valid ? part2_io_OutMat_1_5 : _GEN_467; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_533 = part2_io_Ovalid & io_valid ? part2_io_OutMat_1_6 : _GEN_468; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_534 = part2_io_Ovalid & io_valid ? part2_io_OutMat_1_7 : _GEN_469; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_535 = part2_io_Ovalid & io_valid ? part2_io_OutMat_2_0 : _GEN_470; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_536 = part2_io_Ovalid & io_valid ? part2_io_OutMat_2_1 : _GEN_471; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_537 = part2_io_Ovalid & io_valid ? part2_io_OutMat_2_2 : _GEN_472; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_538 = part2_io_Ovalid & io_valid ? part2_io_OutMat_2_3 : _GEN_473; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_539 = part2_io_Ovalid & io_valid ? part2_io_OutMat_2_4 : _GEN_474; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_540 = part2_io_Ovalid & io_valid ? part2_io_OutMat_2_5 : _GEN_475; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_541 = part2_io_Ovalid & io_valid ? part2_io_OutMat_2_6 : _GEN_476; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_542 = part2_io_Ovalid & io_valid ? part2_io_OutMat_2_7 : _GEN_477; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_543 = part2_io_Ovalid & io_valid ? part2_io_OutMat_3_0 : _GEN_478; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_544 = part2_io_Ovalid & io_valid ? part2_io_OutMat_3_1 : _GEN_479; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_545 = part2_io_Ovalid & io_valid ? part2_io_OutMat_3_2 : _GEN_480; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_546 = part2_io_Ovalid & io_valid ? part2_io_OutMat_3_3 : _GEN_481; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_547 = part2_io_Ovalid & io_valid ? part2_io_OutMat_3_4 : _GEN_482; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_548 = part2_io_Ovalid & io_valid ? part2_io_OutMat_3_5 : _GEN_483; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_549 = part2_io_Ovalid & io_valid ? part2_io_OutMat_3_6 : _GEN_484; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_550 = part2_io_Ovalid & io_valid ? part2_io_OutMat_3_7 : _GEN_485; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_551 = part2_io_Ovalid & io_valid ? part2_io_OutMat_4_0 : _GEN_486; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_552 = part2_io_Ovalid & io_valid ? part2_io_OutMat_4_1 : _GEN_487; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_553 = part2_io_Ovalid & io_valid ? part2_io_OutMat_4_2 : _GEN_488; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_554 = part2_io_Ovalid & io_valid ? part2_io_OutMat_4_3 : _GEN_489; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_555 = part2_io_Ovalid & io_valid ? part2_io_OutMat_4_4 : _GEN_490; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_556 = part2_io_Ovalid & io_valid ? part2_io_OutMat_4_5 : _GEN_491; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_557 = part2_io_Ovalid & io_valid ? part2_io_OutMat_4_6 : _GEN_492; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_558 = part2_io_Ovalid & io_valid ? part2_io_OutMat_4_7 : _GEN_493; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_559 = part2_io_Ovalid & io_valid ? part2_io_OutMat_5_0 : _GEN_494; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_560 = part2_io_Ovalid & io_valid ? part2_io_OutMat_5_1 : _GEN_495; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_561 = part2_io_Ovalid & io_valid ? part2_io_OutMat_5_2 : _GEN_496; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_562 = part2_io_Ovalid & io_valid ? part2_io_OutMat_5_3 : _GEN_497; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_563 = part2_io_Ovalid & io_valid ? part2_io_OutMat_5_4 : _GEN_498; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_564 = part2_io_Ovalid & io_valid ? part2_io_OutMat_5_5 : _GEN_499; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_565 = part2_io_Ovalid & io_valid ? part2_io_OutMat_5_6 : _GEN_500; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_566 = part2_io_Ovalid & io_valid ? part2_io_OutMat_5_7 : _GEN_501; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_567 = part2_io_Ovalid & io_valid ? part2_io_OutMat_6_0 : _GEN_502; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_568 = part2_io_Ovalid & io_valid ? part2_io_OutMat_6_1 : _GEN_503; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_569 = part2_io_Ovalid & io_valid ? part2_io_OutMat_6_2 : _GEN_504; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_570 = part2_io_Ovalid & io_valid ? part2_io_OutMat_6_3 : _GEN_505; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_571 = part2_io_Ovalid & io_valid ? part2_io_OutMat_6_4 : _GEN_506; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_572 = part2_io_Ovalid & io_valid ? part2_io_OutMat_6_5 : _GEN_507; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_573 = part2_io_Ovalid & io_valid ? part2_io_OutMat_6_6 : _GEN_508; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_574 = part2_io_Ovalid & io_valid ? part2_io_OutMat_6_7 : _GEN_509; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_575 = part2_io_Ovalid & io_valid ? part2_io_OutMat_7_0 : _GEN_510; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_576 = part2_io_Ovalid & io_valid ? part2_io_OutMat_7_1 : _GEN_511; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_577 = part2_io_Ovalid & io_valid ? part2_io_OutMat_7_2 : _GEN_512; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_578 = part2_io_Ovalid & io_valid ? part2_io_OutMat_7_3 : _GEN_513; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_579 = part2_io_Ovalid & io_valid ? part2_io_OutMat_7_4 : _GEN_514; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_580 = part2_io_Ovalid & io_valid ? part2_io_OutMat_7_5 : _GEN_515; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_581 = part2_io_Ovalid & io_valid ? part2_io_OutMat_7_6 : _GEN_516; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _GEN_582 = part2_io_Ovalid & io_valid ? part2_io_OutMat_7_7 : _GEN_517; // @[Distribution2.scala 109:42 111:20]
  wire [31:0] _i_T_1 = i + 32'h1; // @[Distribution2.scala 239:16]
  wire [31:0] _j_T_1 = j + 32'h1; // @[Distribution2.scala 242:16]
  SingleLoop2 part2 ( // @[Distribution2.scala 75:23]
    .clock(part2_clock),
    .reset(part2_reset),
    .io_IDex(part2_io_IDex),
    .io_JDex(part2_io_JDex),
    .io_valid(part2_io_valid),
    .io_mat_0_0(part2_io_mat_0_0),
    .io_mat_0_1(part2_io_mat_0_1),
    .io_mat_0_2(part2_io_mat_0_2),
    .io_mat_0_3(part2_io_mat_0_3),
    .io_mat_0_4(part2_io_mat_0_4),
    .io_mat_0_5(part2_io_mat_0_5),
    .io_mat_0_6(part2_io_mat_0_6),
    .io_mat_0_7(part2_io_mat_0_7),
    .io_mat_1_0(part2_io_mat_1_0),
    .io_mat_1_1(part2_io_mat_1_1),
    .io_mat_1_2(part2_io_mat_1_2),
    .io_mat_1_3(part2_io_mat_1_3),
    .io_mat_1_4(part2_io_mat_1_4),
    .io_mat_1_5(part2_io_mat_1_5),
    .io_mat_1_6(part2_io_mat_1_6),
    .io_mat_1_7(part2_io_mat_1_7),
    .io_mat_2_0(part2_io_mat_2_0),
    .io_mat_2_1(part2_io_mat_2_1),
    .io_mat_2_2(part2_io_mat_2_2),
    .io_mat_2_3(part2_io_mat_2_3),
    .io_mat_2_4(part2_io_mat_2_4),
    .io_mat_2_5(part2_io_mat_2_5),
    .io_mat_2_6(part2_io_mat_2_6),
    .io_mat_2_7(part2_io_mat_2_7),
    .io_mat_3_0(part2_io_mat_3_0),
    .io_mat_3_1(part2_io_mat_3_1),
    .io_mat_3_2(part2_io_mat_3_2),
    .io_mat_3_3(part2_io_mat_3_3),
    .io_mat_3_4(part2_io_mat_3_4),
    .io_mat_3_5(part2_io_mat_3_5),
    .io_mat_3_6(part2_io_mat_3_6),
    .io_mat_3_7(part2_io_mat_3_7),
    .io_mat_4_0(part2_io_mat_4_0),
    .io_mat_4_1(part2_io_mat_4_1),
    .io_mat_4_2(part2_io_mat_4_2),
    .io_mat_4_3(part2_io_mat_4_3),
    .io_mat_4_4(part2_io_mat_4_4),
    .io_mat_4_5(part2_io_mat_4_5),
    .io_mat_4_6(part2_io_mat_4_6),
    .io_mat_4_7(part2_io_mat_4_7),
    .io_mat_5_0(part2_io_mat_5_0),
    .io_mat_5_1(part2_io_mat_5_1),
    .io_mat_5_2(part2_io_mat_5_2),
    .io_mat_5_3(part2_io_mat_5_3),
    .io_mat_5_4(part2_io_mat_5_4),
    .io_mat_5_5(part2_io_mat_5_5),
    .io_mat_5_6(part2_io_mat_5_6),
    .io_mat_5_7(part2_io_mat_5_7),
    .io_mat_6_0(part2_io_mat_6_0),
    .io_mat_6_1(part2_io_mat_6_1),
    .io_mat_6_2(part2_io_mat_6_2),
    .io_mat_6_3(part2_io_mat_6_3),
    .io_mat_6_4(part2_io_mat_6_4),
    .io_mat_6_5(part2_io_mat_6_5),
    .io_mat_6_6(part2_io_mat_6_6),
    .io_mat_6_7(part2_io_mat_6_7),
    .io_mat_7_0(part2_io_mat_7_0),
    .io_mat_7_1(part2_io_mat_7_1),
    .io_mat_7_2(part2_io_mat_7_2),
    .io_mat_7_3(part2_io_mat_7_3),
    .io_mat_7_4(part2_io_mat_7_4),
    .io_mat_7_5(part2_io_mat_7_5),
    .io_mat_7_6(part2_io_mat_7_6),
    .io_mat_7_7(part2_io_mat_7_7),
    .io_OutMat_0_0(part2_io_OutMat_0_0),
    .io_OutMat_0_1(part2_io_OutMat_0_1),
    .io_OutMat_0_2(part2_io_OutMat_0_2),
    .io_OutMat_0_3(part2_io_OutMat_0_3),
    .io_OutMat_0_4(part2_io_OutMat_0_4),
    .io_OutMat_0_5(part2_io_OutMat_0_5),
    .io_OutMat_0_6(part2_io_OutMat_0_6),
    .io_OutMat_0_7(part2_io_OutMat_0_7),
    .io_OutMat_1_0(part2_io_OutMat_1_0),
    .io_OutMat_1_1(part2_io_OutMat_1_1),
    .io_OutMat_1_2(part2_io_OutMat_1_2),
    .io_OutMat_1_3(part2_io_OutMat_1_3),
    .io_OutMat_1_4(part2_io_OutMat_1_4),
    .io_OutMat_1_5(part2_io_OutMat_1_5),
    .io_OutMat_1_6(part2_io_OutMat_1_6),
    .io_OutMat_1_7(part2_io_OutMat_1_7),
    .io_OutMat_2_0(part2_io_OutMat_2_0),
    .io_OutMat_2_1(part2_io_OutMat_2_1),
    .io_OutMat_2_2(part2_io_OutMat_2_2),
    .io_OutMat_2_3(part2_io_OutMat_2_3),
    .io_OutMat_2_4(part2_io_OutMat_2_4),
    .io_OutMat_2_5(part2_io_OutMat_2_5),
    .io_OutMat_2_6(part2_io_OutMat_2_6),
    .io_OutMat_2_7(part2_io_OutMat_2_7),
    .io_OutMat_3_0(part2_io_OutMat_3_0),
    .io_OutMat_3_1(part2_io_OutMat_3_1),
    .io_OutMat_3_2(part2_io_OutMat_3_2),
    .io_OutMat_3_3(part2_io_OutMat_3_3),
    .io_OutMat_3_4(part2_io_OutMat_3_4),
    .io_OutMat_3_5(part2_io_OutMat_3_5),
    .io_OutMat_3_6(part2_io_OutMat_3_6),
    .io_OutMat_3_7(part2_io_OutMat_3_7),
    .io_OutMat_4_0(part2_io_OutMat_4_0),
    .io_OutMat_4_1(part2_io_OutMat_4_1),
    .io_OutMat_4_2(part2_io_OutMat_4_2),
    .io_OutMat_4_3(part2_io_OutMat_4_3),
    .io_OutMat_4_4(part2_io_OutMat_4_4),
    .io_OutMat_4_5(part2_io_OutMat_4_5),
    .io_OutMat_4_6(part2_io_OutMat_4_6),
    .io_OutMat_4_7(part2_io_OutMat_4_7),
    .io_OutMat_5_0(part2_io_OutMat_5_0),
    .io_OutMat_5_1(part2_io_OutMat_5_1),
    .io_OutMat_5_2(part2_io_OutMat_5_2),
    .io_OutMat_5_3(part2_io_OutMat_5_3),
    .io_OutMat_5_4(part2_io_OutMat_5_4),
    .io_OutMat_5_5(part2_io_OutMat_5_5),
    .io_OutMat_5_6(part2_io_OutMat_5_6),
    .io_OutMat_5_7(part2_io_OutMat_5_7),
    .io_OutMat_6_0(part2_io_OutMat_6_0),
    .io_OutMat_6_1(part2_io_OutMat_6_1),
    .io_OutMat_6_2(part2_io_OutMat_6_2),
    .io_OutMat_6_3(part2_io_OutMat_6_3),
    .io_OutMat_6_4(part2_io_OutMat_6_4),
    .io_OutMat_6_5(part2_io_OutMat_6_5),
    .io_OutMat_6_6(part2_io_OutMat_6_6),
    .io_OutMat_6_7(part2_io_OutMat_6_7),
    .io_OutMat_7_0(part2_io_OutMat_7_0),
    .io_OutMat_7_1(part2_io_OutMat_7_1),
    .io_OutMat_7_2(part2_io_OutMat_7_2),
    .io_OutMat_7_3(part2_io_OutMat_7_3),
    .io_OutMat_7_4(part2_io_OutMat_7_4),
    .io_OutMat_7_5(part2_io_OutMat_7_5),
    .io_OutMat_7_6(part2_io_OutMat_7_6),
    .io_OutMat_7_7(part2_io_OutMat_7_7),
    .io_Ovalid(part2_io_Ovalid),
    .io_ProcessValid(part2_io_ProcessValid)
  );
  MergeDistribution2 part3 ( // @[Distribution2.scala 90:23]
    .clock(part3_clock),
    .reset(part3_reset),
    .io_IDex(part3_io_IDex),
    .io_mat_0_0(part3_io_mat_0_0),
    .io_mat_0_1(part3_io_mat_0_1),
    .io_mat_0_2(part3_io_mat_0_2),
    .io_mat_0_3(part3_io_mat_0_3),
    .io_mat_0_4(part3_io_mat_0_4),
    .io_mat_0_5(part3_io_mat_0_5),
    .io_mat_0_6(part3_io_mat_0_6),
    .io_mat_0_7(part3_io_mat_0_7),
    .io_mat_1_0(part3_io_mat_1_0),
    .io_mat_1_1(part3_io_mat_1_1),
    .io_mat_1_2(part3_io_mat_1_2),
    .io_mat_1_3(part3_io_mat_1_3),
    .io_mat_1_4(part3_io_mat_1_4),
    .io_mat_1_5(part3_io_mat_1_5),
    .io_mat_1_6(part3_io_mat_1_6),
    .io_mat_1_7(part3_io_mat_1_7),
    .io_mat_2_0(part3_io_mat_2_0),
    .io_mat_2_1(part3_io_mat_2_1),
    .io_mat_2_2(part3_io_mat_2_2),
    .io_mat_2_3(part3_io_mat_2_3),
    .io_mat_2_4(part3_io_mat_2_4),
    .io_mat_2_5(part3_io_mat_2_5),
    .io_mat_2_6(part3_io_mat_2_6),
    .io_mat_2_7(part3_io_mat_2_7),
    .io_mat_3_0(part3_io_mat_3_0),
    .io_mat_3_1(part3_io_mat_3_1),
    .io_mat_3_2(part3_io_mat_3_2),
    .io_mat_3_3(part3_io_mat_3_3),
    .io_mat_3_4(part3_io_mat_3_4),
    .io_mat_3_5(part3_io_mat_3_5),
    .io_mat_3_6(part3_io_mat_3_6),
    .io_mat_3_7(part3_io_mat_3_7),
    .io_mat_4_0(part3_io_mat_4_0),
    .io_mat_4_1(part3_io_mat_4_1),
    .io_mat_4_2(part3_io_mat_4_2),
    .io_mat_4_3(part3_io_mat_4_3),
    .io_mat_4_4(part3_io_mat_4_4),
    .io_mat_4_5(part3_io_mat_4_5),
    .io_mat_4_6(part3_io_mat_4_6),
    .io_mat_4_7(part3_io_mat_4_7),
    .io_mat_5_0(part3_io_mat_5_0),
    .io_mat_5_1(part3_io_mat_5_1),
    .io_mat_5_2(part3_io_mat_5_2),
    .io_mat_5_3(part3_io_mat_5_3),
    .io_mat_5_4(part3_io_mat_5_4),
    .io_mat_5_5(part3_io_mat_5_5),
    .io_mat_5_6(part3_io_mat_5_6),
    .io_mat_5_7(part3_io_mat_5_7),
    .io_mat_6_0(part3_io_mat_6_0),
    .io_mat_6_1(part3_io_mat_6_1),
    .io_mat_6_2(part3_io_mat_6_2),
    .io_mat_6_3(part3_io_mat_6_3),
    .io_mat_6_4(part3_io_mat_6_4),
    .io_mat_6_5(part3_io_mat_6_5),
    .io_mat_6_6(part3_io_mat_6_6),
    .io_mat_6_7(part3_io_mat_6_7),
    .io_mat_7_0(part3_io_mat_7_0),
    .io_mat_7_1(part3_io_mat_7_1),
    .io_mat_7_2(part3_io_mat_7_2),
    .io_mat_7_3(part3_io_mat_7_3),
    .io_mat_7_4(part3_io_mat_7_4),
    .io_mat_7_5(part3_io_mat_7_5),
    .io_mat_7_6(part3_io_mat_7_6),
    .io_mat_7_7(part3_io_mat_7_7),
    .io_i_valid(part3_io_i_valid),
    .io_valid(part3_io_valid),
    .io_Omat_0_0(part3_io_Omat_0_0),
    .io_Omat_0_1(part3_io_Omat_0_1),
    .io_Omat_0_2(part3_io_Omat_0_2),
    .io_Omat_0_3(part3_io_Omat_0_3),
    .io_Omat_0_4(part3_io_Omat_0_4),
    .io_Omat_0_5(part3_io_Omat_0_5),
    .io_Omat_0_6(part3_io_Omat_0_6),
    .io_Omat_0_7(part3_io_Omat_0_7),
    .io_Omat_1_0(part3_io_Omat_1_0),
    .io_Omat_1_1(part3_io_Omat_1_1),
    .io_Omat_1_2(part3_io_Omat_1_2),
    .io_Omat_1_3(part3_io_Omat_1_3),
    .io_Omat_1_4(part3_io_Omat_1_4),
    .io_Omat_1_5(part3_io_Omat_1_5),
    .io_Omat_1_6(part3_io_Omat_1_6),
    .io_Omat_1_7(part3_io_Omat_1_7),
    .io_Omat_2_0(part3_io_Omat_2_0),
    .io_Omat_2_1(part3_io_Omat_2_1),
    .io_Omat_2_2(part3_io_Omat_2_2),
    .io_Omat_2_3(part3_io_Omat_2_3),
    .io_Omat_2_4(part3_io_Omat_2_4),
    .io_Omat_2_5(part3_io_Omat_2_5),
    .io_Omat_2_6(part3_io_Omat_2_6),
    .io_Omat_2_7(part3_io_Omat_2_7),
    .io_Omat_3_0(part3_io_Omat_3_0),
    .io_Omat_3_1(part3_io_Omat_3_1),
    .io_Omat_3_2(part3_io_Omat_3_2),
    .io_Omat_3_3(part3_io_Omat_3_3),
    .io_Omat_3_4(part3_io_Omat_3_4),
    .io_Omat_3_5(part3_io_Omat_3_5),
    .io_Omat_3_6(part3_io_Omat_3_6),
    .io_Omat_3_7(part3_io_Omat_3_7),
    .io_Omat_4_0(part3_io_Omat_4_0),
    .io_Omat_4_1(part3_io_Omat_4_1),
    .io_Omat_4_2(part3_io_Omat_4_2),
    .io_Omat_4_3(part3_io_Omat_4_3),
    .io_Omat_4_4(part3_io_Omat_4_4),
    .io_Omat_4_5(part3_io_Omat_4_5),
    .io_Omat_4_6(part3_io_Omat_4_6),
    .io_Omat_4_7(part3_io_Omat_4_7),
    .io_Omat_5_0(part3_io_Omat_5_0),
    .io_Omat_5_1(part3_io_Omat_5_1),
    .io_Omat_5_2(part3_io_Omat_5_2),
    .io_Omat_5_3(part3_io_Omat_5_3),
    .io_Omat_5_4(part3_io_Omat_5_4),
    .io_Omat_5_5(part3_io_Omat_5_5),
    .io_Omat_5_6(part3_io_Omat_5_6),
    .io_Omat_5_7(part3_io_Omat_5_7),
    .io_Omat_6_0(part3_io_Omat_6_0),
    .io_Omat_6_1(part3_io_Omat_6_1),
    .io_Omat_6_2(part3_io_Omat_6_2),
    .io_Omat_6_3(part3_io_Omat_6_3),
    .io_Omat_6_4(part3_io_Omat_6_4),
    .io_Omat_6_5(part3_io_Omat_6_5),
    .io_Omat_6_6(part3_io_Omat_6_6),
    .io_Omat_6_7(part3_io_Omat_6_7),
    .io_Omat_7_0(part3_io_Omat_7_0),
    .io_Omat_7_1(part3_io_Omat_7_1),
    .io_Omat_7_2(part3_io_Omat_7_2),
    .io_Omat_7_3(part3_io_Omat_7_3),
    .io_Omat_7_4(part3_io_Omat_7_4),
    .io_Omat_7_5(part3_io_Omat_7_5),
    .io_Omat_7_6(part3_io_Omat_7_6),
    .io_Omat_7_7(part3_io_Omat_7_7)
  );
  FinalMerge Final ( // @[Distribution2.scala 114:31]
    .clock(Final_clock),
    .reset(Final_reset),
    .io_IDex(Final_io_IDex),
    .io_PreMat_0_0(Final_io_PreMat_0_0),
    .io_PreMat_0_1(Final_io_PreMat_0_1),
    .io_PreMat_0_2(Final_io_PreMat_0_2),
    .io_PreMat_0_3(Final_io_PreMat_0_3),
    .io_PreMat_0_4(Final_io_PreMat_0_4),
    .io_PreMat_0_5(Final_io_PreMat_0_5),
    .io_PreMat_0_6(Final_io_PreMat_0_6),
    .io_PreMat_0_7(Final_io_PreMat_0_7),
    .io_PreMat_1_0(Final_io_PreMat_1_0),
    .io_PreMat_1_1(Final_io_PreMat_1_1),
    .io_PreMat_1_2(Final_io_PreMat_1_2),
    .io_PreMat_1_3(Final_io_PreMat_1_3),
    .io_PreMat_1_4(Final_io_PreMat_1_4),
    .io_PreMat_1_5(Final_io_PreMat_1_5),
    .io_PreMat_1_6(Final_io_PreMat_1_6),
    .io_PreMat_1_7(Final_io_PreMat_1_7),
    .io_PreMat_2_0(Final_io_PreMat_2_0),
    .io_PreMat_2_1(Final_io_PreMat_2_1),
    .io_PreMat_2_2(Final_io_PreMat_2_2),
    .io_PreMat_2_3(Final_io_PreMat_2_3),
    .io_PreMat_2_4(Final_io_PreMat_2_4),
    .io_PreMat_2_5(Final_io_PreMat_2_5),
    .io_PreMat_2_6(Final_io_PreMat_2_6),
    .io_PreMat_2_7(Final_io_PreMat_2_7),
    .io_PreMat_3_0(Final_io_PreMat_3_0),
    .io_PreMat_3_1(Final_io_PreMat_3_1),
    .io_PreMat_3_2(Final_io_PreMat_3_2),
    .io_PreMat_3_3(Final_io_PreMat_3_3),
    .io_PreMat_3_4(Final_io_PreMat_3_4),
    .io_PreMat_3_5(Final_io_PreMat_3_5),
    .io_PreMat_3_6(Final_io_PreMat_3_6),
    .io_PreMat_3_7(Final_io_PreMat_3_7),
    .io_PreMat_4_0(Final_io_PreMat_4_0),
    .io_PreMat_4_1(Final_io_PreMat_4_1),
    .io_PreMat_4_2(Final_io_PreMat_4_2),
    .io_PreMat_4_3(Final_io_PreMat_4_3),
    .io_PreMat_4_4(Final_io_PreMat_4_4),
    .io_PreMat_4_5(Final_io_PreMat_4_5),
    .io_PreMat_4_6(Final_io_PreMat_4_6),
    .io_PreMat_4_7(Final_io_PreMat_4_7),
    .io_PreMat_5_0(Final_io_PreMat_5_0),
    .io_PreMat_5_1(Final_io_PreMat_5_1),
    .io_PreMat_5_2(Final_io_PreMat_5_2),
    .io_PreMat_5_3(Final_io_PreMat_5_3),
    .io_PreMat_5_4(Final_io_PreMat_5_4),
    .io_PreMat_5_5(Final_io_PreMat_5_5),
    .io_PreMat_5_6(Final_io_PreMat_5_6),
    .io_PreMat_5_7(Final_io_PreMat_5_7),
    .io_PreMat_6_0(Final_io_PreMat_6_0),
    .io_PreMat_6_1(Final_io_PreMat_6_1),
    .io_PreMat_6_2(Final_io_PreMat_6_2),
    .io_PreMat_6_3(Final_io_PreMat_6_3),
    .io_PreMat_6_4(Final_io_PreMat_6_4),
    .io_PreMat_6_5(Final_io_PreMat_6_5),
    .io_PreMat_6_6(Final_io_PreMat_6_6),
    .io_PreMat_6_7(Final_io_PreMat_6_7),
    .io_PreMat_7_0(Final_io_PreMat_7_0),
    .io_PreMat_7_1(Final_io_PreMat_7_1),
    .io_PreMat_7_2(Final_io_PreMat_7_2),
    .io_PreMat_7_3(Final_io_PreMat_7_3),
    .io_PreMat_7_4(Final_io_PreMat_7_4),
    .io_PreMat_7_5(Final_io_PreMat_7_5),
    .io_PreMat_7_6(Final_io_PreMat_7_6),
    .io_PreMat_7_7(Final_io_PreMat_7_7),
    .io_lastMat_0_0(Final_io_lastMat_0_0),
    .io_lastMat_0_1(Final_io_lastMat_0_1),
    .io_lastMat_0_2(Final_io_lastMat_0_2),
    .io_lastMat_0_3(Final_io_lastMat_0_3),
    .io_lastMat_0_4(Final_io_lastMat_0_4),
    .io_lastMat_0_5(Final_io_lastMat_0_5),
    .io_lastMat_0_6(Final_io_lastMat_0_6),
    .io_lastMat_0_7(Final_io_lastMat_0_7),
    .io_lastMat_1_0(Final_io_lastMat_1_0),
    .io_lastMat_1_1(Final_io_lastMat_1_1),
    .io_lastMat_1_2(Final_io_lastMat_1_2),
    .io_lastMat_1_3(Final_io_lastMat_1_3),
    .io_lastMat_1_4(Final_io_lastMat_1_4),
    .io_lastMat_1_5(Final_io_lastMat_1_5),
    .io_lastMat_1_6(Final_io_lastMat_1_6),
    .io_lastMat_1_7(Final_io_lastMat_1_7),
    .io_lastMat_2_0(Final_io_lastMat_2_0),
    .io_lastMat_2_1(Final_io_lastMat_2_1),
    .io_lastMat_2_2(Final_io_lastMat_2_2),
    .io_lastMat_2_3(Final_io_lastMat_2_3),
    .io_lastMat_2_4(Final_io_lastMat_2_4),
    .io_lastMat_2_5(Final_io_lastMat_2_5),
    .io_lastMat_2_6(Final_io_lastMat_2_6),
    .io_lastMat_2_7(Final_io_lastMat_2_7),
    .io_lastMat_3_0(Final_io_lastMat_3_0),
    .io_lastMat_3_1(Final_io_lastMat_3_1),
    .io_lastMat_3_2(Final_io_lastMat_3_2),
    .io_lastMat_3_3(Final_io_lastMat_3_3),
    .io_lastMat_3_4(Final_io_lastMat_3_4),
    .io_lastMat_3_5(Final_io_lastMat_3_5),
    .io_lastMat_3_6(Final_io_lastMat_3_6),
    .io_lastMat_3_7(Final_io_lastMat_3_7),
    .io_lastMat_4_0(Final_io_lastMat_4_0),
    .io_lastMat_4_1(Final_io_lastMat_4_1),
    .io_lastMat_4_2(Final_io_lastMat_4_2),
    .io_lastMat_4_3(Final_io_lastMat_4_3),
    .io_lastMat_4_4(Final_io_lastMat_4_4),
    .io_lastMat_4_5(Final_io_lastMat_4_5),
    .io_lastMat_4_6(Final_io_lastMat_4_6),
    .io_lastMat_4_7(Final_io_lastMat_4_7),
    .io_lastMat_5_0(Final_io_lastMat_5_0),
    .io_lastMat_5_1(Final_io_lastMat_5_1),
    .io_lastMat_5_2(Final_io_lastMat_5_2),
    .io_lastMat_5_3(Final_io_lastMat_5_3),
    .io_lastMat_5_4(Final_io_lastMat_5_4),
    .io_lastMat_5_5(Final_io_lastMat_5_5),
    .io_lastMat_5_6(Final_io_lastMat_5_6),
    .io_lastMat_5_7(Final_io_lastMat_5_7),
    .io_lastMat_6_0(Final_io_lastMat_6_0),
    .io_lastMat_6_1(Final_io_lastMat_6_1),
    .io_lastMat_6_2(Final_io_lastMat_6_2),
    .io_lastMat_6_3(Final_io_lastMat_6_3),
    .io_lastMat_6_4(Final_io_lastMat_6_4),
    .io_lastMat_6_5(Final_io_lastMat_6_5),
    .io_lastMat_6_6(Final_io_lastMat_6_6),
    .io_lastMat_6_7(Final_io_lastMat_6_7),
    .io_lastMat_7_0(Final_io_lastMat_7_0),
    .io_lastMat_7_1(Final_io_lastMat_7_1),
    .io_lastMat_7_2(Final_io_lastMat_7_2),
    .io_lastMat_7_3(Final_io_lastMat_7_3),
    .io_lastMat_7_4(Final_io_lastMat_7_4),
    .io_lastMat_7_5(Final_io_lastMat_7_5),
    .io_lastMat_7_6(Final_io_lastMat_7_6),
    .io_lastMat_7_7(Final_io_lastMat_7_7),
    .io_valid(Final_io_valid),
    .io_Ovalid(Final_io_Ovalid),
    .io_omat_0_0(Final_io_omat_0_0),
    .io_omat_0_1(Final_io_omat_0_1),
    .io_omat_0_2(Final_io_omat_0_2),
    .io_omat_0_3(Final_io_omat_0_3),
    .io_omat_0_4(Final_io_omat_0_4),
    .io_omat_0_5(Final_io_omat_0_5),
    .io_omat_0_6(Final_io_omat_0_6),
    .io_omat_0_7(Final_io_omat_0_7),
    .io_omat_1_0(Final_io_omat_1_0),
    .io_omat_1_1(Final_io_omat_1_1),
    .io_omat_1_2(Final_io_omat_1_2),
    .io_omat_1_3(Final_io_omat_1_3),
    .io_omat_1_4(Final_io_omat_1_4),
    .io_omat_1_5(Final_io_omat_1_5),
    .io_omat_1_6(Final_io_omat_1_6),
    .io_omat_1_7(Final_io_omat_1_7),
    .io_omat_2_0(Final_io_omat_2_0),
    .io_omat_2_1(Final_io_omat_2_1),
    .io_omat_2_2(Final_io_omat_2_2),
    .io_omat_2_3(Final_io_omat_2_3),
    .io_omat_2_4(Final_io_omat_2_4),
    .io_omat_2_5(Final_io_omat_2_5),
    .io_omat_2_6(Final_io_omat_2_6),
    .io_omat_2_7(Final_io_omat_2_7),
    .io_omat_3_0(Final_io_omat_3_0),
    .io_omat_3_1(Final_io_omat_3_1),
    .io_omat_3_2(Final_io_omat_3_2),
    .io_omat_3_3(Final_io_omat_3_3),
    .io_omat_3_4(Final_io_omat_3_4),
    .io_omat_3_5(Final_io_omat_3_5),
    .io_omat_3_6(Final_io_omat_3_6),
    .io_omat_3_7(Final_io_omat_3_7),
    .io_omat_4_0(Final_io_omat_4_0),
    .io_omat_4_1(Final_io_omat_4_1),
    .io_omat_4_2(Final_io_omat_4_2),
    .io_omat_4_3(Final_io_omat_4_3),
    .io_omat_4_4(Final_io_omat_4_4),
    .io_omat_4_5(Final_io_omat_4_5),
    .io_omat_4_6(Final_io_omat_4_6),
    .io_omat_4_7(Final_io_omat_4_7),
    .io_omat_5_0(Final_io_omat_5_0),
    .io_omat_5_1(Final_io_omat_5_1),
    .io_omat_5_2(Final_io_omat_5_2),
    .io_omat_5_3(Final_io_omat_5_3),
    .io_omat_5_4(Final_io_omat_5_4),
    .io_omat_5_5(Final_io_omat_5_5),
    .io_omat_5_6(Final_io_omat_5_6),
    .io_omat_5_7(Final_io_omat_5_7),
    .io_omat_6_0(Final_io_omat_6_0),
    .io_omat_6_1(Final_io_omat_6_1),
    .io_omat_6_2(Final_io_omat_6_2),
    .io_omat_6_3(Final_io_omat_6_3),
    .io_omat_6_4(Final_io_omat_6_4),
    .io_omat_6_5(Final_io_omat_6_5),
    .io_omat_6_6(Final_io_omat_6_6),
    .io_omat_6_7(Final_io_omat_6_7),
    .io_omat_7_0(Final_io_omat_7_0),
    .io_omat_7_1(Final_io_omat_7_1),
    .io_omat_7_2(Final_io_omat_7_2),
    .io_omat_7_3(Final_io_omat_7_3),
    .io_omat_7_4(Final_io_omat_7_4),
    .io_omat_7_5(Final_io_omat_7_5),
    .io_omat_7_6(Final_io_omat_7_6),
    .io_omat_7_7(Final_io_omat_7_7)
  );
  assign io_out_0_0 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_519 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_0_1 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_520 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_0_2 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_521 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_0_3 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_522 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_0_4 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_523 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_0_5 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_524 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_0_6 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_525 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_0_7 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_526 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_1_0 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_527 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_1_1 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_528 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_1_2 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_529 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_1_3 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_530 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_1_4 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_531 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_1_5 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_532 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_1_6 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_533 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_1_7 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_534 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_2_0 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_535 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_2_1 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_536 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_2_2 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_537 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_2_3 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_538 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_2_4 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_539 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_2_5 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_540 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_2_6 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_541 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_2_7 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_542 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_3_0 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_543 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_3_1 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_544 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_3_2 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_545 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_3_3 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_546 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_3_4 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_547 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_3_5 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_548 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_3_6 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_549 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_3_7 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_550 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_4_0 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_551 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_4_1 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_552 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_4_2 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_553 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_4_3 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_554 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_4_4 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_555 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_4_5 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_556 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_4_6 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_557 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_4_7 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_558 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_5_0 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_559 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_5_1 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_560 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_5_2 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_561 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_5_3 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_562 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_5_4 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_563 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_5_5 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_564 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_5_6 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_565 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_5_7 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_566 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_6_0 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_567 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_6_1 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_568 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_6_2 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_569 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_6_3 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_570 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_6_4 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_571 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_6_5 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_572 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_6_6 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_573 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_6_7 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_574 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_7_0 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_575 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_7_1 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_576 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_7_2 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_577 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_7_3 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_578 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_7_4 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_579 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_7_5 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_580 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_7_6 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_581 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_out_7_7 = ~(_complete_T_2 & _T_25 < io_s) ? _GEN_582 : 32'h0; // @[Distribution2.scala 107:99 196:16]
  assign io_ProcessValid = ~(_complete_T_2 & _T_25 < io_s) & _GEN_518; // @[Distribution2.scala 107:99 197:25]
  assign part2_clock = clock;
  assign part2_reset = reset;
  assign part2_io_IDex = complete ? _GEN_370 : 32'h0; // @[Distribution2.scala 82:20 83:23 86:23]
  assign part2_io_JDex = complete ? _GEN_386 : 32'h0; // @[Distribution2.scala 82:20 84:23 87:23]
  assign part2_io_valid = complete; // @[Distribution2.scala 80:20]
  assign part2_io_mat_0_0 = io_matrix_0_0; // @[Distribution2.scala 76:18]
  assign part2_io_mat_0_1 = io_matrix_0_1; // @[Distribution2.scala 76:18]
  assign part2_io_mat_0_2 = io_matrix_0_2; // @[Distribution2.scala 76:18]
  assign part2_io_mat_0_3 = io_matrix_0_3; // @[Distribution2.scala 76:18]
  assign part2_io_mat_0_4 = io_matrix_0_4; // @[Distribution2.scala 76:18]
  assign part2_io_mat_0_5 = io_matrix_0_5; // @[Distribution2.scala 76:18]
  assign part2_io_mat_0_6 = io_matrix_0_6; // @[Distribution2.scala 76:18]
  assign part2_io_mat_0_7 = io_matrix_0_7; // @[Distribution2.scala 76:18]
  assign part2_io_mat_1_0 = io_matrix_1_0; // @[Distribution2.scala 76:18]
  assign part2_io_mat_1_1 = io_matrix_1_1; // @[Distribution2.scala 76:18]
  assign part2_io_mat_1_2 = io_matrix_1_2; // @[Distribution2.scala 76:18]
  assign part2_io_mat_1_3 = io_matrix_1_3; // @[Distribution2.scala 76:18]
  assign part2_io_mat_1_4 = io_matrix_1_4; // @[Distribution2.scala 76:18]
  assign part2_io_mat_1_5 = io_matrix_1_5; // @[Distribution2.scala 76:18]
  assign part2_io_mat_1_6 = io_matrix_1_6; // @[Distribution2.scala 76:18]
  assign part2_io_mat_1_7 = io_matrix_1_7; // @[Distribution2.scala 76:18]
  assign part2_io_mat_2_0 = io_matrix_2_0; // @[Distribution2.scala 76:18]
  assign part2_io_mat_2_1 = io_matrix_2_1; // @[Distribution2.scala 76:18]
  assign part2_io_mat_2_2 = io_matrix_2_2; // @[Distribution2.scala 76:18]
  assign part2_io_mat_2_3 = io_matrix_2_3; // @[Distribution2.scala 76:18]
  assign part2_io_mat_2_4 = io_matrix_2_4; // @[Distribution2.scala 76:18]
  assign part2_io_mat_2_5 = io_matrix_2_5; // @[Distribution2.scala 76:18]
  assign part2_io_mat_2_6 = io_matrix_2_6; // @[Distribution2.scala 76:18]
  assign part2_io_mat_2_7 = io_matrix_2_7; // @[Distribution2.scala 76:18]
  assign part2_io_mat_3_0 = io_matrix_3_0; // @[Distribution2.scala 76:18]
  assign part2_io_mat_3_1 = io_matrix_3_1; // @[Distribution2.scala 76:18]
  assign part2_io_mat_3_2 = io_matrix_3_2; // @[Distribution2.scala 76:18]
  assign part2_io_mat_3_3 = io_matrix_3_3; // @[Distribution2.scala 76:18]
  assign part2_io_mat_3_4 = io_matrix_3_4; // @[Distribution2.scala 76:18]
  assign part2_io_mat_3_5 = io_matrix_3_5; // @[Distribution2.scala 76:18]
  assign part2_io_mat_3_6 = io_matrix_3_6; // @[Distribution2.scala 76:18]
  assign part2_io_mat_3_7 = io_matrix_3_7; // @[Distribution2.scala 76:18]
  assign part2_io_mat_4_0 = io_matrix_4_0; // @[Distribution2.scala 76:18]
  assign part2_io_mat_4_1 = io_matrix_4_1; // @[Distribution2.scala 76:18]
  assign part2_io_mat_4_2 = io_matrix_4_2; // @[Distribution2.scala 76:18]
  assign part2_io_mat_4_3 = io_matrix_4_3; // @[Distribution2.scala 76:18]
  assign part2_io_mat_4_4 = io_matrix_4_4; // @[Distribution2.scala 76:18]
  assign part2_io_mat_4_5 = io_matrix_4_5; // @[Distribution2.scala 76:18]
  assign part2_io_mat_4_6 = io_matrix_4_6; // @[Distribution2.scala 76:18]
  assign part2_io_mat_4_7 = io_matrix_4_7; // @[Distribution2.scala 76:18]
  assign part2_io_mat_5_0 = io_matrix_5_0; // @[Distribution2.scala 76:18]
  assign part2_io_mat_5_1 = io_matrix_5_1; // @[Distribution2.scala 76:18]
  assign part2_io_mat_5_2 = io_matrix_5_2; // @[Distribution2.scala 76:18]
  assign part2_io_mat_5_3 = io_matrix_5_3; // @[Distribution2.scala 76:18]
  assign part2_io_mat_5_4 = io_matrix_5_4; // @[Distribution2.scala 76:18]
  assign part2_io_mat_5_5 = io_matrix_5_5; // @[Distribution2.scala 76:18]
  assign part2_io_mat_5_6 = io_matrix_5_6; // @[Distribution2.scala 76:18]
  assign part2_io_mat_5_7 = io_matrix_5_7; // @[Distribution2.scala 76:18]
  assign part2_io_mat_6_0 = io_matrix_6_0; // @[Distribution2.scala 76:18]
  assign part2_io_mat_6_1 = io_matrix_6_1; // @[Distribution2.scala 76:18]
  assign part2_io_mat_6_2 = io_matrix_6_2; // @[Distribution2.scala 76:18]
  assign part2_io_mat_6_3 = io_matrix_6_3; // @[Distribution2.scala 76:18]
  assign part2_io_mat_6_4 = io_matrix_6_4; // @[Distribution2.scala 76:18]
  assign part2_io_mat_6_5 = io_matrix_6_5; // @[Distribution2.scala 76:18]
  assign part2_io_mat_6_6 = io_matrix_6_6; // @[Distribution2.scala 76:18]
  assign part2_io_mat_6_7 = io_matrix_6_7; // @[Distribution2.scala 76:18]
  assign part2_io_mat_7_0 = io_matrix_7_0; // @[Distribution2.scala 76:18]
  assign part2_io_mat_7_1 = io_matrix_7_1; // @[Distribution2.scala 76:18]
  assign part2_io_mat_7_2 = io_matrix_7_2; // @[Distribution2.scala 76:18]
  assign part2_io_mat_7_3 = io_matrix_7_3; // @[Distribution2.scala 76:18]
  assign part2_io_mat_7_4 = io_matrix_7_4; // @[Distribution2.scala 76:18]
  assign part2_io_mat_7_5 = io_matrix_7_5; // @[Distribution2.scala 76:18]
  assign part2_io_mat_7_6 = io_matrix_7_6; // @[Distribution2.scala 76:18]
  assign part2_io_mat_7_7 = io_matrix_7_7; // @[Distribution2.scala 76:18]
  assign part3_clock = clock;
  assign part3_reset = reset;
  assign part3_io_IDex = 4'hf == io_s[3:0] ? Idex_15 : _GEN_369; // @[Distribution2.scala 92:{19,19}]
  assign part3_io_mat_0_0 = io_matrix_0_0; // @[Distribution2.scala 94:18]
  assign part3_io_mat_0_1 = io_matrix_0_1; // @[Distribution2.scala 94:18]
  assign part3_io_mat_0_2 = io_matrix_0_2; // @[Distribution2.scala 94:18]
  assign part3_io_mat_0_3 = io_matrix_0_3; // @[Distribution2.scala 94:18]
  assign part3_io_mat_0_4 = io_matrix_0_4; // @[Distribution2.scala 94:18]
  assign part3_io_mat_0_5 = io_matrix_0_5; // @[Distribution2.scala 94:18]
  assign part3_io_mat_0_6 = io_matrix_0_6; // @[Distribution2.scala 94:18]
  assign part3_io_mat_0_7 = io_matrix_0_7; // @[Distribution2.scala 94:18]
  assign part3_io_mat_1_0 = io_matrix_1_0; // @[Distribution2.scala 94:18]
  assign part3_io_mat_1_1 = io_matrix_1_1; // @[Distribution2.scala 94:18]
  assign part3_io_mat_1_2 = io_matrix_1_2; // @[Distribution2.scala 94:18]
  assign part3_io_mat_1_3 = io_matrix_1_3; // @[Distribution2.scala 94:18]
  assign part3_io_mat_1_4 = io_matrix_1_4; // @[Distribution2.scala 94:18]
  assign part3_io_mat_1_5 = io_matrix_1_5; // @[Distribution2.scala 94:18]
  assign part3_io_mat_1_6 = io_matrix_1_6; // @[Distribution2.scala 94:18]
  assign part3_io_mat_1_7 = io_matrix_1_7; // @[Distribution2.scala 94:18]
  assign part3_io_mat_2_0 = io_matrix_2_0; // @[Distribution2.scala 94:18]
  assign part3_io_mat_2_1 = io_matrix_2_1; // @[Distribution2.scala 94:18]
  assign part3_io_mat_2_2 = io_matrix_2_2; // @[Distribution2.scala 94:18]
  assign part3_io_mat_2_3 = io_matrix_2_3; // @[Distribution2.scala 94:18]
  assign part3_io_mat_2_4 = io_matrix_2_4; // @[Distribution2.scala 94:18]
  assign part3_io_mat_2_5 = io_matrix_2_5; // @[Distribution2.scala 94:18]
  assign part3_io_mat_2_6 = io_matrix_2_6; // @[Distribution2.scala 94:18]
  assign part3_io_mat_2_7 = io_matrix_2_7; // @[Distribution2.scala 94:18]
  assign part3_io_mat_3_0 = io_matrix_3_0; // @[Distribution2.scala 94:18]
  assign part3_io_mat_3_1 = io_matrix_3_1; // @[Distribution2.scala 94:18]
  assign part3_io_mat_3_2 = io_matrix_3_2; // @[Distribution2.scala 94:18]
  assign part3_io_mat_3_3 = io_matrix_3_3; // @[Distribution2.scala 94:18]
  assign part3_io_mat_3_4 = io_matrix_3_4; // @[Distribution2.scala 94:18]
  assign part3_io_mat_3_5 = io_matrix_3_5; // @[Distribution2.scala 94:18]
  assign part3_io_mat_3_6 = io_matrix_3_6; // @[Distribution2.scala 94:18]
  assign part3_io_mat_3_7 = io_matrix_3_7; // @[Distribution2.scala 94:18]
  assign part3_io_mat_4_0 = io_matrix_4_0; // @[Distribution2.scala 94:18]
  assign part3_io_mat_4_1 = io_matrix_4_1; // @[Distribution2.scala 94:18]
  assign part3_io_mat_4_2 = io_matrix_4_2; // @[Distribution2.scala 94:18]
  assign part3_io_mat_4_3 = io_matrix_4_3; // @[Distribution2.scala 94:18]
  assign part3_io_mat_4_4 = io_matrix_4_4; // @[Distribution2.scala 94:18]
  assign part3_io_mat_4_5 = io_matrix_4_5; // @[Distribution2.scala 94:18]
  assign part3_io_mat_4_6 = io_matrix_4_6; // @[Distribution2.scala 94:18]
  assign part3_io_mat_4_7 = io_matrix_4_7; // @[Distribution2.scala 94:18]
  assign part3_io_mat_5_0 = io_matrix_5_0; // @[Distribution2.scala 94:18]
  assign part3_io_mat_5_1 = io_matrix_5_1; // @[Distribution2.scala 94:18]
  assign part3_io_mat_5_2 = io_matrix_5_2; // @[Distribution2.scala 94:18]
  assign part3_io_mat_5_3 = io_matrix_5_3; // @[Distribution2.scala 94:18]
  assign part3_io_mat_5_4 = io_matrix_5_4; // @[Distribution2.scala 94:18]
  assign part3_io_mat_5_5 = io_matrix_5_5; // @[Distribution2.scala 94:18]
  assign part3_io_mat_5_6 = io_matrix_5_6; // @[Distribution2.scala 94:18]
  assign part3_io_mat_5_7 = io_matrix_5_7; // @[Distribution2.scala 94:18]
  assign part3_io_mat_6_0 = io_matrix_6_0; // @[Distribution2.scala 94:18]
  assign part3_io_mat_6_1 = io_matrix_6_1; // @[Distribution2.scala 94:18]
  assign part3_io_mat_6_2 = io_matrix_6_2; // @[Distribution2.scala 94:18]
  assign part3_io_mat_6_3 = io_matrix_6_3; // @[Distribution2.scala 94:18]
  assign part3_io_mat_6_4 = io_matrix_6_4; // @[Distribution2.scala 94:18]
  assign part3_io_mat_6_5 = io_matrix_6_5; // @[Distribution2.scala 94:18]
  assign part3_io_mat_6_6 = io_matrix_6_6; // @[Distribution2.scala 94:18]
  assign part3_io_mat_6_7 = io_matrix_6_7; // @[Distribution2.scala 94:18]
  assign part3_io_mat_7_0 = io_matrix_7_0; // @[Distribution2.scala 94:18]
  assign part3_io_mat_7_1 = io_matrix_7_1; // @[Distribution2.scala 94:18]
  assign part3_io_mat_7_2 = io_matrix_7_2; // @[Distribution2.scala 94:18]
  assign part3_io_mat_7_3 = io_matrix_7_3; // @[Distribution2.scala 94:18]
  assign part3_io_mat_7_4 = io_matrix_7_4; // @[Distribution2.scala 94:18]
  assign part3_io_mat_7_5 = io_matrix_7_5; // @[Distribution2.scala 94:18]
  assign part3_io_mat_7_6 = io_matrix_7_6; // @[Distribution2.scala 94:18]
  assign part3_io_mat_7_7 = io_matrix_7_7; // @[Distribution2.scala 94:18]
  assign part3_io_i_valid = part2_io_ProcessValid; // @[Distribution2.scala 95:22]
  assign Final_clock = clock;
  assign Final_reset = reset;
  assign Final_io_IDex = 4'hf == io_s[3:0] ? Idex_15 : _GEN_369; // @[Distribution2.scala 115:{27,27}]
  assign Final_io_PreMat_0_0 = part2_io_OutMat_0_0; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_0_1 = part2_io_OutMat_0_1; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_0_2 = part2_io_OutMat_0_2; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_0_3 = part2_io_OutMat_0_3; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_0_4 = part2_io_OutMat_0_4; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_0_5 = part2_io_OutMat_0_5; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_0_6 = part2_io_OutMat_0_6; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_0_7 = part2_io_OutMat_0_7; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_1_0 = part2_io_OutMat_1_0; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_1_1 = part2_io_OutMat_1_1; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_1_2 = part2_io_OutMat_1_2; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_1_3 = part2_io_OutMat_1_3; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_1_4 = part2_io_OutMat_1_4; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_1_5 = part2_io_OutMat_1_5; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_1_6 = part2_io_OutMat_1_6; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_1_7 = part2_io_OutMat_1_7; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_2_0 = part2_io_OutMat_2_0; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_2_1 = part2_io_OutMat_2_1; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_2_2 = part2_io_OutMat_2_2; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_2_3 = part2_io_OutMat_2_3; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_2_4 = part2_io_OutMat_2_4; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_2_5 = part2_io_OutMat_2_5; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_2_6 = part2_io_OutMat_2_6; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_2_7 = part2_io_OutMat_2_7; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_3_0 = part2_io_OutMat_3_0; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_3_1 = part2_io_OutMat_3_1; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_3_2 = part2_io_OutMat_3_2; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_3_3 = part2_io_OutMat_3_3; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_3_4 = part2_io_OutMat_3_4; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_3_5 = part2_io_OutMat_3_5; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_3_6 = part2_io_OutMat_3_6; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_3_7 = part2_io_OutMat_3_7; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_4_0 = part2_io_OutMat_4_0; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_4_1 = part2_io_OutMat_4_1; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_4_2 = part2_io_OutMat_4_2; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_4_3 = part2_io_OutMat_4_3; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_4_4 = part2_io_OutMat_4_4; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_4_5 = part2_io_OutMat_4_5; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_4_6 = part2_io_OutMat_4_6; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_4_7 = part2_io_OutMat_4_7; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_5_0 = part2_io_OutMat_5_0; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_5_1 = part2_io_OutMat_5_1; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_5_2 = part2_io_OutMat_5_2; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_5_3 = part2_io_OutMat_5_3; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_5_4 = part2_io_OutMat_5_4; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_5_5 = part2_io_OutMat_5_5; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_5_6 = part2_io_OutMat_5_6; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_5_7 = part2_io_OutMat_5_7; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_6_0 = part2_io_OutMat_6_0; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_6_1 = part2_io_OutMat_6_1; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_6_2 = part2_io_OutMat_6_2; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_6_3 = part2_io_OutMat_6_3; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_6_4 = part2_io_OutMat_6_4; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_6_5 = part2_io_OutMat_6_5; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_6_6 = part2_io_OutMat_6_6; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_6_7 = part2_io_OutMat_6_7; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_7_0 = part2_io_OutMat_7_0; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_7_1 = part2_io_OutMat_7_1; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_7_2 = part2_io_OutMat_7_2; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_7_3 = part2_io_OutMat_7_3; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_7_4 = part2_io_OutMat_7_4; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_7_5 = part2_io_OutMat_7_5; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_7_6 = part2_io_OutMat_7_6; // @[Distribution2.scala 117:29]
  assign Final_io_PreMat_7_7 = part2_io_OutMat_7_7; // @[Distribution2.scala 117:29]
  assign Final_io_lastMat_0_0 = part3_io_Omat_0_0; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_0_1 = part3_io_Omat_0_1; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_0_2 = part3_io_Omat_0_2; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_0_3 = part3_io_Omat_0_3; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_0_4 = part3_io_Omat_0_4; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_0_5 = part3_io_Omat_0_5; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_0_6 = part3_io_Omat_0_6; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_0_7 = part3_io_Omat_0_7; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_1_0 = part3_io_Omat_1_0; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_1_1 = part3_io_Omat_1_1; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_1_2 = part3_io_Omat_1_2; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_1_3 = part3_io_Omat_1_3; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_1_4 = part3_io_Omat_1_4; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_1_5 = part3_io_Omat_1_5; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_1_6 = part3_io_Omat_1_6; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_1_7 = part3_io_Omat_1_7; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_2_0 = part3_io_Omat_2_0; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_2_1 = part3_io_Omat_2_1; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_2_2 = part3_io_Omat_2_2; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_2_3 = part3_io_Omat_2_3; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_2_4 = part3_io_Omat_2_4; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_2_5 = part3_io_Omat_2_5; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_2_6 = part3_io_Omat_2_6; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_2_7 = part3_io_Omat_2_7; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_3_0 = part3_io_Omat_3_0; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_3_1 = part3_io_Omat_3_1; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_3_2 = part3_io_Omat_3_2; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_3_3 = part3_io_Omat_3_3; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_3_4 = part3_io_Omat_3_4; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_3_5 = part3_io_Omat_3_5; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_3_6 = part3_io_Omat_3_6; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_3_7 = part3_io_Omat_3_7; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_4_0 = part3_io_Omat_4_0; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_4_1 = part3_io_Omat_4_1; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_4_2 = part3_io_Omat_4_2; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_4_3 = part3_io_Omat_4_3; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_4_4 = part3_io_Omat_4_4; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_4_5 = part3_io_Omat_4_5; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_4_6 = part3_io_Omat_4_6; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_4_7 = part3_io_Omat_4_7; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_5_0 = part3_io_Omat_5_0; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_5_1 = part3_io_Omat_5_1; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_5_2 = part3_io_Omat_5_2; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_5_3 = part3_io_Omat_5_3; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_5_4 = part3_io_Omat_5_4; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_5_5 = part3_io_Omat_5_5; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_5_6 = part3_io_Omat_5_6; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_5_7 = part3_io_Omat_5_7; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_6_0 = part3_io_Omat_6_0; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_6_1 = part3_io_Omat_6_1; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_6_2 = part3_io_Omat_6_2; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_6_3 = part3_io_Omat_6_3; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_6_4 = part3_io_Omat_6_4; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_6_5 = part3_io_Omat_6_5; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_6_6 = part3_io_Omat_6_6; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_6_7 = part3_io_Omat_6_7; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_7_0 = part3_io_Omat_7_0; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_7_1 = part3_io_Omat_7_1; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_7_2 = part3_io_Omat_7_2; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_7_3 = part3_io_Omat_7_3; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_7_4 = part3_io_Omat_7_4; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_7_5 = part3_io_Omat_7_5; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_7_6 = part3_io_Omat_7_6; // @[Distribution2.scala 119:30]
  assign Final_io_lastMat_7_7 = part3_io_Omat_7_7; // @[Distribution2.scala 119:30]
  assign Final_io_valid = part3_io_valid; // @[Distribution2.scala 118:28]
  always @(posedge clock) begin
    if (reset) begin // @[Distribution2.scala 22:20]
      i <= 32'h0; // @[Distribution2.scala 22:20]
    end else if (io_valid) begin // @[Distribution2.scala 237:20]
      if (i < 32'h7 & _T_17) begin // @[Distribution2.scala 238:69]
        i <= _i_T_1; // @[Distribution2.scala 239:11]
      end
    end
    if (reset) begin // @[Distribution2.scala 23:20]
      j <= 32'h0; // @[Distribution2.scala 23:20]
    end else if (io_valid) begin // @[Distribution2.scala 237:20]
      if (i <= 32'h7 & j < 32'h7) begin // @[Distribution2.scala 241:68]
        j <= _j_T_1; // @[Distribution2.scala 242:11]
      end else if (!(_complete_T_2)) begin // @[Distribution2.scala 243:75]
        j <= 32'h0; // @[Distribution2.scala 246:11]
      end
    end
    if (reset) begin // @[Distribution2.scala 24:24]
      count <= 32'h0; // @[Distribution2.scala 24:24]
    end else if (io_valid) begin // @[Distribution2.scala 60:20]
      if (_T_2 & (i != 32'h7 | j != 32'h7)) begin // @[Distribution2.scala 61:103]
        count <= _count_T_1; // @[Distribution2.scala 62:15]
      end
    end
    if (reset) begin // @[Distribution2.scala 25:23]
      Idex_0 <= 32'h0; // @[Distribution2.scala 25:23]
    end else if (io_valid) begin // @[Distribution2.scala 60:20]
      if (_T_2 & (i != 32'h7 | j != 32'h7)) begin // @[Distribution2.scala 61:103]
        Idex_0 <= _GEN_129;
      end else if (_T_2 & i == 32'h7 & j == 32'h7) begin // @[Distribution2.scala 65:106]
        Idex_0 <= _GEN_129;
      end
    end
    if (reset) begin // @[Distribution2.scala 25:23]
      Idex_1 <= 32'h0; // @[Distribution2.scala 25:23]
    end else if (io_valid) begin // @[Distribution2.scala 60:20]
      if (_T_2 & (i != 32'h7 | j != 32'h7)) begin // @[Distribution2.scala 61:103]
        Idex_1 <= _GEN_130;
      end else if (_T_2 & i == 32'h7 & j == 32'h7) begin // @[Distribution2.scala 65:106]
        Idex_1 <= _GEN_130;
      end
    end
    if (reset) begin // @[Distribution2.scala 25:23]
      Idex_2 <= 32'h0; // @[Distribution2.scala 25:23]
    end else if (io_valid) begin // @[Distribution2.scala 60:20]
      if (_T_2 & (i != 32'h7 | j != 32'h7)) begin // @[Distribution2.scala 61:103]
        Idex_2 <= _GEN_131;
      end else if (_T_2 & i == 32'h7 & j == 32'h7) begin // @[Distribution2.scala 65:106]
        Idex_2 <= _GEN_131;
      end
    end
    if (reset) begin // @[Distribution2.scala 25:23]
      Idex_3 <= 32'h0; // @[Distribution2.scala 25:23]
    end else if (io_valid) begin // @[Distribution2.scala 60:20]
      if (_T_2 & (i != 32'h7 | j != 32'h7)) begin // @[Distribution2.scala 61:103]
        Idex_3 <= _GEN_132;
      end else if (_T_2 & i == 32'h7 & j == 32'h7) begin // @[Distribution2.scala 65:106]
        Idex_3 <= _GEN_132;
      end
    end
    if (reset) begin // @[Distribution2.scala 25:23]
      Idex_4 <= 32'h0; // @[Distribution2.scala 25:23]
    end else if (io_valid) begin // @[Distribution2.scala 60:20]
      if (_T_2 & (i != 32'h7 | j != 32'h7)) begin // @[Distribution2.scala 61:103]
        Idex_4 <= _GEN_133;
      end else if (_T_2 & i == 32'h7 & j == 32'h7) begin // @[Distribution2.scala 65:106]
        Idex_4 <= _GEN_133;
      end
    end
    if (reset) begin // @[Distribution2.scala 25:23]
      Idex_5 <= 32'h0; // @[Distribution2.scala 25:23]
    end else if (io_valid) begin // @[Distribution2.scala 60:20]
      if (_T_2 & (i != 32'h7 | j != 32'h7)) begin // @[Distribution2.scala 61:103]
        Idex_5 <= _GEN_134;
      end else if (_T_2 & i == 32'h7 & j == 32'h7) begin // @[Distribution2.scala 65:106]
        Idex_5 <= _GEN_134;
      end
    end
    if (reset) begin // @[Distribution2.scala 25:23]
      Idex_6 <= 32'h0; // @[Distribution2.scala 25:23]
    end else if (io_valid) begin // @[Distribution2.scala 60:20]
      if (_T_2 & (i != 32'h7 | j != 32'h7)) begin // @[Distribution2.scala 61:103]
        Idex_6 <= _GEN_135;
      end else if (_T_2 & i == 32'h7 & j == 32'h7) begin // @[Distribution2.scala 65:106]
        Idex_6 <= _GEN_135;
      end
    end
    if (reset) begin // @[Distribution2.scala 25:23]
      Idex_7 <= 32'h0; // @[Distribution2.scala 25:23]
    end else if (io_valid) begin // @[Distribution2.scala 60:20]
      if (_T_2 & (i != 32'h7 | j != 32'h7)) begin // @[Distribution2.scala 61:103]
        Idex_7 <= _GEN_136;
      end else if (_T_2 & i == 32'h7 & j == 32'h7) begin // @[Distribution2.scala 65:106]
        Idex_7 <= _GEN_136;
      end
    end
    if (reset) begin // @[Distribution2.scala 25:23]
      Idex_8 <= 32'h0; // @[Distribution2.scala 25:23]
    end else if (io_valid) begin // @[Distribution2.scala 60:20]
      if (_T_2 & (i != 32'h7 | j != 32'h7)) begin // @[Distribution2.scala 61:103]
        Idex_8 <= _GEN_137;
      end else if (_T_2 & i == 32'h7 & j == 32'h7) begin // @[Distribution2.scala 65:106]
        Idex_8 <= _GEN_137;
      end
    end
    if (reset) begin // @[Distribution2.scala 25:23]
      Idex_9 <= 32'h0; // @[Distribution2.scala 25:23]
    end else if (io_valid) begin // @[Distribution2.scala 60:20]
      if (_T_2 & (i != 32'h7 | j != 32'h7)) begin // @[Distribution2.scala 61:103]
        Idex_9 <= _GEN_138;
      end else if (_T_2 & i == 32'h7 & j == 32'h7) begin // @[Distribution2.scala 65:106]
        Idex_9 <= _GEN_138;
      end
    end
    if (reset) begin // @[Distribution2.scala 25:23]
      Idex_10 <= 32'h0; // @[Distribution2.scala 25:23]
    end else if (io_valid) begin // @[Distribution2.scala 60:20]
      if (_T_2 & (i != 32'h7 | j != 32'h7)) begin // @[Distribution2.scala 61:103]
        Idex_10 <= _GEN_139;
      end else if (_T_2 & i == 32'h7 & j == 32'h7) begin // @[Distribution2.scala 65:106]
        Idex_10 <= _GEN_139;
      end
    end
    if (reset) begin // @[Distribution2.scala 25:23]
      Idex_11 <= 32'h0; // @[Distribution2.scala 25:23]
    end else if (io_valid) begin // @[Distribution2.scala 60:20]
      if (_T_2 & (i != 32'h7 | j != 32'h7)) begin // @[Distribution2.scala 61:103]
        Idex_11 <= _GEN_140;
      end else if (_T_2 & i == 32'h7 & j == 32'h7) begin // @[Distribution2.scala 65:106]
        Idex_11 <= _GEN_140;
      end
    end
    if (reset) begin // @[Distribution2.scala 25:23]
      Idex_12 <= 32'h0; // @[Distribution2.scala 25:23]
    end else if (io_valid) begin // @[Distribution2.scala 60:20]
      if (_T_2 & (i != 32'h7 | j != 32'h7)) begin // @[Distribution2.scala 61:103]
        Idex_12 <= _GEN_141;
      end else if (_T_2 & i == 32'h7 & j == 32'h7) begin // @[Distribution2.scala 65:106]
        Idex_12 <= _GEN_141;
      end
    end
    if (reset) begin // @[Distribution2.scala 25:23]
      Idex_13 <= 32'h0; // @[Distribution2.scala 25:23]
    end else if (io_valid) begin // @[Distribution2.scala 60:20]
      if (_T_2 & (i != 32'h7 | j != 32'h7)) begin // @[Distribution2.scala 61:103]
        Idex_13 <= _GEN_142;
      end else if (_T_2 & i == 32'h7 & j == 32'h7) begin // @[Distribution2.scala 65:106]
        Idex_13 <= _GEN_142;
      end
    end
    if (reset) begin // @[Distribution2.scala 25:23]
      Idex_14 <= 32'h0; // @[Distribution2.scala 25:23]
    end else if (io_valid) begin // @[Distribution2.scala 60:20]
      if (_T_2 & (i != 32'h7 | j != 32'h7)) begin // @[Distribution2.scala 61:103]
        Idex_14 <= _GEN_143;
      end else if (_T_2 & i == 32'h7 & j == 32'h7) begin // @[Distribution2.scala 65:106]
        Idex_14 <= _GEN_143;
      end
    end
    if (reset) begin // @[Distribution2.scala 25:23]
      Idex_15 <= 32'h0; // @[Distribution2.scala 25:23]
    end else if (io_valid) begin // @[Distribution2.scala 60:20]
      if (_T_2 & (i != 32'h7 | j != 32'h7)) begin // @[Distribution2.scala 61:103]
        Idex_15 <= _GEN_144;
      end else if (_T_2 & i == 32'h7 & j == 32'h7) begin // @[Distribution2.scala 65:106]
        Idex_15 <= _GEN_144;
      end
    end
    if (reset) begin // @[Distribution2.scala 26:23]
      Jdex_0 <= 32'h0; // @[Distribution2.scala 26:23]
    end else if (io_valid) begin // @[Distribution2.scala 60:20]
      if (_T_2 & (i != 32'h7 | j != 32'h7)) begin // @[Distribution2.scala 61:103]
        Jdex_0 <= _GEN_145;
      end else if (_T_2 & i == 32'h7 & j == 32'h7) begin // @[Distribution2.scala 65:106]
        Jdex_0 <= _GEN_145;
      end
    end
    if (reset) begin // @[Distribution2.scala 26:23]
      Jdex_1 <= 32'h0; // @[Distribution2.scala 26:23]
    end else if (io_valid) begin // @[Distribution2.scala 60:20]
      if (_T_2 & (i != 32'h7 | j != 32'h7)) begin // @[Distribution2.scala 61:103]
        Jdex_1 <= _GEN_146;
      end else if (_T_2 & i == 32'h7 & j == 32'h7) begin // @[Distribution2.scala 65:106]
        Jdex_1 <= _GEN_146;
      end
    end
    if (reset) begin // @[Distribution2.scala 26:23]
      Jdex_2 <= 32'h0; // @[Distribution2.scala 26:23]
    end else if (io_valid) begin // @[Distribution2.scala 60:20]
      if (_T_2 & (i != 32'h7 | j != 32'h7)) begin // @[Distribution2.scala 61:103]
        Jdex_2 <= _GEN_147;
      end else if (_T_2 & i == 32'h7 & j == 32'h7) begin // @[Distribution2.scala 65:106]
        Jdex_2 <= _GEN_147;
      end
    end
    if (reset) begin // @[Distribution2.scala 26:23]
      Jdex_3 <= 32'h0; // @[Distribution2.scala 26:23]
    end else if (io_valid) begin // @[Distribution2.scala 60:20]
      if (_T_2 & (i != 32'h7 | j != 32'h7)) begin // @[Distribution2.scala 61:103]
        Jdex_3 <= _GEN_148;
      end else if (_T_2 & i == 32'h7 & j == 32'h7) begin // @[Distribution2.scala 65:106]
        Jdex_3 <= _GEN_148;
      end
    end
    if (reset) begin // @[Distribution2.scala 26:23]
      Jdex_4 <= 32'h0; // @[Distribution2.scala 26:23]
    end else if (io_valid) begin // @[Distribution2.scala 60:20]
      if (_T_2 & (i != 32'h7 | j != 32'h7)) begin // @[Distribution2.scala 61:103]
        Jdex_4 <= _GEN_149;
      end else if (_T_2 & i == 32'h7 & j == 32'h7) begin // @[Distribution2.scala 65:106]
        Jdex_4 <= _GEN_149;
      end
    end
    if (reset) begin // @[Distribution2.scala 26:23]
      Jdex_5 <= 32'h0; // @[Distribution2.scala 26:23]
    end else if (io_valid) begin // @[Distribution2.scala 60:20]
      if (_T_2 & (i != 32'h7 | j != 32'h7)) begin // @[Distribution2.scala 61:103]
        Jdex_5 <= _GEN_150;
      end else if (_T_2 & i == 32'h7 & j == 32'h7) begin // @[Distribution2.scala 65:106]
        Jdex_5 <= _GEN_150;
      end
    end
    if (reset) begin // @[Distribution2.scala 26:23]
      Jdex_6 <= 32'h0; // @[Distribution2.scala 26:23]
    end else if (io_valid) begin // @[Distribution2.scala 60:20]
      if (_T_2 & (i != 32'h7 | j != 32'h7)) begin // @[Distribution2.scala 61:103]
        Jdex_6 <= _GEN_151;
      end else if (_T_2 & i == 32'h7 & j == 32'h7) begin // @[Distribution2.scala 65:106]
        Jdex_6 <= _GEN_151;
      end
    end
    if (reset) begin // @[Distribution2.scala 26:23]
      Jdex_7 <= 32'h0; // @[Distribution2.scala 26:23]
    end else if (io_valid) begin // @[Distribution2.scala 60:20]
      if (_T_2 & (i != 32'h7 | j != 32'h7)) begin // @[Distribution2.scala 61:103]
        Jdex_7 <= _GEN_152;
      end else if (_T_2 & i == 32'h7 & j == 32'h7) begin // @[Distribution2.scala 65:106]
        Jdex_7 <= _GEN_152;
      end
    end
    if (reset) begin // @[Distribution2.scala 26:23]
      Jdex_8 <= 32'h0; // @[Distribution2.scala 26:23]
    end else if (io_valid) begin // @[Distribution2.scala 60:20]
      if (_T_2 & (i != 32'h7 | j != 32'h7)) begin // @[Distribution2.scala 61:103]
        Jdex_8 <= _GEN_153;
      end else if (_T_2 & i == 32'h7 & j == 32'h7) begin // @[Distribution2.scala 65:106]
        Jdex_8 <= _GEN_153;
      end
    end
    if (reset) begin // @[Distribution2.scala 26:23]
      Jdex_9 <= 32'h0; // @[Distribution2.scala 26:23]
    end else if (io_valid) begin // @[Distribution2.scala 60:20]
      if (_T_2 & (i != 32'h7 | j != 32'h7)) begin // @[Distribution2.scala 61:103]
        Jdex_9 <= _GEN_154;
      end else if (_T_2 & i == 32'h7 & j == 32'h7) begin // @[Distribution2.scala 65:106]
        Jdex_9 <= _GEN_154;
      end
    end
    if (reset) begin // @[Distribution2.scala 26:23]
      Jdex_10 <= 32'h0; // @[Distribution2.scala 26:23]
    end else if (io_valid) begin // @[Distribution2.scala 60:20]
      if (_T_2 & (i != 32'h7 | j != 32'h7)) begin // @[Distribution2.scala 61:103]
        Jdex_10 <= _GEN_155;
      end else if (_T_2 & i == 32'h7 & j == 32'h7) begin // @[Distribution2.scala 65:106]
        Jdex_10 <= _GEN_155;
      end
    end
    if (reset) begin // @[Distribution2.scala 26:23]
      Jdex_11 <= 32'h0; // @[Distribution2.scala 26:23]
    end else if (io_valid) begin // @[Distribution2.scala 60:20]
      if (_T_2 & (i != 32'h7 | j != 32'h7)) begin // @[Distribution2.scala 61:103]
        Jdex_11 <= _GEN_156;
      end else if (_T_2 & i == 32'h7 & j == 32'h7) begin // @[Distribution2.scala 65:106]
        Jdex_11 <= _GEN_156;
      end
    end
    if (reset) begin // @[Distribution2.scala 26:23]
      Jdex_12 <= 32'h0; // @[Distribution2.scala 26:23]
    end else if (io_valid) begin // @[Distribution2.scala 60:20]
      if (_T_2 & (i != 32'h7 | j != 32'h7)) begin // @[Distribution2.scala 61:103]
        Jdex_12 <= _GEN_157;
      end else if (_T_2 & i == 32'h7 & j == 32'h7) begin // @[Distribution2.scala 65:106]
        Jdex_12 <= _GEN_157;
      end
    end
    if (reset) begin // @[Distribution2.scala 26:23]
      Jdex_13 <= 32'h0; // @[Distribution2.scala 26:23]
    end else if (io_valid) begin // @[Distribution2.scala 60:20]
      if (_T_2 & (i != 32'h7 | j != 32'h7)) begin // @[Distribution2.scala 61:103]
        Jdex_13 <= _GEN_158;
      end else if (_T_2 & i == 32'h7 & j == 32'h7) begin // @[Distribution2.scala 65:106]
        Jdex_13 <= _GEN_158;
      end
    end
    if (reset) begin // @[Distribution2.scala 26:23]
      Jdex_14 <= 32'h0; // @[Distribution2.scala 26:23]
    end else if (io_valid) begin // @[Distribution2.scala 60:20]
      if (_T_2 & (i != 32'h7 | j != 32'h7)) begin // @[Distribution2.scala 61:103]
        Jdex_14 <= _GEN_159;
      end else if (_T_2 & i == 32'h7 & j == 32'h7) begin // @[Distribution2.scala 65:106]
        Jdex_14 <= _GEN_159;
      end
    end
    if (reset) begin // @[Distribution2.scala 26:23]
      Jdex_15 <= 32'h0; // @[Distribution2.scala 26:23]
    end else if (io_valid) begin // @[Distribution2.scala 60:20]
      if (_T_2 & (i != 32'h7 | j != 32'h7)) begin // @[Distribution2.scala 61:103]
        Jdex_15 <= _GEN_160;
      end else if (_T_2 & i == 32'h7 & j == 32'h7) begin // @[Distribution2.scala 65:106]
        Jdex_15 <= _GEN_160;
      end
    end
    complete <= _T_15 & _T_17; // @[Distribution2.scala 78:55]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  i = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  j = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  count = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  Idex_0 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  Idex_1 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  Idex_2 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  Idex_3 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  Idex_4 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  Idex_5 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  Idex_6 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  Idex_7 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  Idex_8 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  Idex_9 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  Idex_10 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  Idex_11 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  Idex_12 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  Idex_13 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  Idex_14 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  Idex_15 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  Jdex_0 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  Jdex_1 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  Jdex_2 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  Jdex_3 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  Jdex_4 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  Jdex_5 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  Jdex_6 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  Jdex_7 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  Jdex_8 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  Jdex_9 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  Jdex_10 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  Jdex_11 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  Jdex_12 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  Jdex_13 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  Jdex_14 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  Jdex_15 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  complete = _RAND_35[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PathFinder(
  input         clock,
  input         reset,
  input  [15:0] io_Stationary_matrix_0_0,
  input  [15:0] io_Stationary_matrix_0_1,
  input  [15:0] io_Stationary_matrix_0_2,
  input  [15:0] io_Stationary_matrix_0_3,
  input  [15:0] io_Stationary_matrix_0_4,
  input  [15:0] io_Stationary_matrix_0_5,
  input  [15:0] io_Stationary_matrix_0_6,
  input  [15:0] io_Stationary_matrix_0_7,
  input  [15:0] io_Stationary_matrix_1_0,
  input  [15:0] io_Stationary_matrix_1_1,
  input  [15:0] io_Stationary_matrix_1_2,
  input  [15:0] io_Stationary_matrix_1_3,
  input  [15:0] io_Stationary_matrix_1_4,
  input  [15:0] io_Stationary_matrix_1_5,
  input  [15:0] io_Stationary_matrix_1_6,
  input  [15:0] io_Stationary_matrix_1_7,
  input  [15:0] io_Stationary_matrix_2_0,
  input  [15:0] io_Stationary_matrix_2_1,
  input  [15:0] io_Stationary_matrix_2_2,
  input  [15:0] io_Stationary_matrix_2_3,
  input  [15:0] io_Stationary_matrix_2_4,
  input  [15:0] io_Stationary_matrix_2_5,
  input  [15:0] io_Stationary_matrix_2_6,
  input  [15:0] io_Stationary_matrix_2_7,
  input  [15:0] io_Stationary_matrix_3_0,
  input  [15:0] io_Stationary_matrix_3_1,
  input  [15:0] io_Stationary_matrix_3_2,
  input  [15:0] io_Stationary_matrix_3_3,
  input  [15:0] io_Stationary_matrix_3_4,
  input  [15:0] io_Stationary_matrix_3_5,
  input  [15:0] io_Stationary_matrix_3_6,
  input  [15:0] io_Stationary_matrix_3_7,
  input  [15:0] io_Stationary_matrix_4_0,
  input  [15:0] io_Stationary_matrix_4_1,
  input  [15:0] io_Stationary_matrix_4_2,
  input  [15:0] io_Stationary_matrix_4_3,
  input  [15:0] io_Stationary_matrix_4_4,
  input  [15:0] io_Stationary_matrix_4_5,
  input  [15:0] io_Stationary_matrix_4_6,
  input  [15:0] io_Stationary_matrix_4_7,
  input  [15:0] io_Stationary_matrix_5_0,
  input  [15:0] io_Stationary_matrix_5_1,
  input  [15:0] io_Stationary_matrix_5_2,
  input  [15:0] io_Stationary_matrix_5_3,
  input  [15:0] io_Stationary_matrix_5_4,
  input  [15:0] io_Stationary_matrix_5_5,
  input  [15:0] io_Stationary_matrix_5_6,
  input  [15:0] io_Stationary_matrix_5_7,
  input  [15:0] io_Stationary_matrix_6_0,
  input  [15:0] io_Stationary_matrix_6_1,
  input  [15:0] io_Stationary_matrix_6_2,
  input  [15:0] io_Stationary_matrix_6_3,
  input  [15:0] io_Stationary_matrix_6_4,
  input  [15:0] io_Stationary_matrix_6_5,
  input  [15:0] io_Stationary_matrix_6_6,
  input  [15:0] io_Stationary_matrix_6_7,
  input  [15:0] io_Stationary_matrix_7_0,
  input  [15:0] io_Stationary_matrix_7_1,
  input  [15:0] io_Stationary_matrix_7_2,
  input  [15:0] io_Stationary_matrix_7_3,
  input  [15:0] io_Stationary_matrix_7_4,
  input  [15:0] io_Stationary_matrix_7_5,
  input  [15:0] io_Stationary_matrix_7_6,
  input  [15:0] io_Stationary_matrix_7_7,
  input  [15:0] io_Streaming_matrix_0,
  input  [15:0] io_Streaming_matrix_1,
  input  [15:0] io_Streaming_matrix_2,
  input  [15:0] io_Streaming_matrix_3,
  input  [15:0] io_Streaming_matrix_4,
  input  [15:0] io_Streaming_matrix_5,
  input  [15:0] io_Streaming_matrix_6,
  input  [15:0] io_Streaming_matrix_7,
  output [3:0]  io_i_mux_bus_0,
  output [3:0]  io_i_mux_bus_1,
  output [3:0]  io_i_mux_bus_2,
  output [3:0]  io_i_mux_bus_3,
  output [15:0] io_Source_0,
  output [15:0] io_Source_1,
  output [15:0] io_Source_2,
  output [15:0] io_Source_3,
  output        io_PF_Valid,
  input  [31:0] io_NoDPE,
  input         io_DataValid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  myMuxes_clock; // @[PathFinder.scala 25:23]
  wire  myMuxes_reset; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_0_0; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_0_1; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_0_2; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_0_3; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_0_4; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_0_5; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_0_6; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_0_7; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_1_0; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_1_1; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_1_2; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_1_3; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_1_4; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_1_5; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_1_6; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_1_7; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_2_0; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_2_1; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_2_2; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_2_3; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_2_4; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_2_5; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_2_6; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_2_7; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_3_0; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_3_1; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_3_2; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_3_3; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_3_4; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_3_5; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_3_6; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_3_7; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_4_0; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_4_1; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_4_2; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_4_3; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_4_4; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_4_5; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_4_6; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_4_7; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_5_0; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_5_1; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_5_2; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_5_3; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_5_4; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_5_5; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_5_6; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_5_7; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_6_0; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_6_1; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_6_2; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_6_3; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_6_4; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_6_5; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_6_6; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_6_7; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_7_0; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_7_1; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_7_2; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_7_3; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_7_4; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_7_5; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_7_6; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat1_7_7; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat2_0; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat2_1; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat2_2; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat2_3; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat2_4; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat2_5; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat2_6; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_mat2_7; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_0_0; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_0_1; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_0_2; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_0_3; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_0_4; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_0_5; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_0_6; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_0_7; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_1_0; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_1_1; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_1_2; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_1_3; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_1_4; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_1_5; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_1_6; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_1_7; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_2_0; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_2_1; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_2_2; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_2_3; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_2_4; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_2_5; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_2_6; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_2_7; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_3_0; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_3_1; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_3_2; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_3_3; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_3_4; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_3_5; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_3_6; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_3_7; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_4_0; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_4_1; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_4_2; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_4_3; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_4_4; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_4_5; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_4_6; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_4_7; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_5_0; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_5_1; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_5_2; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_5_3; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_5_4; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_5_5; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_5_6; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_5_7; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_6_0; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_6_1; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_6_2; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_6_3; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_6_4; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_6_5; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_6_6; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_6_7; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_7_0; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_7_1; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_7_2; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_7_3; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_7_4; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_7_5; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_7_6; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix1_7_7; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix2_0; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix2_1; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix2_2; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix2_3; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix2_4; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix2_5; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix2_6; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_counterMatrix2_7; // @[PathFinder.scala 25:23]
  wire [3:0] myMuxes_io_i_mux_bus_0; // @[PathFinder.scala 25:23]
  wire [3:0] myMuxes_io_i_mux_bus_1; // @[PathFinder.scala 25:23]
  wire [3:0] myMuxes_io_i_mux_bus_2; // @[PathFinder.scala 25:23]
  wire [3:0] myMuxes_io_i_mux_bus_3; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_Source_0; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_Source_1; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_Source_2; // @[PathFinder.scala 25:23]
  wire [15:0] myMuxes_io_Source_3; // @[PathFinder.scala 25:23]
  wire  myMuxes_io_valid; // @[PathFinder.scala 25:23]
  wire  myCounter_clock; // @[PathFinder.scala 31:25]
  wire  myCounter_reset; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_0_0; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_0_1; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_0_2; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_0_3; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_0_4; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_0_5; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_0_6; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_0_7; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_1_0; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_1_1; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_1_2; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_1_3; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_1_4; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_1_5; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_1_6; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_1_7; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_2_0; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_2_1; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_2_2; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_2_3; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_2_4; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_2_5; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_2_6; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_2_7; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_3_0; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_3_1; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_3_2; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_3_3; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_3_4; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_3_5; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_3_6; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_3_7; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_4_0; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_4_1; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_4_2; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_4_3; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_4_4; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_4_5; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_4_6; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_4_7; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_5_0; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_5_1; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_5_2; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_5_3; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_5_4; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_5_5; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_5_6; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_5_7; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_6_0; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_6_1; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_6_2; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_6_3; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_6_4; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_6_5; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_6_6; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_6_7; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_7_0; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_7_1; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_7_2; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_7_3; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_7_4; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_7_5; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_7_6; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Stationary_matrix_7_7; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Streaming_matrix_0; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Streaming_matrix_1; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Streaming_matrix_2; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Streaming_matrix_3; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Streaming_matrix_4; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Streaming_matrix_5; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Streaming_matrix_6; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_Streaming_matrix_7; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_0_0; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_0_1; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_0_2; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_0_3; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_0_4; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_0_5; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_0_6; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_0_7; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_1_0; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_1_1; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_1_2; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_1_3; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_1_4; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_1_5; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_1_6; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_1_7; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_2_0; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_2_1; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_2_2; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_2_3; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_2_4; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_2_5; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_2_6; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_2_7; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_3_0; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_3_1; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_3_2; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_3_3; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_3_4; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_3_5; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_3_6; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_3_7; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_4_0; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_4_1; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_4_2; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_4_3; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_4_4; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_4_5; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_4_6; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_4_7; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_5_0; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_5_1; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_5_2; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_5_3; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_5_4; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_5_5; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_5_6; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_5_7; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_6_0; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_6_1; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_6_2; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_6_3; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_6_4; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_6_5; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_6_6; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_6_7; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_7_0; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_7_1; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_7_2; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_7_3; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_7_4; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_7_5; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_7_6; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix1_bits_7_7; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix2_bits_0; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix2_bits_1; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix2_bits_2; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix2_bits_3; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix2_bits_4; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix2_bits_5; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix2_bits_6; // @[PathFinder.scala 31:25]
  wire [15:0] myCounter_io_counterMatrix2_bits_7; // @[PathFinder.scala 31:25]
  wire  myCounter_io_valid; // @[PathFinder.scala 31:25]
  wire  myCounter_io_start; // @[PathFinder.scala 31:25]
  wire  Distribution_clock; // @[PathFinder.scala 50:28]
  wire  Distribution_reset; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_0_0; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_0_1; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_0_2; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_0_3; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_0_4; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_0_5; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_0_6; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_0_7; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_1_0; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_1_1; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_1_2; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_1_3; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_1_4; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_1_5; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_1_6; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_1_7; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_2_0; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_2_1; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_2_2; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_2_3; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_2_4; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_2_5; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_2_6; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_2_7; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_3_0; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_3_1; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_3_2; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_3_3; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_3_4; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_3_5; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_3_6; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_3_7; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_4_0; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_4_1; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_4_2; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_4_3; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_4_4; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_4_5; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_4_6; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_4_7; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_5_0; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_5_1; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_5_2; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_5_3; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_5_4; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_5_5; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_5_6; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_5_7; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_6_0; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_6_1; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_6_2; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_6_3; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_6_4; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_6_5; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_6_6; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_6_7; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_7_0; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_7_1; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_7_2; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_7_3; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_7_4; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_7_5; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_7_6; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_matrix_7_7; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_s; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_0_0; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_0_1; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_0_2; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_0_3; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_0_4; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_0_5; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_0_6; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_0_7; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_1_0; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_1_1; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_1_2; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_1_3; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_1_4; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_1_5; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_1_6; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_1_7; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_2_0; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_2_1; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_2_2; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_2_3; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_2_4; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_2_5; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_2_6; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_2_7; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_3_0; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_3_1; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_3_2; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_3_3; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_3_4; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_3_5; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_3_6; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_3_7; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_4_0; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_4_1; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_4_2; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_4_3; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_4_4; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_4_5; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_4_6; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_4_7; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_5_0; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_5_1; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_5_2; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_5_3; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_5_4; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_5_5; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_5_6; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_5_7; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_6_0; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_6_1; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_6_2; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_6_3; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_6_4; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_6_5; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_6_6; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_6_7; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_7_0; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_7_1; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_7_2; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_7_3; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_7_4; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_7_5; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_7_6; // @[PathFinder.scala 50:28]
  wire [31:0] Distribution_io_out_7_7; // @[PathFinder.scala 50:28]
  wire  Distribution_io_ProcessValid; // @[PathFinder.scala 50:28]
  wire  Distribution_io_valid; // @[PathFinder.scala 50:28]
  reg [31:0] delay; // @[PathFinder.scala 24:22]
  reg  high; // @[PathFinder.scala 26:21]
  reg  myCounter_io_start_REG; // @[PathFinder.scala 32:32]
  reg  high2; // @[PathFinder.scala 36:22]
  wire  _T_1 = delay < 32'h40 & high2; // @[PathFinder.scala 41:62]
  wire [31:0] _delay_T_1 = delay + 32'h1; // @[PathFinder.scala 42:20]
  wire  _GEN_2 = delay < 32'h40 & high2 & high2; // @[PathFinder.scala 36:22 41:72 47:11]
  wire  _GEN_3 = myCounter_io_valid | _GEN_2; // @[PathFinder.scala 39:28 40:11]
  wire [31:0] _GEN_79 = Distribution_io_ProcessValid ? Distribution_io_out_0_0 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_80 = Distribution_io_ProcessValid ? Distribution_io_out_0_1 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_81 = Distribution_io_ProcessValid ? Distribution_io_out_0_2 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_82 = Distribution_io_ProcessValid ? Distribution_io_out_0_3 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_83 = Distribution_io_ProcessValid ? Distribution_io_out_0_4 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_84 = Distribution_io_ProcessValid ? Distribution_io_out_0_5 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_85 = Distribution_io_ProcessValid ? Distribution_io_out_0_6 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_86 = Distribution_io_ProcessValid ? Distribution_io_out_0_7 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_87 = Distribution_io_ProcessValid ? Distribution_io_out_1_0 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_88 = Distribution_io_ProcessValid ? Distribution_io_out_1_1 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_89 = Distribution_io_ProcessValid ? Distribution_io_out_1_2 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_90 = Distribution_io_ProcessValid ? Distribution_io_out_1_3 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_91 = Distribution_io_ProcessValid ? Distribution_io_out_1_4 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_92 = Distribution_io_ProcessValid ? Distribution_io_out_1_5 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_93 = Distribution_io_ProcessValid ? Distribution_io_out_1_6 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_94 = Distribution_io_ProcessValid ? Distribution_io_out_1_7 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_95 = Distribution_io_ProcessValid ? Distribution_io_out_2_0 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_96 = Distribution_io_ProcessValid ? Distribution_io_out_2_1 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_97 = Distribution_io_ProcessValid ? Distribution_io_out_2_2 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_98 = Distribution_io_ProcessValid ? Distribution_io_out_2_3 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_99 = Distribution_io_ProcessValid ? Distribution_io_out_2_4 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_100 = Distribution_io_ProcessValid ? Distribution_io_out_2_5 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_101 = Distribution_io_ProcessValid ? Distribution_io_out_2_6 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_102 = Distribution_io_ProcessValid ? Distribution_io_out_2_7 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_103 = Distribution_io_ProcessValid ? Distribution_io_out_3_0 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_104 = Distribution_io_ProcessValid ? Distribution_io_out_3_1 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_105 = Distribution_io_ProcessValid ? Distribution_io_out_3_2 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_106 = Distribution_io_ProcessValid ? Distribution_io_out_3_3 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_107 = Distribution_io_ProcessValid ? Distribution_io_out_3_4 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_108 = Distribution_io_ProcessValid ? Distribution_io_out_3_5 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_109 = Distribution_io_ProcessValid ? Distribution_io_out_3_6 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_110 = Distribution_io_ProcessValid ? Distribution_io_out_3_7 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_111 = Distribution_io_ProcessValid ? Distribution_io_out_4_0 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_112 = Distribution_io_ProcessValid ? Distribution_io_out_4_1 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_113 = Distribution_io_ProcessValid ? Distribution_io_out_4_2 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_114 = Distribution_io_ProcessValid ? Distribution_io_out_4_3 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_115 = Distribution_io_ProcessValid ? Distribution_io_out_4_4 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_116 = Distribution_io_ProcessValid ? Distribution_io_out_4_5 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_117 = Distribution_io_ProcessValid ? Distribution_io_out_4_6 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_118 = Distribution_io_ProcessValid ? Distribution_io_out_4_7 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_119 = Distribution_io_ProcessValid ? Distribution_io_out_5_0 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_120 = Distribution_io_ProcessValid ? Distribution_io_out_5_1 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_121 = Distribution_io_ProcessValid ? Distribution_io_out_5_2 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_122 = Distribution_io_ProcessValid ? Distribution_io_out_5_3 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_123 = Distribution_io_ProcessValid ? Distribution_io_out_5_4 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_124 = Distribution_io_ProcessValid ? Distribution_io_out_5_5 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_125 = Distribution_io_ProcessValid ? Distribution_io_out_5_6 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_126 = Distribution_io_ProcessValid ? Distribution_io_out_5_7 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_127 = Distribution_io_ProcessValid ? Distribution_io_out_6_0 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_128 = Distribution_io_ProcessValid ? Distribution_io_out_6_1 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_129 = Distribution_io_ProcessValid ? Distribution_io_out_6_2 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_130 = Distribution_io_ProcessValid ? Distribution_io_out_6_3 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_131 = Distribution_io_ProcessValid ? Distribution_io_out_6_4 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_132 = Distribution_io_ProcessValid ? Distribution_io_out_6_5 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_133 = Distribution_io_ProcessValid ? Distribution_io_out_6_6 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_134 = Distribution_io_ProcessValid ? Distribution_io_out_6_7 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_135 = Distribution_io_ProcessValid ? Distribution_io_out_7_0 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_136 = Distribution_io_ProcessValid ? Distribution_io_out_7_1 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_137 = Distribution_io_ProcessValid ? Distribution_io_out_7_2 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_138 = Distribution_io_ProcessValid ? Distribution_io_out_7_3 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_139 = Distribution_io_ProcessValid ? Distribution_io_out_7_4 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_140 = Distribution_io_ProcessValid ? Distribution_io_out_7_5 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_141 = Distribution_io_ProcessValid ? Distribution_io_out_7_6 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_142 = Distribution_io_ProcessValid ? Distribution_io_out_7_7 : 32'h0; // @[PathFinder.scala 65:40 71:31 80:31]
  wire [31:0] _GEN_152 = io_DataValid ? {{28'd0}, myMuxes_io_i_mux_bus_0} : 32'h0; // @[PathFinder.scala 19:20 88:16 94:16]
  wire [31:0] _GEN_153 = io_DataValid ? {{28'd0}, myMuxes_io_i_mux_bus_1} : 32'h0; // @[PathFinder.scala 19:20 88:16 94:16]
  wire [31:0] _GEN_154 = io_DataValid ? {{28'd0}, myMuxes_io_i_mux_bus_2} : 32'h0; // @[PathFinder.scala 19:20 88:16 94:16]
  wire [31:0] _GEN_155 = io_DataValid ? {{28'd0}, myMuxes_io_i_mux_bus_3} : 32'h0; // @[PathFinder.scala 19:20 88:16 94:16]
  wire [31:0] _GEN_156 = io_DataValid ? {{16'd0}, myMuxes_io_Source_0} : 32'h0; // @[PathFinder.scala 19:20 89:13 95:13]
  wire [31:0] _GEN_157 = io_DataValid ? {{16'd0}, myMuxes_io_Source_1} : 32'h0; // @[PathFinder.scala 19:20 89:13 95:13]
  wire [31:0] _GEN_158 = io_DataValid ? {{16'd0}, myMuxes_io_Source_2} : 32'h0; // @[PathFinder.scala 19:20 89:13 95:13]
  wire [31:0] _GEN_159 = io_DataValid ? {{16'd0}, myMuxes_io_Source_3} : 32'h0; // @[PathFinder.scala 19:20 89:13 95:13]
  Muxes myMuxes ( // @[PathFinder.scala 25:23]
    .clock(myMuxes_clock),
    .reset(myMuxes_reset),
    .io_mat1_0_0(myMuxes_io_mat1_0_0),
    .io_mat1_0_1(myMuxes_io_mat1_0_1),
    .io_mat1_0_2(myMuxes_io_mat1_0_2),
    .io_mat1_0_3(myMuxes_io_mat1_0_3),
    .io_mat1_0_4(myMuxes_io_mat1_0_4),
    .io_mat1_0_5(myMuxes_io_mat1_0_5),
    .io_mat1_0_6(myMuxes_io_mat1_0_6),
    .io_mat1_0_7(myMuxes_io_mat1_0_7),
    .io_mat1_1_0(myMuxes_io_mat1_1_0),
    .io_mat1_1_1(myMuxes_io_mat1_1_1),
    .io_mat1_1_2(myMuxes_io_mat1_1_2),
    .io_mat1_1_3(myMuxes_io_mat1_1_3),
    .io_mat1_1_4(myMuxes_io_mat1_1_4),
    .io_mat1_1_5(myMuxes_io_mat1_1_5),
    .io_mat1_1_6(myMuxes_io_mat1_1_6),
    .io_mat1_1_7(myMuxes_io_mat1_1_7),
    .io_mat1_2_0(myMuxes_io_mat1_2_0),
    .io_mat1_2_1(myMuxes_io_mat1_2_1),
    .io_mat1_2_2(myMuxes_io_mat1_2_2),
    .io_mat1_2_3(myMuxes_io_mat1_2_3),
    .io_mat1_2_4(myMuxes_io_mat1_2_4),
    .io_mat1_2_5(myMuxes_io_mat1_2_5),
    .io_mat1_2_6(myMuxes_io_mat1_2_6),
    .io_mat1_2_7(myMuxes_io_mat1_2_7),
    .io_mat1_3_0(myMuxes_io_mat1_3_0),
    .io_mat1_3_1(myMuxes_io_mat1_3_1),
    .io_mat1_3_2(myMuxes_io_mat1_3_2),
    .io_mat1_3_3(myMuxes_io_mat1_3_3),
    .io_mat1_3_4(myMuxes_io_mat1_3_4),
    .io_mat1_3_5(myMuxes_io_mat1_3_5),
    .io_mat1_3_6(myMuxes_io_mat1_3_6),
    .io_mat1_3_7(myMuxes_io_mat1_3_7),
    .io_mat1_4_0(myMuxes_io_mat1_4_0),
    .io_mat1_4_1(myMuxes_io_mat1_4_1),
    .io_mat1_4_2(myMuxes_io_mat1_4_2),
    .io_mat1_4_3(myMuxes_io_mat1_4_3),
    .io_mat1_4_4(myMuxes_io_mat1_4_4),
    .io_mat1_4_5(myMuxes_io_mat1_4_5),
    .io_mat1_4_6(myMuxes_io_mat1_4_6),
    .io_mat1_4_7(myMuxes_io_mat1_4_7),
    .io_mat1_5_0(myMuxes_io_mat1_5_0),
    .io_mat1_5_1(myMuxes_io_mat1_5_1),
    .io_mat1_5_2(myMuxes_io_mat1_5_2),
    .io_mat1_5_3(myMuxes_io_mat1_5_3),
    .io_mat1_5_4(myMuxes_io_mat1_5_4),
    .io_mat1_5_5(myMuxes_io_mat1_5_5),
    .io_mat1_5_6(myMuxes_io_mat1_5_6),
    .io_mat1_5_7(myMuxes_io_mat1_5_7),
    .io_mat1_6_0(myMuxes_io_mat1_6_0),
    .io_mat1_6_1(myMuxes_io_mat1_6_1),
    .io_mat1_6_2(myMuxes_io_mat1_6_2),
    .io_mat1_6_3(myMuxes_io_mat1_6_3),
    .io_mat1_6_4(myMuxes_io_mat1_6_4),
    .io_mat1_6_5(myMuxes_io_mat1_6_5),
    .io_mat1_6_6(myMuxes_io_mat1_6_6),
    .io_mat1_6_7(myMuxes_io_mat1_6_7),
    .io_mat1_7_0(myMuxes_io_mat1_7_0),
    .io_mat1_7_1(myMuxes_io_mat1_7_1),
    .io_mat1_7_2(myMuxes_io_mat1_7_2),
    .io_mat1_7_3(myMuxes_io_mat1_7_3),
    .io_mat1_7_4(myMuxes_io_mat1_7_4),
    .io_mat1_7_5(myMuxes_io_mat1_7_5),
    .io_mat1_7_6(myMuxes_io_mat1_7_6),
    .io_mat1_7_7(myMuxes_io_mat1_7_7),
    .io_mat2_0(myMuxes_io_mat2_0),
    .io_mat2_1(myMuxes_io_mat2_1),
    .io_mat2_2(myMuxes_io_mat2_2),
    .io_mat2_3(myMuxes_io_mat2_3),
    .io_mat2_4(myMuxes_io_mat2_4),
    .io_mat2_5(myMuxes_io_mat2_5),
    .io_mat2_6(myMuxes_io_mat2_6),
    .io_mat2_7(myMuxes_io_mat2_7),
    .io_counterMatrix1_0_0(myMuxes_io_counterMatrix1_0_0),
    .io_counterMatrix1_0_1(myMuxes_io_counterMatrix1_0_1),
    .io_counterMatrix1_0_2(myMuxes_io_counterMatrix1_0_2),
    .io_counterMatrix1_0_3(myMuxes_io_counterMatrix1_0_3),
    .io_counterMatrix1_0_4(myMuxes_io_counterMatrix1_0_4),
    .io_counterMatrix1_0_5(myMuxes_io_counterMatrix1_0_5),
    .io_counterMatrix1_0_6(myMuxes_io_counterMatrix1_0_6),
    .io_counterMatrix1_0_7(myMuxes_io_counterMatrix1_0_7),
    .io_counterMatrix1_1_0(myMuxes_io_counterMatrix1_1_0),
    .io_counterMatrix1_1_1(myMuxes_io_counterMatrix1_1_1),
    .io_counterMatrix1_1_2(myMuxes_io_counterMatrix1_1_2),
    .io_counterMatrix1_1_3(myMuxes_io_counterMatrix1_1_3),
    .io_counterMatrix1_1_4(myMuxes_io_counterMatrix1_1_4),
    .io_counterMatrix1_1_5(myMuxes_io_counterMatrix1_1_5),
    .io_counterMatrix1_1_6(myMuxes_io_counterMatrix1_1_6),
    .io_counterMatrix1_1_7(myMuxes_io_counterMatrix1_1_7),
    .io_counterMatrix1_2_0(myMuxes_io_counterMatrix1_2_0),
    .io_counterMatrix1_2_1(myMuxes_io_counterMatrix1_2_1),
    .io_counterMatrix1_2_2(myMuxes_io_counterMatrix1_2_2),
    .io_counterMatrix1_2_3(myMuxes_io_counterMatrix1_2_3),
    .io_counterMatrix1_2_4(myMuxes_io_counterMatrix1_2_4),
    .io_counterMatrix1_2_5(myMuxes_io_counterMatrix1_2_5),
    .io_counterMatrix1_2_6(myMuxes_io_counterMatrix1_2_6),
    .io_counterMatrix1_2_7(myMuxes_io_counterMatrix1_2_7),
    .io_counterMatrix1_3_0(myMuxes_io_counterMatrix1_3_0),
    .io_counterMatrix1_3_1(myMuxes_io_counterMatrix1_3_1),
    .io_counterMatrix1_3_2(myMuxes_io_counterMatrix1_3_2),
    .io_counterMatrix1_3_3(myMuxes_io_counterMatrix1_3_3),
    .io_counterMatrix1_3_4(myMuxes_io_counterMatrix1_3_4),
    .io_counterMatrix1_3_5(myMuxes_io_counterMatrix1_3_5),
    .io_counterMatrix1_3_6(myMuxes_io_counterMatrix1_3_6),
    .io_counterMatrix1_3_7(myMuxes_io_counterMatrix1_3_7),
    .io_counterMatrix1_4_0(myMuxes_io_counterMatrix1_4_0),
    .io_counterMatrix1_4_1(myMuxes_io_counterMatrix1_4_1),
    .io_counterMatrix1_4_2(myMuxes_io_counterMatrix1_4_2),
    .io_counterMatrix1_4_3(myMuxes_io_counterMatrix1_4_3),
    .io_counterMatrix1_4_4(myMuxes_io_counterMatrix1_4_4),
    .io_counterMatrix1_4_5(myMuxes_io_counterMatrix1_4_5),
    .io_counterMatrix1_4_6(myMuxes_io_counterMatrix1_4_6),
    .io_counterMatrix1_4_7(myMuxes_io_counterMatrix1_4_7),
    .io_counterMatrix1_5_0(myMuxes_io_counterMatrix1_5_0),
    .io_counterMatrix1_5_1(myMuxes_io_counterMatrix1_5_1),
    .io_counterMatrix1_5_2(myMuxes_io_counterMatrix1_5_2),
    .io_counterMatrix1_5_3(myMuxes_io_counterMatrix1_5_3),
    .io_counterMatrix1_5_4(myMuxes_io_counterMatrix1_5_4),
    .io_counterMatrix1_5_5(myMuxes_io_counterMatrix1_5_5),
    .io_counterMatrix1_5_6(myMuxes_io_counterMatrix1_5_6),
    .io_counterMatrix1_5_7(myMuxes_io_counterMatrix1_5_7),
    .io_counterMatrix1_6_0(myMuxes_io_counterMatrix1_6_0),
    .io_counterMatrix1_6_1(myMuxes_io_counterMatrix1_6_1),
    .io_counterMatrix1_6_2(myMuxes_io_counterMatrix1_6_2),
    .io_counterMatrix1_6_3(myMuxes_io_counterMatrix1_6_3),
    .io_counterMatrix1_6_4(myMuxes_io_counterMatrix1_6_4),
    .io_counterMatrix1_6_5(myMuxes_io_counterMatrix1_6_5),
    .io_counterMatrix1_6_6(myMuxes_io_counterMatrix1_6_6),
    .io_counterMatrix1_6_7(myMuxes_io_counterMatrix1_6_7),
    .io_counterMatrix1_7_0(myMuxes_io_counterMatrix1_7_0),
    .io_counterMatrix1_7_1(myMuxes_io_counterMatrix1_7_1),
    .io_counterMatrix1_7_2(myMuxes_io_counterMatrix1_7_2),
    .io_counterMatrix1_7_3(myMuxes_io_counterMatrix1_7_3),
    .io_counterMatrix1_7_4(myMuxes_io_counterMatrix1_7_4),
    .io_counterMatrix1_7_5(myMuxes_io_counterMatrix1_7_5),
    .io_counterMatrix1_7_6(myMuxes_io_counterMatrix1_7_6),
    .io_counterMatrix1_7_7(myMuxes_io_counterMatrix1_7_7),
    .io_counterMatrix2_0(myMuxes_io_counterMatrix2_0),
    .io_counterMatrix2_1(myMuxes_io_counterMatrix2_1),
    .io_counterMatrix2_2(myMuxes_io_counterMatrix2_2),
    .io_counterMatrix2_3(myMuxes_io_counterMatrix2_3),
    .io_counterMatrix2_4(myMuxes_io_counterMatrix2_4),
    .io_counterMatrix2_5(myMuxes_io_counterMatrix2_5),
    .io_counterMatrix2_6(myMuxes_io_counterMatrix2_6),
    .io_counterMatrix2_7(myMuxes_io_counterMatrix2_7),
    .io_i_mux_bus_0(myMuxes_io_i_mux_bus_0),
    .io_i_mux_bus_1(myMuxes_io_i_mux_bus_1),
    .io_i_mux_bus_2(myMuxes_io_i_mux_bus_2),
    .io_i_mux_bus_3(myMuxes_io_i_mux_bus_3),
    .io_Source_0(myMuxes_io_Source_0),
    .io_Source_1(myMuxes_io_Source_1),
    .io_Source_2(myMuxes_io_Source_2),
    .io_Source_3(myMuxes_io_Source_3),
    .io_valid(myMuxes_io_valid)
  );
  SourceDestination myCounter ( // @[PathFinder.scala 31:25]
    .clock(myCounter_clock),
    .reset(myCounter_reset),
    .io_Stationary_matrix_0_0(myCounter_io_Stationary_matrix_0_0),
    .io_Stationary_matrix_0_1(myCounter_io_Stationary_matrix_0_1),
    .io_Stationary_matrix_0_2(myCounter_io_Stationary_matrix_0_2),
    .io_Stationary_matrix_0_3(myCounter_io_Stationary_matrix_0_3),
    .io_Stationary_matrix_0_4(myCounter_io_Stationary_matrix_0_4),
    .io_Stationary_matrix_0_5(myCounter_io_Stationary_matrix_0_5),
    .io_Stationary_matrix_0_6(myCounter_io_Stationary_matrix_0_6),
    .io_Stationary_matrix_0_7(myCounter_io_Stationary_matrix_0_7),
    .io_Stationary_matrix_1_0(myCounter_io_Stationary_matrix_1_0),
    .io_Stationary_matrix_1_1(myCounter_io_Stationary_matrix_1_1),
    .io_Stationary_matrix_1_2(myCounter_io_Stationary_matrix_1_2),
    .io_Stationary_matrix_1_3(myCounter_io_Stationary_matrix_1_3),
    .io_Stationary_matrix_1_4(myCounter_io_Stationary_matrix_1_4),
    .io_Stationary_matrix_1_5(myCounter_io_Stationary_matrix_1_5),
    .io_Stationary_matrix_1_6(myCounter_io_Stationary_matrix_1_6),
    .io_Stationary_matrix_1_7(myCounter_io_Stationary_matrix_1_7),
    .io_Stationary_matrix_2_0(myCounter_io_Stationary_matrix_2_0),
    .io_Stationary_matrix_2_1(myCounter_io_Stationary_matrix_2_1),
    .io_Stationary_matrix_2_2(myCounter_io_Stationary_matrix_2_2),
    .io_Stationary_matrix_2_3(myCounter_io_Stationary_matrix_2_3),
    .io_Stationary_matrix_2_4(myCounter_io_Stationary_matrix_2_4),
    .io_Stationary_matrix_2_5(myCounter_io_Stationary_matrix_2_5),
    .io_Stationary_matrix_2_6(myCounter_io_Stationary_matrix_2_6),
    .io_Stationary_matrix_2_7(myCounter_io_Stationary_matrix_2_7),
    .io_Stationary_matrix_3_0(myCounter_io_Stationary_matrix_3_0),
    .io_Stationary_matrix_3_1(myCounter_io_Stationary_matrix_3_1),
    .io_Stationary_matrix_3_2(myCounter_io_Stationary_matrix_3_2),
    .io_Stationary_matrix_3_3(myCounter_io_Stationary_matrix_3_3),
    .io_Stationary_matrix_3_4(myCounter_io_Stationary_matrix_3_4),
    .io_Stationary_matrix_3_5(myCounter_io_Stationary_matrix_3_5),
    .io_Stationary_matrix_3_6(myCounter_io_Stationary_matrix_3_6),
    .io_Stationary_matrix_3_7(myCounter_io_Stationary_matrix_3_7),
    .io_Stationary_matrix_4_0(myCounter_io_Stationary_matrix_4_0),
    .io_Stationary_matrix_4_1(myCounter_io_Stationary_matrix_4_1),
    .io_Stationary_matrix_4_2(myCounter_io_Stationary_matrix_4_2),
    .io_Stationary_matrix_4_3(myCounter_io_Stationary_matrix_4_3),
    .io_Stationary_matrix_4_4(myCounter_io_Stationary_matrix_4_4),
    .io_Stationary_matrix_4_5(myCounter_io_Stationary_matrix_4_5),
    .io_Stationary_matrix_4_6(myCounter_io_Stationary_matrix_4_6),
    .io_Stationary_matrix_4_7(myCounter_io_Stationary_matrix_4_7),
    .io_Stationary_matrix_5_0(myCounter_io_Stationary_matrix_5_0),
    .io_Stationary_matrix_5_1(myCounter_io_Stationary_matrix_5_1),
    .io_Stationary_matrix_5_2(myCounter_io_Stationary_matrix_5_2),
    .io_Stationary_matrix_5_3(myCounter_io_Stationary_matrix_5_3),
    .io_Stationary_matrix_5_4(myCounter_io_Stationary_matrix_5_4),
    .io_Stationary_matrix_5_5(myCounter_io_Stationary_matrix_5_5),
    .io_Stationary_matrix_5_6(myCounter_io_Stationary_matrix_5_6),
    .io_Stationary_matrix_5_7(myCounter_io_Stationary_matrix_5_7),
    .io_Stationary_matrix_6_0(myCounter_io_Stationary_matrix_6_0),
    .io_Stationary_matrix_6_1(myCounter_io_Stationary_matrix_6_1),
    .io_Stationary_matrix_6_2(myCounter_io_Stationary_matrix_6_2),
    .io_Stationary_matrix_6_3(myCounter_io_Stationary_matrix_6_3),
    .io_Stationary_matrix_6_4(myCounter_io_Stationary_matrix_6_4),
    .io_Stationary_matrix_6_5(myCounter_io_Stationary_matrix_6_5),
    .io_Stationary_matrix_6_6(myCounter_io_Stationary_matrix_6_6),
    .io_Stationary_matrix_6_7(myCounter_io_Stationary_matrix_6_7),
    .io_Stationary_matrix_7_0(myCounter_io_Stationary_matrix_7_0),
    .io_Stationary_matrix_7_1(myCounter_io_Stationary_matrix_7_1),
    .io_Stationary_matrix_7_2(myCounter_io_Stationary_matrix_7_2),
    .io_Stationary_matrix_7_3(myCounter_io_Stationary_matrix_7_3),
    .io_Stationary_matrix_7_4(myCounter_io_Stationary_matrix_7_4),
    .io_Stationary_matrix_7_5(myCounter_io_Stationary_matrix_7_5),
    .io_Stationary_matrix_7_6(myCounter_io_Stationary_matrix_7_6),
    .io_Stationary_matrix_7_7(myCounter_io_Stationary_matrix_7_7),
    .io_Streaming_matrix_0(myCounter_io_Streaming_matrix_0),
    .io_Streaming_matrix_1(myCounter_io_Streaming_matrix_1),
    .io_Streaming_matrix_2(myCounter_io_Streaming_matrix_2),
    .io_Streaming_matrix_3(myCounter_io_Streaming_matrix_3),
    .io_Streaming_matrix_4(myCounter_io_Streaming_matrix_4),
    .io_Streaming_matrix_5(myCounter_io_Streaming_matrix_5),
    .io_Streaming_matrix_6(myCounter_io_Streaming_matrix_6),
    .io_Streaming_matrix_7(myCounter_io_Streaming_matrix_7),
    .io_counterMatrix1_bits_0_0(myCounter_io_counterMatrix1_bits_0_0),
    .io_counterMatrix1_bits_0_1(myCounter_io_counterMatrix1_bits_0_1),
    .io_counterMatrix1_bits_0_2(myCounter_io_counterMatrix1_bits_0_2),
    .io_counterMatrix1_bits_0_3(myCounter_io_counterMatrix1_bits_0_3),
    .io_counterMatrix1_bits_0_4(myCounter_io_counterMatrix1_bits_0_4),
    .io_counterMatrix1_bits_0_5(myCounter_io_counterMatrix1_bits_0_5),
    .io_counterMatrix1_bits_0_6(myCounter_io_counterMatrix1_bits_0_6),
    .io_counterMatrix1_bits_0_7(myCounter_io_counterMatrix1_bits_0_7),
    .io_counterMatrix1_bits_1_0(myCounter_io_counterMatrix1_bits_1_0),
    .io_counterMatrix1_bits_1_1(myCounter_io_counterMatrix1_bits_1_1),
    .io_counterMatrix1_bits_1_2(myCounter_io_counterMatrix1_bits_1_2),
    .io_counterMatrix1_bits_1_3(myCounter_io_counterMatrix1_bits_1_3),
    .io_counterMatrix1_bits_1_4(myCounter_io_counterMatrix1_bits_1_4),
    .io_counterMatrix1_bits_1_5(myCounter_io_counterMatrix1_bits_1_5),
    .io_counterMatrix1_bits_1_6(myCounter_io_counterMatrix1_bits_1_6),
    .io_counterMatrix1_bits_1_7(myCounter_io_counterMatrix1_bits_1_7),
    .io_counterMatrix1_bits_2_0(myCounter_io_counterMatrix1_bits_2_0),
    .io_counterMatrix1_bits_2_1(myCounter_io_counterMatrix1_bits_2_1),
    .io_counterMatrix1_bits_2_2(myCounter_io_counterMatrix1_bits_2_2),
    .io_counterMatrix1_bits_2_3(myCounter_io_counterMatrix1_bits_2_3),
    .io_counterMatrix1_bits_2_4(myCounter_io_counterMatrix1_bits_2_4),
    .io_counterMatrix1_bits_2_5(myCounter_io_counterMatrix1_bits_2_5),
    .io_counterMatrix1_bits_2_6(myCounter_io_counterMatrix1_bits_2_6),
    .io_counterMatrix1_bits_2_7(myCounter_io_counterMatrix1_bits_2_7),
    .io_counterMatrix1_bits_3_0(myCounter_io_counterMatrix1_bits_3_0),
    .io_counterMatrix1_bits_3_1(myCounter_io_counterMatrix1_bits_3_1),
    .io_counterMatrix1_bits_3_2(myCounter_io_counterMatrix1_bits_3_2),
    .io_counterMatrix1_bits_3_3(myCounter_io_counterMatrix1_bits_3_3),
    .io_counterMatrix1_bits_3_4(myCounter_io_counterMatrix1_bits_3_4),
    .io_counterMatrix1_bits_3_5(myCounter_io_counterMatrix1_bits_3_5),
    .io_counterMatrix1_bits_3_6(myCounter_io_counterMatrix1_bits_3_6),
    .io_counterMatrix1_bits_3_7(myCounter_io_counterMatrix1_bits_3_7),
    .io_counterMatrix1_bits_4_0(myCounter_io_counterMatrix1_bits_4_0),
    .io_counterMatrix1_bits_4_1(myCounter_io_counterMatrix1_bits_4_1),
    .io_counterMatrix1_bits_4_2(myCounter_io_counterMatrix1_bits_4_2),
    .io_counterMatrix1_bits_4_3(myCounter_io_counterMatrix1_bits_4_3),
    .io_counterMatrix1_bits_4_4(myCounter_io_counterMatrix1_bits_4_4),
    .io_counterMatrix1_bits_4_5(myCounter_io_counterMatrix1_bits_4_5),
    .io_counterMatrix1_bits_4_6(myCounter_io_counterMatrix1_bits_4_6),
    .io_counterMatrix1_bits_4_7(myCounter_io_counterMatrix1_bits_4_7),
    .io_counterMatrix1_bits_5_0(myCounter_io_counterMatrix1_bits_5_0),
    .io_counterMatrix1_bits_5_1(myCounter_io_counterMatrix1_bits_5_1),
    .io_counterMatrix1_bits_5_2(myCounter_io_counterMatrix1_bits_5_2),
    .io_counterMatrix1_bits_5_3(myCounter_io_counterMatrix1_bits_5_3),
    .io_counterMatrix1_bits_5_4(myCounter_io_counterMatrix1_bits_5_4),
    .io_counterMatrix1_bits_5_5(myCounter_io_counterMatrix1_bits_5_5),
    .io_counterMatrix1_bits_5_6(myCounter_io_counterMatrix1_bits_5_6),
    .io_counterMatrix1_bits_5_7(myCounter_io_counterMatrix1_bits_5_7),
    .io_counterMatrix1_bits_6_0(myCounter_io_counterMatrix1_bits_6_0),
    .io_counterMatrix1_bits_6_1(myCounter_io_counterMatrix1_bits_6_1),
    .io_counterMatrix1_bits_6_2(myCounter_io_counterMatrix1_bits_6_2),
    .io_counterMatrix1_bits_6_3(myCounter_io_counterMatrix1_bits_6_3),
    .io_counterMatrix1_bits_6_4(myCounter_io_counterMatrix1_bits_6_4),
    .io_counterMatrix1_bits_6_5(myCounter_io_counterMatrix1_bits_6_5),
    .io_counterMatrix1_bits_6_6(myCounter_io_counterMatrix1_bits_6_6),
    .io_counterMatrix1_bits_6_7(myCounter_io_counterMatrix1_bits_6_7),
    .io_counterMatrix1_bits_7_0(myCounter_io_counterMatrix1_bits_7_0),
    .io_counterMatrix1_bits_7_1(myCounter_io_counterMatrix1_bits_7_1),
    .io_counterMatrix1_bits_7_2(myCounter_io_counterMatrix1_bits_7_2),
    .io_counterMatrix1_bits_7_3(myCounter_io_counterMatrix1_bits_7_3),
    .io_counterMatrix1_bits_7_4(myCounter_io_counterMatrix1_bits_7_4),
    .io_counterMatrix1_bits_7_5(myCounter_io_counterMatrix1_bits_7_5),
    .io_counterMatrix1_bits_7_6(myCounter_io_counterMatrix1_bits_7_6),
    .io_counterMatrix1_bits_7_7(myCounter_io_counterMatrix1_bits_7_7),
    .io_counterMatrix2_bits_0(myCounter_io_counterMatrix2_bits_0),
    .io_counterMatrix2_bits_1(myCounter_io_counterMatrix2_bits_1),
    .io_counterMatrix2_bits_2(myCounter_io_counterMatrix2_bits_2),
    .io_counterMatrix2_bits_3(myCounter_io_counterMatrix2_bits_3),
    .io_counterMatrix2_bits_4(myCounter_io_counterMatrix2_bits_4),
    .io_counterMatrix2_bits_5(myCounter_io_counterMatrix2_bits_5),
    .io_counterMatrix2_bits_6(myCounter_io_counterMatrix2_bits_6),
    .io_counterMatrix2_bits_7(myCounter_io_counterMatrix2_bits_7),
    .io_valid(myCounter_io_valid),
    .io_start(myCounter_io_start)
  );
  Distribution2 Distribution ( // @[PathFinder.scala 50:28]
    .clock(Distribution_clock),
    .reset(Distribution_reset),
    .io_matrix_0_0(Distribution_io_matrix_0_0),
    .io_matrix_0_1(Distribution_io_matrix_0_1),
    .io_matrix_0_2(Distribution_io_matrix_0_2),
    .io_matrix_0_3(Distribution_io_matrix_0_3),
    .io_matrix_0_4(Distribution_io_matrix_0_4),
    .io_matrix_0_5(Distribution_io_matrix_0_5),
    .io_matrix_0_6(Distribution_io_matrix_0_6),
    .io_matrix_0_7(Distribution_io_matrix_0_7),
    .io_matrix_1_0(Distribution_io_matrix_1_0),
    .io_matrix_1_1(Distribution_io_matrix_1_1),
    .io_matrix_1_2(Distribution_io_matrix_1_2),
    .io_matrix_1_3(Distribution_io_matrix_1_3),
    .io_matrix_1_4(Distribution_io_matrix_1_4),
    .io_matrix_1_5(Distribution_io_matrix_1_5),
    .io_matrix_1_6(Distribution_io_matrix_1_6),
    .io_matrix_1_7(Distribution_io_matrix_1_7),
    .io_matrix_2_0(Distribution_io_matrix_2_0),
    .io_matrix_2_1(Distribution_io_matrix_2_1),
    .io_matrix_2_2(Distribution_io_matrix_2_2),
    .io_matrix_2_3(Distribution_io_matrix_2_3),
    .io_matrix_2_4(Distribution_io_matrix_2_4),
    .io_matrix_2_5(Distribution_io_matrix_2_5),
    .io_matrix_2_6(Distribution_io_matrix_2_6),
    .io_matrix_2_7(Distribution_io_matrix_2_7),
    .io_matrix_3_0(Distribution_io_matrix_3_0),
    .io_matrix_3_1(Distribution_io_matrix_3_1),
    .io_matrix_3_2(Distribution_io_matrix_3_2),
    .io_matrix_3_3(Distribution_io_matrix_3_3),
    .io_matrix_3_4(Distribution_io_matrix_3_4),
    .io_matrix_3_5(Distribution_io_matrix_3_5),
    .io_matrix_3_6(Distribution_io_matrix_3_6),
    .io_matrix_3_7(Distribution_io_matrix_3_7),
    .io_matrix_4_0(Distribution_io_matrix_4_0),
    .io_matrix_4_1(Distribution_io_matrix_4_1),
    .io_matrix_4_2(Distribution_io_matrix_4_2),
    .io_matrix_4_3(Distribution_io_matrix_4_3),
    .io_matrix_4_4(Distribution_io_matrix_4_4),
    .io_matrix_4_5(Distribution_io_matrix_4_5),
    .io_matrix_4_6(Distribution_io_matrix_4_6),
    .io_matrix_4_7(Distribution_io_matrix_4_7),
    .io_matrix_5_0(Distribution_io_matrix_5_0),
    .io_matrix_5_1(Distribution_io_matrix_5_1),
    .io_matrix_5_2(Distribution_io_matrix_5_2),
    .io_matrix_5_3(Distribution_io_matrix_5_3),
    .io_matrix_5_4(Distribution_io_matrix_5_4),
    .io_matrix_5_5(Distribution_io_matrix_5_5),
    .io_matrix_5_6(Distribution_io_matrix_5_6),
    .io_matrix_5_7(Distribution_io_matrix_5_7),
    .io_matrix_6_0(Distribution_io_matrix_6_0),
    .io_matrix_6_1(Distribution_io_matrix_6_1),
    .io_matrix_6_2(Distribution_io_matrix_6_2),
    .io_matrix_6_3(Distribution_io_matrix_6_3),
    .io_matrix_6_4(Distribution_io_matrix_6_4),
    .io_matrix_6_5(Distribution_io_matrix_6_5),
    .io_matrix_6_6(Distribution_io_matrix_6_6),
    .io_matrix_6_7(Distribution_io_matrix_6_7),
    .io_matrix_7_0(Distribution_io_matrix_7_0),
    .io_matrix_7_1(Distribution_io_matrix_7_1),
    .io_matrix_7_2(Distribution_io_matrix_7_2),
    .io_matrix_7_3(Distribution_io_matrix_7_3),
    .io_matrix_7_4(Distribution_io_matrix_7_4),
    .io_matrix_7_5(Distribution_io_matrix_7_5),
    .io_matrix_7_6(Distribution_io_matrix_7_6),
    .io_matrix_7_7(Distribution_io_matrix_7_7),
    .io_s(Distribution_io_s),
    .io_out_0_0(Distribution_io_out_0_0),
    .io_out_0_1(Distribution_io_out_0_1),
    .io_out_0_2(Distribution_io_out_0_2),
    .io_out_0_3(Distribution_io_out_0_3),
    .io_out_0_4(Distribution_io_out_0_4),
    .io_out_0_5(Distribution_io_out_0_5),
    .io_out_0_6(Distribution_io_out_0_6),
    .io_out_0_7(Distribution_io_out_0_7),
    .io_out_1_0(Distribution_io_out_1_0),
    .io_out_1_1(Distribution_io_out_1_1),
    .io_out_1_2(Distribution_io_out_1_2),
    .io_out_1_3(Distribution_io_out_1_3),
    .io_out_1_4(Distribution_io_out_1_4),
    .io_out_1_5(Distribution_io_out_1_5),
    .io_out_1_6(Distribution_io_out_1_6),
    .io_out_1_7(Distribution_io_out_1_7),
    .io_out_2_0(Distribution_io_out_2_0),
    .io_out_2_1(Distribution_io_out_2_1),
    .io_out_2_2(Distribution_io_out_2_2),
    .io_out_2_3(Distribution_io_out_2_3),
    .io_out_2_4(Distribution_io_out_2_4),
    .io_out_2_5(Distribution_io_out_2_5),
    .io_out_2_6(Distribution_io_out_2_6),
    .io_out_2_7(Distribution_io_out_2_7),
    .io_out_3_0(Distribution_io_out_3_0),
    .io_out_3_1(Distribution_io_out_3_1),
    .io_out_3_2(Distribution_io_out_3_2),
    .io_out_3_3(Distribution_io_out_3_3),
    .io_out_3_4(Distribution_io_out_3_4),
    .io_out_3_5(Distribution_io_out_3_5),
    .io_out_3_6(Distribution_io_out_3_6),
    .io_out_3_7(Distribution_io_out_3_7),
    .io_out_4_0(Distribution_io_out_4_0),
    .io_out_4_1(Distribution_io_out_4_1),
    .io_out_4_2(Distribution_io_out_4_2),
    .io_out_4_3(Distribution_io_out_4_3),
    .io_out_4_4(Distribution_io_out_4_4),
    .io_out_4_5(Distribution_io_out_4_5),
    .io_out_4_6(Distribution_io_out_4_6),
    .io_out_4_7(Distribution_io_out_4_7),
    .io_out_5_0(Distribution_io_out_5_0),
    .io_out_5_1(Distribution_io_out_5_1),
    .io_out_5_2(Distribution_io_out_5_2),
    .io_out_5_3(Distribution_io_out_5_3),
    .io_out_5_4(Distribution_io_out_5_4),
    .io_out_5_5(Distribution_io_out_5_5),
    .io_out_5_6(Distribution_io_out_5_6),
    .io_out_5_7(Distribution_io_out_5_7),
    .io_out_6_0(Distribution_io_out_6_0),
    .io_out_6_1(Distribution_io_out_6_1),
    .io_out_6_2(Distribution_io_out_6_2),
    .io_out_6_3(Distribution_io_out_6_3),
    .io_out_6_4(Distribution_io_out_6_4),
    .io_out_6_5(Distribution_io_out_6_5),
    .io_out_6_6(Distribution_io_out_6_6),
    .io_out_6_7(Distribution_io_out_6_7),
    .io_out_7_0(Distribution_io_out_7_0),
    .io_out_7_1(Distribution_io_out_7_1),
    .io_out_7_2(Distribution_io_out_7_2),
    .io_out_7_3(Distribution_io_out_7_3),
    .io_out_7_4(Distribution_io_out_7_4),
    .io_out_7_5(Distribution_io_out_7_5),
    .io_out_7_6(Distribution_io_out_7_6),
    .io_out_7_7(Distribution_io_out_7_7),
    .io_ProcessValid(Distribution_io_ProcessValid),
    .io_valid(Distribution_io_valid)
  );
  assign io_i_mux_bus_0 = _GEN_152[3:0];
  assign io_i_mux_bus_1 = _GEN_153[3:0];
  assign io_i_mux_bus_2 = _GEN_154[3:0];
  assign io_i_mux_bus_3 = _GEN_155[3:0];
  assign io_Source_0 = _GEN_156[15:0];
  assign io_Source_1 = _GEN_157[15:0];
  assign io_Source_2 = _GEN_158[15:0];
  assign io_Source_3 = _GEN_159[15:0];
  assign io_PF_Valid = io_DataValid & myMuxes_io_valid; // @[PathFinder.scala 19:20 87:15 93:15]
  assign myMuxes_clock = clock;
  assign myMuxes_reset = reset;
  assign myMuxes_io_mat1_0_0 = Distribution_io_ProcessValid ? io_Stationary_matrix_0_0 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_0_1 = Distribution_io_ProcessValid ? io_Stationary_matrix_0_1 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_0_2 = Distribution_io_ProcessValid ? io_Stationary_matrix_0_2 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_0_3 = Distribution_io_ProcessValid ? io_Stationary_matrix_0_3 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_0_4 = Distribution_io_ProcessValid ? io_Stationary_matrix_0_4 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_0_5 = Distribution_io_ProcessValid ? io_Stationary_matrix_0_5 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_0_6 = Distribution_io_ProcessValid ? io_Stationary_matrix_0_6 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_0_7 = Distribution_io_ProcessValid ? io_Stationary_matrix_0_7 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_1_0 = Distribution_io_ProcessValid ? io_Stationary_matrix_1_0 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_1_1 = Distribution_io_ProcessValid ? io_Stationary_matrix_1_1 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_1_2 = Distribution_io_ProcessValid ? io_Stationary_matrix_1_2 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_1_3 = Distribution_io_ProcessValid ? io_Stationary_matrix_1_3 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_1_4 = Distribution_io_ProcessValid ? io_Stationary_matrix_1_4 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_1_5 = Distribution_io_ProcessValid ? io_Stationary_matrix_1_5 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_1_6 = Distribution_io_ProcessValid ? io_Stationary_matrix_1_6 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_1_7 = Distribution_io_ProcessValid ? io_Stationary_matrix_1_7 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_2_0 = Distribution_io_ProcessValid ? io_Stationary_matrix_2_0 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_2_1 = Distribution_io_ProcessValid ? io_Stationary_matrix_2_1 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_2_2 = Distribution_io_ProcessValid ? io_Stationary_matrix_2_2 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_2_3 = Distribution_io_ProcessValid ? io_Stationary_matrix_2_3 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_2_4 = Distribution_io_ProcessValid ? io_Stationary_matrix_2_4 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_2_5 = Distribution_io_ProcessValid ? io_Stationary_matrix_2_5 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_2_6 = Distribution_io_ProcessValid ? io_Stationary_matrix_2_6 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_2_7 = Distribution_io_ProcessValid ? io_Stationary_matrix_2_7 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_3_0 = Distribution_io_ProcessValid ? io_Stationary_matrix_3_0 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_3_1 = Distribution_io_ProcessValid ? io_Stationary_matrix_3_1 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_3_2 = Distribution_io_ProcessValid ? io_Stationary_matrix_3_2 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_3_3 = Distribution_io_ProcessValid ? io_Stationary_matrix_3_3 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_3_4 = Distribution_io_ProcessValid ? io_Stationary_matrix_3_4 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_3_5 = Distribution_io_ProcessValid ? io_Stationary_matrix_3_5 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_3_6 = Distribution_io_ProcessValid ? io_Stationary_matrix_3_6 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_3_7 = Distribution_io_ProcessValid ? io_Stationary_matrix_3_7 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_4_0 = Distribution_io_ProcessValid ? io_Stationary_matrix_4_0 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_4_1 = Distribution_io_ProcessValid ? io_Stationary_matrix_4_1 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_4_2 = Distribution_io_ProcessValid ? io_Stationary_matrix_4_2 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_4_3 = Distribution_io_ProcessValid ? io_Stationary_matrix_4_3 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_4_4 = Distribution_io_ProcessValid ? io_Stationary_matrix_4_4 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_4_5 = Distribution_io_ProcessValid ? io_Stationary_matrix_4_5 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_4_6 = Distribution_io_ProcessValid ? io_Stationary_matrix_4_6 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_4_7 = Distribution_io_ProcessValid ? io_Stationary_matrix_4_7 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_5_0 = Distribution_io_ProcessValid ? io_Stationary_matrix_5_0 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_5_1 = Distribution_io_ProcessValid ? io_Stationary_matrix_5_1 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_5_2 = Distribution_io_ProcessValid ? io_Stationary_matrix_5_2 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_5_3 = Distribution_io_ProcessValid ? io_Stationary_matrix_5_3 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_5_4 = Distribution_io_ProcessValid ? io_Stationary_matrix_5_4 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_5_5 = Distribution_io_ProcessValid ? io_Stationary_matrix_5_5 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_5_6 = Distribution_io_ProcessValid ? io_Stationary_matrix_5_6 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_5_7 = Distribution_io_ProcessValid ? io_Stationary_matrix_5_7 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_6_0 = Distribution_io_ProcessValid ? io_Stationary_matrix_6_0 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_6_1 = Distribution_io_ProcessValid ? io_Stationary_matrix_6_1 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_6_2 = Distribution_io_ProcessValid ? io_Stationary_matrix_6_2 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_6_3 = Distribution_io_ProcessValid ? io_Stationary_matrix_6_3 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_6_4 = Distribution_io_ProcessValid ? io_Stationary_matrix_6_4 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_6_5 = Distribution_io_ProcessValid ? io_Stationary_matrix_6_5 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_6_6 = Distribution_io_ProcessValid ? io_Stationary_matrix_6_6 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_6_7 = Distribution_io_ProcessValid ? io_Stationary_matrix_6_7 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_7_0 = Distribution_io_ProcessValid ? io_Stationary_matrix_7_0 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_7_1 = Distribution_io_ProcessValid ? io_Stationary_matrix_7_1 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_7_2 = Distribution_io_ProcessValid ? io_Stationary_matrix_7_2 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_7_3 = Distribution_io_ProcessValid ? io_Stationary_matrix_7_3 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_7_4 = Distribution_io_ProcessValid ? io_Stationary_matrix_7_4 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_7_5 = Distribution_io_ProcessValid ? io_Stationary_matrix_7_5 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_7_6 = Distribution_io_ProcessValid ? io_Stationary_matrix_7_6 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat1_7_7 = Distribution_io_ProcessValid ? io_Stationary_matrix_7_7 : 16'h0; // @[PathFinder.scala 65:40 68:21 78:21]
  assign myMuxes_io_mat2_0 = Distribution_io_ProcessValid ? io_Streaming_matrix_0 : 16'h0; // @[PathFinder.scala 65:40 70:21 79:21]
  assign myMuxes_io_mat2_1 = Distribution_io_ProcessValid ? io_Streaming_matrix_1 : 16'h0; // @[PathFinder.scala 65:40 70:21 79:21]
  assign myMuxes_io_mat2_2 = Distribution_io_ProcessValid ? io_Streaming_matrix_2 : 16'h0; // @[PathFinder.scala 65:40 70:21 79:21]
  assign myMuxes_io_mat2_3 = Distribution_io_ProcessValid ? io_Streaming_matrix_3 : 16'h0; // @[PathFinder.scala 65:40 70:21 79:21]
  assign myMuxes_io_mat2_4 = Distribution_io_ProcessValid ? io_Streaming_matrix_4 : 16'h0; // @[PathFinder.scala 65:40 70:21 79:21]
  assign myMuxes_io_mat2_5 = Distribution_io_ProcessValid ? io_Streaming_matrix_5 : 16'h0; // @[PathFinder.scala 65:40 70:21 79:21]
  assign myMuxes_io_mat2_6 = Distribution_io_ProcessValid ? io_Streaming_matrix_6 : 16'h0; // @[PathFinder.scala 65:40 70:21 79:21]
  assign myMuxes_io_mat2_7 = Distribution_io_ProcessValid ? io_Streaming_matrix_7 : 16'h0; // @[PathFinder.scala 65:40 70:21 79:21]
  assign myMuxes_io_counterMatrix1_0_0 = _GEN_79[15:0];
  assign myMuxes_io_counterMatrix1_0_1 = _GEN_80[15:0];
  assign myMuxes_io_counterMatrix1_0_2 = _GEN_81[15:0];
  assign myMuxes_io_counterMatrix1_0_3 = _GEN_82[15:0];
  assign myMuxes_io_counterMatrix1_0_4 = _GEN_83[15:0];
  assign myMuxes_io_counterMatrix1_0_5 = _GEN_84[15:0];
  assign myMuxes_io_counterMatrix1_0_6 = _GEN_85[15:0];
  assign myMuxes_io_counterMatrix1_0_7 = _GEN_86[15:0];
  assign myMuxes_io_counterMatrix1_1_0 = _GEN_87[15:0];
  assign myMuxes_io_counterMatrix1_1_1 = _GEN_88[15:0];
  assign myMuxes_io_counterMatrix1_1_2 = _GEN_89[15:0];
  assign myMuxes_io_counterMatrix1_1_3 = _GEN_90[15:0];
  assign myMuxes_io_counterMatrix1_1_4 = _GEN_91[15:0];
  assign myMuxes_io_counterMatrix1_1_5 = _GEN_92[15:0];
  assign myMuxes_io_counterMatrix1_1_6 = _GEN_93[15:0];
  assign myMuxes_io_counterMatrix1_1_7 = _GEN_94[15:0];
  assign myMuxes_io_counterMatrix1_2_0 = _GEN_95[15:0];
  assign myMuxes_io_counterMatrix1_2_1 = _GEN_96[15:0];
  assign myMuxes_io_counterMatrix1_2_2 = _GEN_97[15:0];
  assign myMuxes_io_counterMatrix1_2_3 = _GEN_98[15:0];
  assign myMuxes_io_counterMatrix1_2_4 = _GEN_99[15:0];
  assign myMuxes_io_counterMatrix1_2_5 = _GEN_100[15:0];
  assign myMuxes_io_counterMatrix1_2_6 = _GEN_101[15:0];
  assign myMuxes_io_counterMatrix1_2_7 = _GEN_102[15:0];
  assign myMuxes_io_counterMatrix1_3_0 = _GEN_103[15:0];
  assign myMuxes_io_counterMatrix1_3_1 = _GEN_104[15:0];
  assign myMuxes_io_counterMatrix1_3_2 = _GEN_105[15:0];
  assign myMuxes_io_counterMatrix1_3_3 = _GEN_106[15:0];
  assign myMuxes_io_counterMatrix1_3_4 = _GEN_107[15:0];
  assign myMuxes_io_counterMatrix1_3_5 = _GEN_108[15:0];
  assign myMuxes_io_counterMatrix1_3_6 = _GEN_109[15:0];
  assign myMuxes_io_counterMatrix1_3_7 = _GEN_110[15:0];
  assign myMuxes_io_counterMatrix1_4_0 = _GEN_111[15:0];
  assign myMuxes_io_counterMatrix1_4_1 = _GEN_112[15:0];
  assign myMuxes_io_counterMatrix1_4_2 = _GEN_113[15:0];
  assign myMuxes_io_counterMatrix1_4_3 = _GEN_114[15:0];
  assign myMuxes_io_counterMatrix1_4_4 = _GEN_115[15:0];
  assign myMuxes_io_counterMatrix1_4_5 = _GEN_116[15:0];
  assign myMuxes_io_counterMatrix1_4_6 = _GEN_117[15:0];
  assign myMuxes_io_counterMatrix1_4_7 = _GEN_118[15:0];
  assign myMuxes_io_counterMatrix1_5_0 = _GEN_119[15:0];
  assign myMuxes_io_counterMatrix1_5_1 = _GEN_120[15:0];
  assign myMuxes_io_counterMatrix1_5_2 = _GEN_121[15:0];
  assign myMuxes_io_counterMatrix1_5_3 = _GEN_122[15:0];
  assign myMuxes_io_counterMatrix1_5_4 = _GEN_123[15:0];
  assign myMuxes_io_counterMatrix1_5_5 = _GEN_124[15:0];
  assign myMuxes_io_counterMatrix1_5_6 = _GEN_125[15:0];
  assign myMuxes_io_counterMatrix1_5_7 = _GEN_126[15:0];
  assign myMuxes_io_counterMatrix1_6_0 = _GEN_127[15:0];
  assign myMuxes_io_counterMatrix1_6_1 = _GEN_128[15:0];
  assign myMuxes_io_counterMatrix1_6_2 = _GEN_129[15:0];
  assign myMuxes_io_counterMatrix1_6_3 = _GEN_130[15:0];
  assign myMuxes_io_counterMatrix1_6_4 = _GEN_131[15:0];
  assign myMuxes_io_counterMatrix1_6_5 = _GEN_132[15:0];
  assign myMuxes_io_counterMatrix1_6_6 = _GEN_133[15:0];
  assign myMuxes_io_counterMatrix1_6_7 = _GEN_134[15:0];
  assign myMuxes_io_counterMatrix1_7_0 = _GEN_135[15:0];
  assign myMuxes_io_counterMatrix1_7_1 = _GEN_136[15:0];
  assign myMuxes_io_counterMatrix1_7_2 = _GEN_137[15:0];
  assign myMuxes_io_counterMatrix1_7_3 = _GEN_138[15:0];
  assign myMuxes_io_counterMatrix1_7_4 = _GEN_139[15:0];
  assign myMuxes_io_counterMatrix1_7_5 = _GEN_140[15:0];
  assign myMuxes_io_counterMatrix1_7_6 = _GEN_141[15:0];
  assign myMuxes_io_counterMatrix1_7_7 = _GEN_142[15:0];
  assign myMuxes_io_counterMatrix2_0 = Distribution_io_ProcessValid ? myCounter_io_counterMatrix2_bits_0 : 16'h0; // @[PathFinder.scala 65:40 72:31 81:31]
  assign myMuxes_io_counterMatrix2_1 = Distribution_io_ProcessValid ? myCounter_io_counterMatrix2_bits_1 : 16'h0; // @[PathFinder.scala 65:40 72:31 81:31]
  assign myMuxes_io_counterMatrix2_2 = Distribution_io_ProcessValid ? myCounter_io_counterMatrix2_bits_2 : 16'h0; // @[PathFinder.scala 65:40 72:31 81:31]
  assign myMuxes_io_counterMatrix2_3 = Distribution_io_ProcessValid ? myCounter_io_counterMatrix2_bits_3 : 16'h0; // @[PathFinder.scala 65:40 72:31 81:31]
  assign myMuxes_io_counterMatrix2_4 = Distribution_io_ProcessValid ? myCounter_io_counterMatrix2_bits_4 : 16'h0; // @[PathFinder.scala 65:40 72:31 81:31]
  assign myMuxes_io_counterMatrix2_5 = Distribution_io_ProcessValid ? myCounter_io_counterMatrix2_bits_5 : 16'h0; // @[PathFinder.scala 65:40 72:31 81:31]
  assign myMuxes_io_counterMatrix2_6 = Distribution_io_ProcessValid ? myCounter_io_counterMatrix2_bits_6 : 16'h0; // @[PathFinder.scala 65:40 72:31 81:31]
  assign myMuxes_io_counterMatrix2_7 = Distribution_io_ProcessValid ? myCounter_io_counterMatrix2_bits_7 : 16'h0; // @[PathFinder.scala 65:40 72:31 81:31]
  assign myCounter_clock = clock;
  assign myCounter_reset = reset;
  assign myCounter_io_Stationary_matrix_0_0 = io_Stationary_matrix_0_0; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_0_1 = io_Stationary_matrix_0_1; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_0_2 = io_Stationary_matrix_0_2; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_0_3 = io_Stationary_matrix_0_3; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_0_4 = io_Stationary_matrix_0_4; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_0_5 = io_Stationary_matrix_0_5; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_0_6 = io_Stationary_matrix_0_6; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_0_7 = io_Stationary_matrix_0_7; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_1_0 = io_Stationary_matrix_1_0; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_1_1 = io_Stationary_matrix_1_1; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_1_2 = io_Stationary_matrix_1_2; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_1_3 = io_Stationary_matrix_1_3; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_1_4 = io_Stationary_matrix_1_4; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_1_5 = io_Stationary_matrix_1_5; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_1_6 = io_Stationary_matrix_1_6; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_1_7 = io_Stationary_matrix_1_7; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_2_0 = io_Stationary_matrix_2_0; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_2_1 = io_Stationary_matrix_2_1; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_2_2 = io_Stationary_matrix_2_2; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_2_3 = io_Stationary_matrix_2_3; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_2_4 = io_Stationary_matrix_2_4; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_2_5 = io_Stationary_matrix_2_5; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_2_6 = io_Stationary_matrix_2_6; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_2_7 = io_Stationary_matrix_2_7; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_3_0 = io_Stationary_matrix_3_0; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_3_1 = io_Stationary_matrix_3_1; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_3_2 = io_Stationary_matrix_3_2; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_3_3 = io_Stationary_matrix_3_3; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_3_4 = io_Stationary_matrix_3_4; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_3_5 = io_Stationary_matrix_3_5; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_3_6 = io_Stationary_matrix_3_6; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_3_7 = io_Stationary_matrix_3_7; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_4_0 = io_Stationary_matrix_4_0; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_4_1 = io_Stationary_matrix_4_1; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_4_2 = io_Stationary_matrix_4_2; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_4_3 = io_Stationary_matrix_4_3; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_4_4 = io_Stationary_matrix_4_4; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_4_5 = io_Stationary_matrix_4_5; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_4_6 = io_Stationary_matrix_4_6; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_4_7 = io_Stationary_matrix_4_7; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_5_0 = io_Stationary_matrix_5_0; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_5_1 = io_Stationary_matrix_5_1; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_5_2 = io_Stationary_matrix_5_2; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_5_3 = io_Stationary_matrix_5_3; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_5_4 = io_Stationary_matrix_5_4; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_5_5 = io_Stationary_matrix_5_5; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_5_6 = io_Stationary_matrix_5_6; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_5_7 = io_Stationary_matrix_5_7; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_6_0 = io_Stationary_matrix_6_0; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_6_1 = io_Stationary_matrix_6_1; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_6_2 = io_Stationary_matrix_6_2; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_6_3 = io_Stationary_matrix_6_3; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_6_4 = io_Stationary_matrix_6_4; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_6_5 = io_Stationary_matrix_6_5; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_6_6 = io_Stationary_matrix_6_6; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_6_7 = io_Stationary_matrix_6_7; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_7_0 = io_Stationary_matrix_7_0; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_7_1 = io_Stationary_matrix_7_1; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_7_2 = io_Stationary_matrix_7_2; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_7_3 = io_Stationary_matrix_7_3; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_7_4 = io_Stationary_matrix_7_4; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_7_5 = io_Stationary_matrix_7_5; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_7_6 = io_Stationary_matrix_7_6; // @[PathFinder.scala 33:34]
  assign myCounter_io_Stationary_matrix_7_7 = io_Stationary_matrix_7_7; // @[PathFinder.scala 33:34]
  assign myCounter_io_Streaming_matrix_0 = io_Streaming_matrix_0; // @[PathFinder.scala 34:33]
  assign myCounter_io_Streaming_matrix_1 = io_Streaming_matrix_1; // @[PathFinder.scala 34:33]
  assign myCounter_io_Streaming_matrix_2 = io_Streaming_matrix_2; // @[PathFinder.scala 34:33]
  assign myCounter_io_Streaming_matrix_3 = io_Streaming_matrix_3; // @[PathFinder.scala 34:33]
  assign myCounter_io_Streaming_matrix_4 = io_Streaming_matrix_4; // @[PathFinder.scala 34:33]
  assign myCounter_io_Streaming_matrix_5 = io_Streaming_matrix_5; // @[PathFinder.scala 34:33]
  assign myCounter_io_Streaming_matrix_6 = io_Streaming_matrix_6; // @[PathFinder.scala 34:33]
  assign myCounter_io_Streaming_matrix_7 = io_Streaming_matrix_7; // @[PathFinder.scala 34:33]
  assign myCounter_io_start = myCounter_io_start_REG; // @[PathFinder.scala 32:22]
  assign Distribution_clock = clock;
  assign Distribution_reset = reset;
  assign Distribution_io_matrix_0_0 = {{16'd0}, myCounter_io_counterMatrix1_bits_0_0}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_0_1 = {{16'd0}, myCounter_io_counterMatrix1_bits_0_1}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_0_2 = {{16'd0}, myCounter_io_counterMatrix1_bits_0_2}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_0_3 = {{16'd0}, myCounter_io_counterMatrix1_bits_0_3}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_0_4 = {{16'd0}, myCounter_io_counterMatrix1_bits_0_4}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_0_5 = {{16'd0}, myCounter_io_counterMatrix1_bits_0_5}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_0_6 = {{16'd0}, myCounter_io_counterMatrix1_bits_0_6}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_0_7 = {{16'd0}, myCounter_io_counterMatrix1_bits_0_7}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_1_0 = {{16'd0}, myCounter_io_counterMatrix1_bits_1_0}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_1_1 = {{16'd0}, myCounter_io_counterMatrix1_bits_1_1}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_1_2 = {{16'd0}, myCounter_io_counterMatrix1_bits_1_2}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_1_3 = {{16'd0}, myCounter_io_counterMatrix1_bits_1_3}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_1_4 = {{16'd0}, myCounter_io_counterMatrix1_bits_1_4}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_1_5 = {{16'd0}, myCounter_io_counterMatrix1_bits_1_5}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_1_6 = {{16'd0}, myCounter_io_counterMatrix1_bits_1_6}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_1_7 = {{16'd0}, myCounter_io_counterMatrix1_bits_1_7}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_2_0 = {{16'd0}, myCounter_io_counterMatrix1_bits_2_0}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_2_1 = {{16'd0}, myCounter_io_counterMatrix1_bits_2_1}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_2_2 = {{16'd0}, myCounter_io_counterMatrix1_bits_2_2}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_2_3 = {{16'd0}, myCounter_io_counterMatrix1_bits_2_3}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_2_4 = {{16'd0}, myCounter_io_counterMatrix1_bits_2_4}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_2_5 = {{16'd0}, myCounter_io_counterMatrix1_bits_2_5}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_2_6 = {{16'd0}, myCounter_io_counterMatrix1_bits_2_6}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_2_7 = {{16'd0}, myCounter_io_counterMatrix1_bits_2_7}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_3_0 = {{16'd0}, myCounter_io_counterMatrix1_bits_3_0}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_3_1 = {{16'd0}, myCounter_io_counterMatrix1_bits_3_1}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_3_2 = {{16'd0}, myCounter_io_counterMatrix1_bits_3_2}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_3_3 = {{16'd0}, myCounter_io_counterMatrix1_bits_3_3}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_3_4 = {{16'd0}, myCounter_io_counterMatrix1_bits_3_4}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_3_5 = {{16'd0}, myCounter_io_counterMatrix1_bits_3_5}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_3_6 = {{16'd0}, myCounter_io_counterMatrix1_bits_3_6}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_3_7 = {{16'd0}, myCounter_io_counterMatrix1_bits_3_7}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_4_0 = {{16'd0}, myCounter_io_counterMatrix1_bits_4_0}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_4_1 = {{16'd0}, myCounter_io_counterMatrix1_bits_4_1}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_4_2 = {{16'd0}, myCounter_io_counterMatrix1_bits_4_2}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_4_3 = {{16'd0}, myCounter_io_counterMatrix1_bits_4_3}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_4_4 = {{16'd0}, myCounter_io_counterMatrix1_bits_4_4}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_4_5 = {{16'd0}, myCounter_io_counterMatrix1_bits_4_5}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_4_6 = {{16'd0}, myCounter_io_counterMatrix1_bits_4_6}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_4_7 = {{16'd0}, myCounter_io_counterMatrix1_bits_4_7}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_5_0 = {{16'd0}, myCounter_io_counterMatrix1_bits_5_0}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_5_1 = {{16'd0}, myCounter_io_counterMatrix1_bits_5_1}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_5_2 = {{16'd0}, myCounter_io_counterMatrix1_bits_5_2}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_5_3 = {{16'd0}, myCounter_io_counterMatrix1_bits_5_3}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_5_4 = {{16'd0}, myCounter_io_counterMatrix1_bits_5_4}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_5_5 = {{16'd0}, myCounter_io_counterMatrix1_bits_5_5}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_5_6 = {{16'd0}, myCounter_io_counterMatrix1_bits_5_6}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_5_7 = {{16'd0}, myCounter_io_counterMatrix1_bits_5_7}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_6_0 = {{16'd0}, myCounter_io_counterMatrix1_bits_6_0}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_6_1 = {{16'd0}, myCounter_io_counterMatrix1_bits_6_1}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_6_2 = {{16'd0}, myCounter_io_counterMatrix1_bits_6_2}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_6_3 = {{16'd0}, myCounter_io_counterMatrix1_bits_6_3}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_6_4 = {{16'd0}, myCounter_io_counterMatrix1_bits_6_4}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_6_5 = {{16'd0}, myCounter_io_counterMatrix1_bits_6_5}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_6_6 = {{16'd0}, myCounter_io_counterMatrix1_bits_6_6}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_6_7 = {{16'd0}, myCounter_io_counterMatrix1_bits_6_7}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_7_0 = {{16'd0}, myCounter_io_counterMatrix1_bits_7_0}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_7_1 = {{16'd0}, myCounter_io_counterMatrix1_bits_7_1}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_7_2 = {{16'd0}, myCounter_io_counterMatrix1_bits_7_2}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_7_3 = {{16'd0}, myCounter_io_counterMatrix1_bits_7_3}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_7_4 = {{16'd0}, myCounter_io_counterMatrix1_bits_7_4}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_7_5 = {{16'd0}, myCounter_io_counterMatrix1_bits_7_5}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_7_6 = {{16'd0}, myCounter_io_counterMatrix1_bits_7_6}; // @[PathFinder.scala 56:26]
  assign Distribution_io_matrix_7_7 = {{16'd0}, myCounter_io_counterMatrix1_bits_7_7}; // @[PathFinder.scala 56:26]
  assign Distribution_io_s = io_NoDPE; // @[PathFinder.scala 53:21]
  assign Distribution_io_valid = high; // @[PathFinder.scala 52:25]
  always @(posedge clock) begin
    if (reset) begin // @[PathFinder.scala 24:22]
      delay <= 32'h0; // @[PathFinder.scala 24:22]
    end else if (!(myCounter_io_valid)) begin // @[PathFinder.scala 39:28]
      if (delay < 32'h40 & high2) begin // @[PathFinder.scala 41:72]
        delay <= _delay_T_1; // @[PathFinder.scala 42:11]
      end
    end
    if (reset) begin // @[PathFinder.scala 26:21]
      high <= 1'h0; // @[PathFinder.scala 26:21]
    end else if (!(myCounter_io_valid)) begin // @[PathFinder.scala 39:28]
      high <= _T_1;
    end
    myCounter_io_start_REG <= io_DataValid; // @[PathFinder.scala 32:32]
    if (reset) begin // @[PathFinder.scala 36:22]
      high2 <= 1'h0; // @[PathFinder.scala 36:22]
    end else begin
      high2 <= _GEN_3;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  delay = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  high = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  myCounter_io_start_REG = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  high2 = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module stationary(
  input         clock,
  input         reset,
  input  [15:0] io_Stationary_matrix_0_0,
  input  [15:0] io_Stationary_matrix_0_1,
  input  [15:0] io_Stationary_matrix_0_2,
  input  [15:0] io_Stationary_matrix_0_3,
  input  [15:0] io_Stationary_matrix_0_4,
  input  [15:0] io_Stationary_matrix_0_5,
  input  [15:0] io_Stationary_matrix_0_6,
  input  [15:0] io_Stationary_matrix_0_7,
  input  [15:0] io_Stationary_matrix_1_0,
  input  [15:0] io_Stationary_matrix_1_1,
  input  [15:0] io_Stationary_matrix_1_2,
  input  [15:0] io_Stationary_matrix_1_3,
  input  [15:0] io_Stationary_matrix_1_4,
  input  [15:0] io_Stationary_matrix_1_5,
  input  [15:0] io_Stationary_matrix_1_6,
  input  [15:0] io_Stationary_matrix_1_7,
  input  [15:0] io_Stationary_matrix_2_0,
  input  [15:0] io_Stationary_matrix_2_1,
  input  [15:0] io_Stationary_matrix_2_2,
  input  [15:0] io_Stationary_matrix_2_3,
  input  [15:0] io_Stationary_matrix_2_4,
  input  [15:0] io_Stationary_matrix_2_5,
  input  [15:0] io_Stationary_matrix_2_6,
  input  [15:0] io_Stationary_matrix_2_7,
  input  [15:0] io_Stationary_matrix_3_0,
  input  [15:0] io_Stationary_matrix_3_1,
  input  [15:0] io_Stationary_matrix_3_2,
  input  [15:0] io_Stationary_matrix_3_3,
  input  [15:0] io_Stationary_matrix_3_4,
  input  [15:0] io_Stationary_matrix_3_5,
  input  [15:0] io_Stationary_matrix_3_6,
  input  [15:0] io_Stationary_matrix_3_7,
  input  [15:0] io_Stationary_matrix_4_0,
  input  [15:0] io_Stationary_matrix_4_1,
  input  [15:0] io_Stationary_matrix_4_2,
  input  [15:0] io_Stationary_matrix_4_3,
  input  [15:0] io_Stationary_matrix_4_4,
  input  [15:0] io_Stationary_matrix_4_5,
  input  [15:0] io_Stationary_matrix_4_6,
  input  [15:0] io_Stationary_matrix_4_7,
  input  [15:0] io_Stationary_matrix_5_0,
  input  [15:0] io_Stationary_matrix_5_1,
  input  [15:0] io_Stationary_matrix_5_2,
  input  [15:0] io_Stationary_matrix_5_3,
  input  [15:0] io_Stationary_matrix_5_4,
  input  [15:0] io_Stationary_matrix_5_5,
  input  [15:0] io_Stationary_matrix_5_6,
  input  [15:0] io_Stationary_matrix_5_7,
  input  [15:0] io_Stationary_matrix_6_0,
  input  [15:0] io_Stationary_matrix_6_1,
  input  [15:0] io_Stationary_matrix_6_2,
  input  [15:0] io_Stationary_matrix_6_3,
  input  [15:0] io_Stationary_matrix_6_4,
  input  [15:0] io_Stationary_matrix_6_5,
  input  [15:0] io_Stationary_matrix_6_6,
  input  [15:0] io_Stationary_matrix_6_7,
  input  [15:0] io_Stationary_matrix_7_0,
  input  [15:0] io_Stationary_matrix_7_1,
  input  [15:0] io_Stationary_matrix_7_2,
  input  [15:0] io_Stationary_matrix_7_3,
  input  [15:0] io_Stationary_matrix_7_4,
  input  [15:0] io_Stationary_matrix_7_5,
  input  [15:0] io_Stationary_matrix_7_6,
  input  [15:0] io_Stationary_matrix_7_7,
  output [15:0] io_o_Stationary_matrix1_0_0,
  output [15:0] io_o_Stationary_matrix1_0_1,
  output [15:0] io_o_Stationary_matrix1_0_2,
  output [15:0] io_o_Stationary_matrix1_0_3,
  output [15:0] io_o_Stationary_matrix1_0_4,
  output [15:0] io_o_Stationary_matrix1_0_5,
  output [15:0] io_o_Stationary_matrix1_0_6,
  output [15:0] io_o_Stationary_matrix1_0_7,
  output [15:0] io_o_Stationary_matrix1_1_0,
  output [15:0] io_o_Stationary_matrix1_1_1,
  output [15:0] io_o_Stationary_matrix1_1_2,
  output [15:0] io_o_Stationary_matrix1_1_3,
  output [15:0] io_o_Stationary_matrix1_1_4,
  output [15:0] io_o_Stationary_matrix1_1_5,
  output [15:0] io_o_Stationary_matrix1_1_6,
  output [15:0] io_o_Stationary_matrix1_1_7,
  output [15:0] io_o_Stationary_matrix1_2_0,
  output [15:0] io_o_Stationary_matrix1_2_1,
  output [15:0] io_o_Stationary_matrix1_2_2,
  output [15:0] io_o_Stationary_matrix1_2_3,
  output [15:0] io_o_Stationary_matrix1_2_4,
  output [15:0] io_o_Stationary_matrix1_2_5,
  output [15:0] io_o_Stationary_matrix1_2_6,
  output [15:0] io_o_Stationary_matrix1_2_7,
  output [15:0] io_o_Stationary_matrix1_3_0,
  output [15:0] io_o_Stationary_matrix1_3_1,
  output [15:0] io_o_Stationary_matrix1_3_2,
  output [15:0] io_o_Stationary_matrix1_3_3,
  output [15:0] io_o_Stationary_matrix1_3_4,
  output [15:0] io_o_Stationary_matrix1_3_5,
  output [15:0] io_o_Stationary_matrix1_3_6,
  output [15:0] io_o_Stationary_matrix1_3_7,
  output [15:0] io_o_Stationary_matrix1_4_0,
  output [15:0] io_o_Stationary_matrix1_4_1,
  output [15:0] io_o_Stationary_matrix1_4_2,
  output [15:0] io_o_Stationary_matrix1_4_3,
  output [15:0] io_o_Stationary_matrix1_4_4,
  output [15:0] io_o_Stationary_matrix1_4_5,
  output [15:0] io_o_Stationary_matrix1_4_6,
  output [15:0] io_o_Stationary_matrix1_4_7,
  output [15:0] io_o_Stationary_matrix1_5_0,
  output [15:0] io_o_Stationary_matrix1_5_1,
  output [15:0] io_o_Stationary_matrix1_5_2,
  output [15:0] io_o_Stationary_matrix1_5_3,
  output [15:0] io_o_Stationary_matrix1_5_4,
  output [15:0] io_o_Stationary_matrix1_5_5,
  output [15:0] io_o_Stationary_matrix1_5_6,
  output [15:0] io_o_Stationary_matrix1_5_7,
  output [15:0] io_o_Stationary_matrix1_6_0,
  output [15:0] io_o_Stationary_matrix1_6_1,
  output [15:0] io_o_Stationary_matrix1_6_2,
  output [15:0] io_o_Stationary_matrix1_6_3,
  output [15:0] io_o_Stationary_matrix1_6_4,
  output [15:0] io_o_Stationary_matrix1_6_5,
  output [15:0] io_o_Stationary_matrix1_6_6,
  output [15:0] io_o_Stationary_matrix1_6_7,
  output [15:0] io_o_Stationary_matrix1_7_0,
  output [15:0] io_o_Stationary_matrix1_7_1,
  output [15:0] io_o_Stationary_matrix1_7_2,
  output [15:0] io_o_Stationary_matrix1_7_3,
  output [15:0] io_o_Stationary_matrix1_7_4,
  output [15:0] io_o_Stationary_matrix1_7_5,
  output [15:0] io_o_Stationary_matrix1_7_6,
  output [15:0] io_o_Stationary_matrix1_7_7,
  output [15:0] io_o_Stationary_matrix2_0_0,
  output [15:0] io_o_Stationary_matrix2_0_1,
  output [15:0] io_o_Stationary_matrix2_0_2,
  output [15:0] io_o_Stationary_matrix2_0_3,
  output [15:0] io_o_Stationary_matrix2_0_4,
  output [15:0] io_o_Stationary_matrix2_0_5,
  output [15:0] io_o_Stationary_matrix2_0_6,
  output [15:0] io_o_Stationary_matrix2_0_7,
  output [15:0] io_o_Stationary_matrix2_1_0,
  output [15:0] io_o_Stationary_matrix2_1_1,
  output [15:0] io_o_Stationary_matrix2_1_2,
  output [15:0] io_o_Stationary_matrix2_1_3,
  output [15:0] io_o_Stationary_matrix2_1_4,
  output [15:0] io_o_Stationary_matrix2_1_5,
  output [15:0] io_o_Stationary_matrix2_1_6,
  output [15:0] io_o_Stationary_matrix2_1_7,
  output [15:0] io_o_Stationary_matrix2_2_0,
  output [15:0] io_o_Stationary_matrix2_2_1,
  output [15:0] io_o_Stationary_matrix2_2_2,
  output [15:0] io_o_Stationary_matrix2_2_3,
  output [15:0] io_o_Stationary_matrix2_2_4,
  output [15:0] io_o_Stationary_matrix2_2_5,
  output [15:0] io_o_Stationary_matrix2_2_6,
  output [15:0] io_o_Stationary_matrix2_2_7,
  output [15:0] io_o_Stationary_matrix2_3_0,
  output [15:0] io_o_Stationary_matrix2_3_1,
  output [15:0] io_o_Stationary_matrix2_3_2,
  output [15:0] io_o_Stationary_matrix2_3_3,
  output [15:0] io_o_Stationary_matrix2_3_4,
  output [15:0] io_o_Stationary_matrix2_3_5,
  output [15:0] io_o_Stationary_matrix2_3_6,
  output [15:0] io_o_Stationary_matrix2_3_7,
  output [15:0] io_o_Stationary_matrix2_4_0,
  output [15:0] io_o_Stationary_matrix2_4_1,
  output [15:0] io_o_Stationary_matrix2_4_2,
  output [15:0] io_o_Stationary_matrix2_4_3,
  output [15:0] io_o_Stationary_matrix2_4_4,
  output [15:0] io_o_Stationary_matrix2_4_5,
  output [15:0] io_o_Stationary_matrix2_4_6,
  output [15:0] io_o_Stationary_matrix2_4_7,
  output [15:0] io_o_Stationary_matrix2_5_0,
  output [15:0] io_o_Stationary_matrix2_5_1,
  output [15:0] io_o_Stationary_matrix2_5_2,
  output [15:0] io_o_Stationary_matrix2_5_3,
  output [15:0] io_o_Stationary_matrix2_5_4,
  output [15:0] io_o_Stationary_matrix2_5_5,
  output [15:0] io_o_Stationary_matrix2_5_6,
  output [15:0] io_o_Stationary_matrix2_5_7,
  output [15:0] io_o_Stationary_matrix2_6_0,
  output [15:0] io_o_Stationary_matrix2_6_1,
  output [15:0] io_o_Stationary_matrix2_6_2,
  output [15:0] io_o_Stationary_matrix2_6_3,
  output [15:0] io_o_Stationary_matrix2_6_4,
  output [15:0] io_o_Stationary_matrix2_6_5,
  output [15:0] io_o_Stationary_matrix2_6_6,
  output [15:0] io_o_Stationary_matrix2_6_7,
  output [15:0] io_o_Stationary_matrix2_7_0,
  output [15:0] io_o_Stationary_matrix2_7_1,
  output [15:0] io_o_Stationary_matrix2_7_2,
  output [15:0] io_o_Stationary_matrix2_7_3,
  output [15:0] io_o_Stationary_matrix2_7_4,
  output [15:0] io_o_Stationary_matrix2_7_5,
  output [15:0] io_o_Stationary_matrix2_7_6,
  output [15:0] io_o_Stationary_matrix2_7_7,
  output [15:0] io_o_Stationary_matrix3_0_0,
  output [15:0] io_o_Stationary_matrix3_0_1,
  output [15:0] io_o_Stationary_matrix3_0_2,
  output [15:0] io_o_Stationary_matrix3_0_3,
  output [15:0] io_o_Stationary_matrix3_0_4,
  output [15:0] io_o_Stationary_matrix3_0_5,
  output [15:0] io_o_Stationary_matrix3_0_6,
  output [15:0] io_o_Stationary_matrix3_0_7,
  output [15:0] io_o_Stationary_matrix3_1_0,
  output [15:0] io_o_Stationary_matrix3_1_1,
  output [15:0] io_o_Stationary_matrix3_1_2,
  output [15:0] io_o_Stationary_matrix3_1_3,
  output [15:0] io_o_Stationary_matrix3_1_4,
  output [15:0] io_o_Stationary_matrix3_1_5,
  output [15:0] io_o_Stationary_matrix3_1_6,
  output [15:0] io_o_Stationary_matrix3_1_7,
  output [15:0] io_o_Stationary_matrix3_2_0,
  output [15:0] io_o_Stationary_matrix3_2_1,
  output [15:0] io_o_Stationary_matrix3_2_2,
  output [15:0] io_o_Stationary_matrix3_2_3,
  output [15:0] io_o_Stationary_matrix3_2_4,
  output [15:0] io_o_Stationary_matrix3_2_5,
  output [15:0] io_o_Stationary_matrix3_2_6,
  output [15:0] io_o_Stationary_matrix3_2_7,
  output [15:0] io_o_Stationary_matrix3_3_0,
  output [15:0] io_o_Stationary_matrix3_3_1,
  output [15:0] io_o_Stationary_matrix3_3_2,
  output [15:0] io_o_Stationary_matrix3_3_3,
  output [15:0] io_o_Stationary_matrix3_3_4,
  output [15:0] io_o_Stationary_matrix3_3_5,
  output [15:0] io_o_Stationary_matrix3_3_6,
  output [15:0] io_o_Stationary_matrix3_3_7,
  output [15:0] io_o_Stationary_matrix3_4_0,
  output [15:0] io_o_Stationary_matrix3_4_1,
  output [15:0] io_o_Stationary_matrix3_4_2,
  output [15:0] io_o_Stationary_matrix3_4_3,
  output [15:0] io_o_Stationary_matrix3_4_4,
  output [15:0] io_o_Stationary_matrix3_4_5,
  output [15:0] io_o_Stationary_matrix3_4_6,
  output [15:0] io_o_Stationary_matrix3_4_7,
  output [15:0] io_o_Stationary_matrix3_5_0,
  output [15:0] io_o_Stationary_matrix3_5_1,
  output [15:0] io_o_Stationary_matrix3_5_2,
  output [15:0] io_o_Stationary_matrix3_5_3,
  output [15:0] io_o_Stationary_matrix3_5_4,
  output [15:0] io_o_Stationary_matrix3_5_5,
  output [15:0] io_o_Stationary_matrix3_5_6,
  output [15:0] io_o_Stationary_matrix3_5_7,
  output [15:0] io_o_Stationary_matrix3_6_0,
  output [15:0] io_o_Stationary_matrix3_6_1,
  output [15:0] io_o_Stationary_matrix3_6_2,
  output [15:0] io_o_Stationary_matrix3_6_3,
  output [15:0] io_o_Stationary_matrix3_6_4,
  output [15:0] io_o_Stationary_matrix3_6_5,
  output [15:0] io_o_Stationary_matrix3_6_6,
  output [15:0] io_o_Stationary_matrix3_6_7,
  output [15:0] io_o_Stationary_matrix3_7_0,
  output [15:0] io_o_Stationary_matrix3_7_1,
  output [15:0] io_o_Stationary_matrix3_7_2,
  output [15:0] io_o_Stationary_matrix3_7_3,
  output [15:0] io_o_Stationary_matrix3_7_4,
  output [15:0] io_o_Stationary_matrix3_7_5,
  output [15:0] io_o_Stationary_matrix3_7_6,
  output [15:0] io_o_Stationary_matrix3_7_7,
  output [15:0] io_o_Stationary_matrix4_0_0,
  output [15:0] io_o_Stationary_matrix4_0_1,
  output [15:0] io_o_Stationary_matrix4_0_2,
  output [15:0] io_o_Stationary_matrix4_0_3,
  output [15:0] io_o_Stationary_matrix4_0_4,
  output [15:0] io_o_Stationary_matrix4_0_5,
  output [15:0] io_o_Stationary_matrix4_0_6,
  output [15:0] io_o_Stationary_matrix4_0_7,
  output [15:0] io_o_Stationary_matrix4_1_0,
  output [15:0] io_o_Stationary_matrix4_1_1,
  output [15:0] io_o_Stationary_matrix4_1_2,
  output [15:0] io_o_Stationary_matrix4_1_3,
  output [15:0] io_o_Stationary_matrix4_1_4,
  output [15:0] io_o_Stationary_matrix4_1_5,
  output [15:0] io_o_Stationary_matrix4_1_6,
  output [15:0] io_o_Stationary_matrix4_1_7,
  output [15:0] io_o_Stationary_matrix4_2_0,
  output [15:0] io_o_Stationary_matrix4_2_1,
  output [15:0] io_o_Stationary_matrix4_2_2,
  output [15:0] io_o_Stationary_matrix4_2_3,
  output [15:0] io_o_Stationary_matrix4_2_4,
  output [15:0] io_o_Stationary_matrix4_2_5,
  output [15:0] io_o_Stationary_matrix4_2_6,
  output [15:0] io_o_Stationary_matrix4_2_7,
  output [15:0] io_o_Stationary_matrix4_3_0,
  output [15:0] io_o_Stationary_matrix4_3_1,
  output [15:0] io_o_Stationary_matrix4_3_2,
  output [15:0] io_o_Stationary_matrix4_3_3,
  output [15:0] io_o_Stationary_matrix4_3_4,
  output [15:0] io_o_Stationary_matrix4_3_5,
  output [15:0] io_o_Stationary_matrix4_3_6,
  output [15:0] io_o_Stationary_matrix4_3_7,
  output [15:0] io_o_Stationary_matrix4_4_0,
  output [15:0] io_o_Stationary_matrix4_4_1,
  output [15:0] io_o_Stationary_matrix4_4_2,
  output [15:0] io_o_Stationary_matrix4_4_3,
  output [15:0] io_o_Stationary_matrix4_4_4,
  output [15:0] io_o_Stationary_matrix4_4_5,
  output [15:0] io_o_Stationary_matrix4_4_6,
  output [15:0] io_o_Stationary_matrix4_4_7,
  output [15:0] io_o_Stationary_matrix4_5_0,
  output [15:0] io_o_Stationary_matrix4_5_1,
  output [15:0] io_o_Stationary_matrix4_5_2,
  output [15:0] io_o_Stationary_matrix4_5_3,
  output [15:0] io_o_Stationary_matrix4_5_4,
  output [15:0] io_o_Stationary_matrix4_5_5,
  output [15:0] io_o_Stationary_matrix4_5_6,
  output [15:0] io_o_Stationary_matrix4_5_7,
  output [15:0] io_o_Stationary_matrix4_6_0,
  output [15:0] io_o_Stationary_matrix4_6_1,
  output [15:0] io_o_Stationary_matrix4_6_2,
  output [15:0] io_o_Stationary_matrix4_6_3,
  output [15:0] io_o_Stationary_matrix4_6_4,
  output [15:0] io_o_Stationary_matrix4_6_5,
  output [15:0] io_o_Stationary_matrix4_6_6,
  output [15:0] io_o_Stationary_matrix4_6_7,
  output [15:0] io_o_Stationary_matrix4_7_0,
  output [15:0] io_o_Stationary_matrix4_7_1,
  output [15:0] io_o_Stationary_matrix4_7_2,
  output [15:0] io_o_Stationary_matrix4_7_3,
  output [15:0] io_o_Stationary_matrix4_7_4,
  output [15:0] io_o_Stationary_matrix4_7_5,
  output [15:0] io_o_Stationary_matrix4_7_6,
  output [15:0] io_o_Stationary_matrix4_7_7,
  output [15:0] io_o_Stationary_matrix5_0_0,
  output [15:0] io_o_Stationary_matrix5_0_1,
  output [15:0] io_o_Stationary_matrix5_0_2,
  output [15:0] io_o_Stationary_matrix5_0_3,
  output [15:0] io_o_Stationary_matrix5_0_4,
  output [15:0] io_o_Stationary_matrix5_0_5,
  output [15:0] io_o_Stationary_matrix5_0_6,
  output [15:0] io_o_Stationary_matrix5_0_7,
  output [15:0] io_o_Stationary_matrix5_1_0,
  output [15:0] io_o_Stationary_matrix5_1_1,
  output [15:0] io_o_Stationary_matrix5_1_2,
  output [15:0] io_o_Stationary_matrix5_1_3,
  output [15:0] io_o_Stationary_matrix5_1_4,
  output [15:0] io_o_Stationary_matrix5_1_5,
  output [15:0] io_o_Stationary_matrix5_1_6,
  output [15:0] io_o_Stationary_matrix5_1_7,
  output [15:0] io_o_Stationary_matrix5_2_0,
  output [15:0] io_o_Stationary_matrix5_2_1,
  output [15:0] io_o_Stationary_matrix5_2_2,
  output [15:0] io_o_Stationary_matrix5_2_3,
  output [15:0] io_o_Stationary_matrix5_2_4,
  output [15:0] io_o_Stationary_matrix5_2_5,
  output [15:0] io_o_Stationary_matrix5_2_6,
  output [15:0] io_o_Stationary_matrix5_2_7,
  output [15:0] io_o_Stationary_matrix5_3_0,
  output [15:0] io_o_Stationary_matrix5_3_1,
  output [15:0] io_o_Stationary_matrix5_3_2,
  output [15:0] io_o_Stationary_matrix5_3_3,
  output [15:0] io_o_Stationary_matrix5_3_4,
  output [15:0] io_o_Stationary_matrix5_3_5,
  output [15:0] io_o_Stationary_matrix5_3_6,
  output [15:0] io_o_Stationary_matrix5_3_7,
  output [15:0] io_o_Stationary_matrix5_4_0,
  output [15:0] io_o_Stationary_matrix5_4_1,
  output [15:0] io_o_Stationary_matrix5_4_2,
  output [15:0] io_o_Stationary_matrix5_4_3,
  output [15:0] io_o_Stationary_matrix5_4_4,
  output [15:0] io_o_Stationary_matrix5_4_5,
  output [15:0] io_o_Stationary_matrix5_4_6,
  output [15:0] io_o_Stationary_matrix5_4_7,
  output [15:0] io_o_Stationary_matrix5_5_0,
  output [15:0] io_o_Stationary_matrix5_5_1,
  output [15:0] io_o_Stationary_matrix5_5_2,
  output [15:0] io_o_Stationary_matrix5_5_3,
  output [15:0] io_o_Stationary_matrix5_5_4,
  output [15:0] io_o_Stationary_matrix5_5_5,
  output [15:0] io_o_Stationary_matrix5_5_6,
  output [15:0] io_o_Stationary_matrix5_5_7,
  output [15:0] io_o_Stationary_matrix5_6_0,
  output [15:0] io_o_Stationary_matrix5_6_1,
  output [15:0] io_o_Stationary_matrix5_6_2,
  output [15:0] io_o_Stationary_matrix5_6_3,
  output [15:0] io_o_Stationary_matrix5_6_4,
  output [15:0] io_o_Stationary_matrix5_6_5,
  output [15:0] io_o_Stationary_matrix5_6_6,
  output [15:0] io_o_Stationary_matrix5_6_7,
  output [15:0] io_o_Stationary_matrix5_7_0,
  output [15:0] io_o_Stationary_matrix5_7_1,
  output [15:0] io_o_Stationary_matrix5_7_2,
  output [15:0] io_o_Stationary_matrix5_7_3,
  output [15:0] io_o_Stationary_matrix5_7_4,
  output [15:0] io_o_Stationary_matrix5_7_5,
  output [15:0] io_o_Stationary_matrix5_7_6,
  output [15:0] io_o_Stationary_matrix5_7_7,
  output [15:0] io_o_Stationary_matrix6_0_0,
  output [15:0] io_o_Stationary_matrix6_0_1,
  output [15:0] io_o_Stationary_matrix6_0_2,
  output [15:0] io_o_Stationary_matrix6_0_3,
  output [15:0] io_o_Stationary_matrix6_0_4,
  output [15:0] io_o_Stationary_matrix6_0_5,
  output [15:0] io_o_Stationary_matrix6_0_6,
  output [15:0] io_o_Stationary_matrix6_0_7,
  output [15:0] io_o_Stationary_matrix6_1_0,
  output [15:0] io_o_Stationary_matrix6_1_1,
  output [15:0] io_o_Stationary_matrix6_1_2,
  output [15:0] io_o_Stationary_matrix6_1_3,
  output [15:0] io_o_Stationary_matrix6_1_4,
  output [15:0] io_o_Stationary_matrix6_1_5,
  output [15:0] io_o_Stationary_matrix6_1_6,
  output [15:0] io_o_Stationary_matrix6_1_7,
  output [15:0] io_o_Stationary_matrix6_2_0,
  output [15:0] io_o_Stationary_matrix6_2_1,
  output [15:0] io_o_Stationary_matrix6_2_2,
  output [15:0] io_o_Stationary_matrix6_2_3,
  output [15:0] io_o_Stationary_matrix6_2_4,
  output [15:0] io_o_Stationary_matrix6_2_5,
  output [15:0] io_o_Stationary_matrix6_2_6,
  output [15:0] io_o_Stationary_matrix6_2_7,
  output [15:0] io_o_Stationary_matrix6_3_0,
  output [15:0] io_o_Stationary_matrix6_3_1,
  output [15:0] io_o_Stationary_matrix6_3_2,
  output [15:0] io_o_Stationary_matrix6_3_3,
  output [15:0] io_o_Stationary_matrix6_3_4,
  output [15:0] io_o_Stationary_matrix6_3_5,
  output [15:0] io_o_Stationary_matrix6_3_6,
  output [15:0] io_o_Stationary_matrix6_3_7,
  output [15:0] io_o_Stationary_matrix6_4_0,
  output [15:0] io_o_Stationary_matrix6_4_1,
  output [15:0] io_o_Stationary_matrix6_4_2,
  output [15:0] io_o_Stationary_matrix6_4_3,
  output [15:0] io_o_Stationary_matrix6_4_4,
  output [15:0] io_o_Stationary_matrix6_4_5,
  output [15:0] io_o_Stationary_matrix6_4_6,
  output [15:0] io_o_Stationary_matrix6_4_7,
  output [15:0] io_o_Stationary_matrix6_5_0,
  output [15:0] io_o_Stationary_matrix6_5_1,
  output [15:0] io_o_Stationary_matrix6_5_2,
  output [15:0] io_o_Stationary_matrix6_5_3,
  output [15:0] io_o_Stationary_matrix6_5_4,
  output [15:0] io_o_Stationary_matrix6_5_5,
  output [15:0] io_o_Stationary_matrix6_5_6,
  output [15:0] io_o_Stationary_matrix6_5_7,
  output [15:0] io_o_Stationary_matrix6_6_0,
  output [15:0] io_o_Stationary_matrix6_6_1,
  output [15:0] io_o_Stationary_matrix6_6_2,
  output [15:0] io_o_Stationary_matrix6_6_3,
  output [15:0] io_o_Stationary_matrix6_6_4,
  output [15:0] io_o_Stationary_matrix6_6_5,
  output [15:0] io_o_Stationary_matrix6_6_6,
  output [15:0] io_o_Stationary_matrix6_6_7,
  output [15:0] io_o_Stationary_matrix6_7_0,
  output [15:0] io_o_Stationary_matrix6_7_1,
  output [15:0] io_o_Stationary_matrix6_7_2,
  output [15:0] io_o_Stationary_matrix6_7_3,
  output [15:0] io_o_Stationary_matrix6_7_4,
  output [15:0] io_o_Stationary_matrix6_7_5,
  output [15:0] io_o_Stationary_matrix6_7_6,
  output [15:0] io_o_Stationary_matrix6_7_7,
  output [15:0] io_o_Stationary_matrix7_0_0,
  output [15:0] io_o_Stationary_matrix7_0_1,
  output [15:0] io_o_Stationary_matrix7_0_2,
  output [15:0] io_o_Stationary_matrix7_0_3,
  output [15:0] io_o_Stationary_matrix7_0_4,
  output [15:0] io_o_Stationary_matrix7_0_5,
  output [15:0] io_o_Stationary_matrix7_0_6,
  output [15:0] io_o_Stationary_matrix7_0_7,
  output [15:0] io_o_Stationary_matrix7_1_0,
  output [15:0] io_o_Stationary_matrix7_1_1,
  output [15:0] io_o_Stationary_matrix7_1_2,
  output [15:0] io_o_Stationary_matrix7_1_3,
  output [15:0] io_o_Stationary_matrix7_1_4,
  output [15:0] io_o_Stationary_matrix7_1_5,
  output [15:0] io_o_Stationary_matrix7_1_6,
  output [15:0] io_o_Stationary_matrix7_1_7,
  output [15:0] io_o_Stationary_matrix7_2_0,
  output [15:0] io_o_Stationary_matrix7_2_1,
  output [15:0] io_o_Stationary_matrix7_2_2,
  output [15:0] io_o_Stationary_matrix7_2_3,
  output [15:0] io_o_Stationary_matrix7_2_4,
  output [15:0] io_o_Stationary_matrix7_2_5,
  output [15:0] io_o_Stationary_matrix7_2_6,
  output [15:0] io_o_Stationary_matrix7_2_7,
  output [15:0] io_o_Stationary_matrix7_3_0,
  output [15:0] io_o_Stationary_matrix7_3_1,
  output [15:0] io_o_Stationary_matrix7_3_2,
  output [15:0] io_o_Stationary_matrix7_3_3,
  output [15:0] io_o_Stationary_matrix7_3_4,
  output [15:0] io_o_Stationary_matrix7_3_5,
  output [15:0] io_o_Stationary_matrix7_3_6,
  output [15:0] io_o_Stationary_matrix7_3_7,
  output [15:0] io_o_Stationary_matrix7_4_0,
  output [15:0] io_o_Stationary_matrix7_4_1,
  output [15:0] io_o_Stationary_matrix7_4_2,
  output [15:0] io_o_Stationary_matrix7_4_3,
  output [15:0] io_o_Stationary_matrix7_4_4,
  output [15:0] io_o_Stationary_matrix7_4_5,
  output [15:0] io_o_Stationary_matrix7_4_6,
  output [15:0] io_o_Stationary_matrix7_4_7,
  output [15:0] io_o_Stationary_matrix7_5_0,
  output [15:0] io_o_Stationary_matrix7_5_1,
  output [15:0] io_o_Stationary_matrix7_5_2,
  output [15:0] io_o_Stationary_matrix7_5_3,
  output [15:0] io_o_Stationary_matrix7_5_4,
  output [15:0] io_o_Stationary_matrix7_5_5,
  output [15:0] io_o_Stationary_matrix7_5_6,
  output [15:0] io_o_Stationary_matrix7_5_7,
  output [15:0] io_o_Stationary_matrix7_6_0,
  output [15:0] io_o_Stationary_matrix7_6_1,
  output [15:0] io_o_Stationary_matrix7_6_2,
  output [15:0] io_o_Stationary_matrix7_6_3,
  output [15:0] io_o_Stationary_matrix7_6_4,
  output [15:0] io_o_Stationary_matrix7_6_5,
  output [15:0] io_o_Stationary_matrix7_6_6,
  output [15:0] io_o_Stationary_matrix7_6_7,
  output [15:0] io_o_Stationary_matrix7_7_0,
  output [15:0] io_o_Stationary_matrix7_7_1,
  output [15:0] io_o_Stationary_matrix7_7_2,
  output [15:0] io_o_Stationary_matrix7_7_3,
  output [15:0] io_o_Stationary_matrix7_7_4,
  output [15:0] io_o_Stationary_matrix7_7_5,
  output [15:0] io_o_Stationary_matrix7_7_6,
  output [15:0] io_o_Stationary_matrix7_7_7,
  output [15:0] io_o_Stationary_matrix8_0_0,
  output [15:0] io_o_Stationary_matrix8_0_1,
  output [15:0] io_o_Stationary_matrix8_0_2,
  output [15:0] io_o_Stationary_matrix8_0_3,
  output [15:0] io_o_Stationary_matrix8_0_4,
  output [15:0] io_o_Stationary_matrix8_0_5,
  output [15:0] io_o_Stationary_matrix8_0_6,
  output [15:0] io_o_Stationary_matrix8_0_7,
  output [15:0] io_o_Stationary_matrix8_1_0,
  output [15:0] io_o_Stationary_matrix8_1_1,
  output [15:0] io_o_Stationary_matrix8_1_2,
  output [15:0] io_o_Stationary_matrix8_1_3,
  output [15:0] io_o_Stationary_matrix8_1_4,
  output [15:0] io_o_Stationary_matrix8_1_5,
  output [15:0] io_o_Stationary_matrix8_1_6,
  output [15:0] io_o_Stationary_matrix8_1_7,
  output [15:0] io_o_Stationary_matrix8_2_0,
  output [15:0] io_o_Stationary_matrix8_2_1,
  output [15:0] io_o_Stationary_matrix8_2_2,
  output [15:0] io_o_Stationary_matrix8_2_3,
  output [15:0] io_o_Stationary_matrix8_2_4,
  output [15:0] io_o_Stationary_matrix8_2_5,
  output [15:0] io_o_Stationary_matrix8_2_6,
  output [15:0] io_o_Stationary_matrix8_2_7,
  output [15:0] io_o_Stationary_matrix8_3_0,
  output [15:0] io_o_Stationary_matrix8_3_1,
  output [15:0] io_o_Stationary_matrix8_3_2,
  output [15:0] io_o_Stationary_matrix8_3_3,
  output [15:0] io_o_Stationary_matrix8_3_4,
  output [15:0] io_o_Stationary_matrix8_3_5,
  output [15:0] io_o_Stationary_matrix8_3_6,
  output [15:0] io_o_Stationary_matrix8_3_7,
  output [15:0] io_o_Stationary_matrix8_4_0,
  output [15:0] io_o_Stationary_matrix8_4_1,
  output [15:0] io_o_Stationary_matrix8_4_2,
  output [15:0] io_o_Stationary_matrix8_4_3,
  output [15:0] io_o_Stationary_matrix8_4_4,
  output [15:0] io_o_Stationary_matrix8_4_5,
  output [15:0] io_o_Stationary_matrix8_4_6,
  output [15:0] io_o_Stationary_matrix8_4_7,
  output [15:0] io_o_Stationary_matrix8_5_0,
  output [15:0] io_o_Stationary_matrix8_5_1,
  output [15:0] io_o_Stationary_matrix8_5_2,
  output [15:0] io_o_Stationary_matrix8_5_3,
  output [15:0] io_o_Stationary_matrix8_5_4,
  output [15:0] io_o_Stationary_matrix8_5_5,
  output [15:0] io_o_Stationary_matrix8_5_6,
  output [15:0] io_o_Stationary_matrix8_5_7,
  output [15:0] io_o_Stationary_matrix8_6_0,
  output [15:0] io_o_Stationary_matrix8_6_1,
  output [15:0] io_o_Stationary_matrix8_6_2,
  output [15:0] io_o_Stationary_matrix8_6_3,
  output [15:0] io_o_Stationary_matrix8_6_4,
  output [15:0] io_o_Stationary_matrix8_6_5,
  output [15:0] io_o_Stationary_matrix8_6_6,
  output [15:0] io_o_Stationary_matrix8_6_7,
  output [15:0] io_o_Stationary_matrix8_7_0,
  output [15:0] io_o_Stationary_matrix8_7_1,
  output [15:0] io_o_Stationary_matrix8_7_2,
  output [15:0] io_o_Stationary_matrix8_7_3,
  output [15:0] io_o_Stationary_matrix8_7_4,
  output [15:0] io_o_Stationary_matrix8_7_5,
  output [15:0] io_o_Stationary_matrix8_7_6,
  output [15:0] io_o_Stationary_matrix8_7_7
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] count; // @[stationary_dpe.scala 23:27]
  reg [15:0] Station2_0_0; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_0_1; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_0_2; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_0_3; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_0_4; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_0_5; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_0_6; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_0_7; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_1_0; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_1_1; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_1_2; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_1_3; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_1_4; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_1_5; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_1_6; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_1_7; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_2_0; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_2_1; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_2_2; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_2_3; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_2_4; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_2_5; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_2_6; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_2_7; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_3_0; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_3_1; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_3_2; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_3_3; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_3_4; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_3_5; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_3_6; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_3_7; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_4_0; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_4_1; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_4_2; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_4_3; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_4_4; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_4_5; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_4_6; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_4_7; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_5_0; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_5_1; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_5_2; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_5_3; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_5_4; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_5_5; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_5_6; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_5_7; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_6_0; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_6_1; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_6_2; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_6_3; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_6_4; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_6_5; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_6_6; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_6_7; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_7_0; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_7_1; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_7_2; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_7_3; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_7_4; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_7_5; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_7_6; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station2_7_7; // @[stationary_dpe.scala 26:25]
  reg [15:0] Station3_0_0; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_0_1; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_0_2; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_0_3; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_0_4; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_0_5; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_0_6; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_0_7; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_1_0; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_1_1; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_1_2; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_1_3; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_1_4; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_1_5; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_1_6; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_1_7; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_2_0; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_2_1; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_2_2; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_2_3; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_2_4; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_2_5; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_2_6; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_2_7; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_3_0; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_3_1; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_3_2; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_3_3; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_3_4; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_3_5; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_3_6; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_3_7; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_4_0; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_4_1; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_4_2; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_4_3; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_4_4; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_4_5; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_4_6; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_4_7; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_5_0; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_5_1; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_5_2; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_5_3; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_5_4; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_5_5; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_5_6; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_5_7; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_6_0; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_6_1; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_6_2; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_6_3; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_6_4; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_6_5; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_6_6; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_6_7; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_7_0; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_7_1; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_7_2; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_7_3; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_7_4; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_7_5; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_7_6; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station3_7_7; // @[stationary_dpe.scala 27:26]
  reg [15:0] Station4_0_0; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_0_1; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_0_2; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_0_3; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_0_4; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_0_5; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_0_6; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_0_7; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_1_0; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_1_1; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_1_2; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_1_3; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_1_4; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_1_5; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_1_6; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_1_7; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_2_0; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_2_1; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_2_2; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_2_3; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_2_4; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_2_5; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_2_6; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_2_7; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_3_0; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_3_1; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_3_2; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_3_3; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_3_4; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_3_5; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_3_6; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_3_7; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_4_0; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_4_1; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_4_2; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_4_3; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_4_4; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_4_5; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_4_6; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_4_7; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_5_0; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_5_1; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_5_2; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_5_3; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_5_4; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_5_5; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_5_6; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_5_7; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_6_0; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_6_1; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_6_2; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_6_3; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_6_4; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_6_5; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_6_6; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_6_7; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_7_0; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_7_1; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_7_2; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_7_3; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_7_4; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_7_5; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_7_6; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station4_7_7; // @[stationary_dpe.scala 28:27]
  reg [15:0] Station5_0_0; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_0_1; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_0_2; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_0_3; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_0_4; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_0_5; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_0_6; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_0_7; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_1_0; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_1_1; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_1_2; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_1_3; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_1_4; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_1_5; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_1_6; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_1_7; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_2_0; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_2_1; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_2_2; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_2_3; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_2_4; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_2_5; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_2_6; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_2_7; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_3_0; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_3_1; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_3_2; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_3_3; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_3_4; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_3_5; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_3_6; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_3_7; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_4_0; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_4_1; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_4_2; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_4_3; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_4_4; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_4_5; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_4_6; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_4_7; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_5_0; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_5_1; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_5_2; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_5_3; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_5_4; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_5_5; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_5_6; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_5_7; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_6_0; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_6_1; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_6_2; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_6_3; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_6_4; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_6_5; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_6_6; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_6_7; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_7_0; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_7_1; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_7_2; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_7_3; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_7_4; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_7_5; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_7_6; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station5_7_7; // @[stationary_dpe.scala 29:28]
  reg [15:0] Station6_0_0; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_0_1; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_0_2; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_0_3; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_0_4; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_0_5; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_0_6; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_0_7; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_1_0; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_1_1; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_1_2; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_1_3; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_1_4; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_1_5; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_1_6; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_1_7; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_2_0; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_2_1; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_2_2; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_2_3; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_2_4; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_2_5; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_2_6; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_2_7; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_3_0; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_3_1; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_3_2; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_3_3; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_3_4; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_3_5; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_3_6; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_3_7; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_4_0; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_4_1; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_4_2; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_4_3; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_4_4; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_4_5; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_4_6; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_4_7; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_5_0; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_5_1; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_5_2; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_5_3; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_5_4; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_5_5; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_5_6; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_5_7; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_6_0; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_6_1; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_6_2; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_6_3; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_6_4; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_6_5; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_6_6; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_6_7; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_7_0; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_7_1; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_7_2; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_7_3; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_7_4; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_7_5; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_7_6; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station6_7_7; // @[stationary_dpe.scala 30:29]
  reg [15:0] Station7_0_0; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_0_1; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_0_2; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_0_3; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_0_4; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_0_5; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_0_6; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_0_7; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_1_0; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_1_1; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_1_2; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_1_3; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_1_4; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_1_5; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_1_6; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_1_7; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_2_0; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_2_1; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_2_2; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_2_3; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_2_4; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_2_5; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_2_6; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_2_7; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_3_0; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_3_1; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_3_2; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_3_3; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_3_4; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_3_5; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_3_6; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_3_7; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_4_0; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_4_1; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_4_2; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_4_3; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_4_4; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_4_5; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_4_6; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_4_7; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_5_0; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_5_1; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_5_2; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_5_3; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_5_4; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_5_5; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_5_6; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_5_7; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_6_0; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_6_1; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_6_2; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_6_3; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_6_4; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_6_5; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_6_6; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_6_7; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_7_0; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_7_1; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_7_2; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_7_3; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_7_4; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_7_5; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_7_6; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station7_7_7; // @[stationary_dpe.scala 31:30]
  reg [15:0] Station8_0_0; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_0_1; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_0_2; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_0_3; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_0_4; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_0_5; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_0_6; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_0_7; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_1_0; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_1_1; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_1_2; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_1_3; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_1_4; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_1_5; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_1_6; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_1_7; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_2_0; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_2_1; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_2_2; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_2_3; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_2_4; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_2_5; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_2_6; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_2_7; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_3_0; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_3_1; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_3_2; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_3_3; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_3_4; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_3_5; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_3_6; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_3_7; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_4_0; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_4_1; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_4_2; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_4_3; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_4_4; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_4_5; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_4_6; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_4_7; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_5_0; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_5_1; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_5_2; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_5_3; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_5_4; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_5_5; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_5_6; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_5_7; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_6_0; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_6_1; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_6_2; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_6_3; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_6_4; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_6_5; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_6_6; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_6_7; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_7_0; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_7_1; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_7_2; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_7_3; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_7_4; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_7_5; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_7_6; // @[stationary_dpe.scala 32:31]
  reg [15:0] Station8_7_7; // @[stationary_dpe.scala 32:31]
  wire [15:0] _GEN_0 = count == 32'h0 ? io_Stationary_matrix_0_0 : Station2_0_0; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_1 = count == 32'h0 ? io_Stationary_matrix_0_1 : Station2_0_1; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_2 = count == 32'h0 ? io_Stationary_matrix_0_2 : Station2_0_2; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_3 = count == 32'h0 ? io_Stationary_matrix_0_3 : Station2_0_3; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_4 = count == 32'h0 ? io_Stationary_matrix_0_4 : Station2_0_4; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_5 = count == 32'h0 ? io_Stationary_matrix_0_5 : Station2_0_5; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_6 = count == 32'h0 ? io_Stationary_matrix_0_6 : Station2_0_6; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_7 = count == 32'h0 ? io_Stationary_matrix_0_7 : Station2_0_7; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_8 = count == 32'h0 ? io_Stationary_matrix_1_0 : Station2_1_0; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_9 = count == 32'h0 ? io_Stationary_matrix_1_1 : Station2_1_1; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_10 = count == 32'h0 ? io_Stationary_matrix_1_2 : Station2_1_2; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_11 = count == 32'h0 ? io_Stationary_matrix_1_3 : Station2_1_3; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_12 = count == 32'h0 ? io_Stationary_matrix_1_4 : Station2_1_4; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_13 = count == 32'h0 ? io_Stationary_matrix_1_5 : Station2_1_5; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_14 = count == 32'h0 ? io_Stationary_matrix_1_6 : Station2_1_6; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_15 = count == 32'h0 ? io_Stationary_matrix_1_7 : Station2_1_7; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_16 = count == 32'h0 ? io_Stationary_matrix_2_0 : Station2_2_0; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_17 = count == 32'h0 ? io_Stationary_matrix_2_1 : Station2_2_1; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_18 = count == 32'h0 ? io_Stationary_matrix_2_2 : Station2_2_2; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_19 = count == 32'h0 ? io_Stationary_matrix_2_3 : Station2_2_3; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_20 = count == 32'h0 ? io_Stationary_matrix_2_4 : Station2_2_4; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_21 = count == 32'h0 ? io_Stationary_matrix_2_5 : Station2_2_5; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_22 = count == 32'h0 ? io_Stationary_matrix_2_6 : Station2_2_6; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_23 = count == 32'h0 ? io_Stationary_matrix_2_7 : Station2_2_7; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_24 = count == 32'h0 ? io_Stationary_matrix_3_0 : Station2_3_0; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_25 = count == 32'h0 ? io_Stationary_matrix_3_1 : Station2_3_1; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_26 = count == 32'h0 ? io_Stationary_matrix_3_2 : Station2_3_2; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_27 = count == 32'h0 ? io_Stationary_matrix_3_3 : Station2_3_3; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_28 = count == 32'h0 ? io_Stationary_matrix_3_4 : Station2_3_4; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_29 = count == 32'h0 ? io_Stationary_matrix_3_5 : Station2_3_5; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_30 = count == 32'h0 ? io_Stationary_matrix_3_6 : Station2_3_6; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_31 = count == 32'h0 ? io_Stationary_matrix_3_7 : Station2_3_7; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_32 = count == 32'h0 ? io_Stationary_matrix_4_0 : Station2_4_0; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_33 = count == 32'h0 ? io_Stationary_matrix_4_1 : Station2_4_1; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_34 = count == 32'h0 ? io_Stationary_matrix_4_2 : Station2_4_2; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_35 = count == 32'h0 ? io_Stationary_matrix_4_3 : Station2_4_3; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_36 = count == 32'h0 ? io_Stationary_matrix_4_4 : Station2_4_4; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_37 = count == 32'h0 ? io_Stationary_matrix_4_5 : Station2_4_5; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_38 = count == 32'h0 ? io_Stationary_matrix_4_6 : Station2_4_6; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_39 = count == 32'h0 ? io_Stationary_matrix_4_7 : Station2_4_7; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_40 = count == 32'h0 ? io_Stationary_matrix_5_0 : Station2_5_0; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_41 = count == 32'h0 ? io_Stationary_matrix_5_1 : Station2_5_1; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_42 = count == 32'h0 ? io_Stationary_matrix_5_2 : Station2_5_2; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_43 = count == 32'h0 ? io_Stationary_matrix_5_3 : Station2_5_3; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_44 = count == 32'h0 ? io_Stationary_matrix_5_4 : Station2_5_4; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_45 = count == 32'h0 ? io_Stationary_matrix_5_5 : Station2_5_5; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_46 = count == 32'h0 ? io_Stationary_matrix_5_6 : Station2_5_6; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_47 = count == 32'h0 ? io_Stationary_matrix_5_7 : Station2_5_7; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_48 = count == 32'h0 ? io_Stationary_matrix_6_0 : Station2_6_0; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_49 = count == 32'h0 ? io_Stationary_matrix_6_1 : Station2_6_1; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_50 = count == 32'h0 ? io_Stationary_matrix_6_2 : Station2_6_2; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_51 = count == 32'h0 ? io_Stationary_matrix_6_3 : Station2_6_3; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_52 = count == 32'h0 ? io_Stationary_matrix_6_4 : Station2_6_4; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_53 = count == 32'h0 ? io_Stationary_matrix_6_5 : Station2_6_5; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_54 = count == 32'h0 ? io_Stationary_matrix_6_6 : Station2_6_6; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_55 = count == 32'h0 ? io_Stationary_matrix_6_7 : Station2_6_7; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_56 = count == 32'h0 ? io_Stationary_matrix_7_0 : Station2_7_0; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_57 = count == 32'h0 ? io_Stationary_matrix_7_1 : Station2_7_1; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_58 = count == 32'h0 ? io_Stationary_matrix_7_2 : Station2_7_2; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_59 = count == 32'h0 ? io_Stationary_matrix_7_3 : Station2_7_3; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_60 = count == 32'h0 ? io_Stationary_matrix_7_4 : Station2_7_4; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_61 = count == 32'h0 ? io_Stationary_matrix_7_5 : Station2_7_5; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_62 = count == 32'h0 ? io_Stationary_matrix_7_6 : Station2_7_6; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_63 = count == 32'h0 ? io_Stationary_matrix_7_7 : Station2_7_7; // @[stationary_dpe.scala 45:24 46:15 26:25]
  wire [15:0] _GEN_64 = count == 32'h8 ? Station2_0_0 : Station3_0_0; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_65 = count == 32'h8 ? Station2_0_1 : Station3_0_1; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_66 = count == 32'h8 ? Station2_0_2 : Station3_0_2; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_67 = count == 32'h8 ? Station2_0_3 : Station3_0_3; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_68 = count == 32'h8 ? Station2_0_4 : Station3_0_4; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_69 = count == 32'h8 ? Station2_0_5 : Station3_0_5; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_70 = count == 32'h8 ? Station2_0_6 : Station3_0_6; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_71 = count == 32'h8 ? Station2_0_7 : Station3_0_7; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_72 = count == 32'h8 ? Station2_1_0 : Station3_1_0; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_73 = count == 32'h8 ? Station2_1_1 : Station3_1_1; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_74 = count == 32'h8 ? Station2_1_2 : Station3_1_2; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_75 = count == 32'h8 ? Station2_1_3 : Station3_1_3; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_76 = count == 32'h8 ? Station2_1_4 : Station3_1_4; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_77 = count == 32'h8 ? Station2_1_5 : Station3_1_5; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_78 = count == 32'h8 ? Station2_1_6 : Station3_1_6; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_79 = count == 32'h8 ? Station2_1_7 : Station3_1_7; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_80 = count == 32'h8 ? Station2_2_0 : Station3_2_0; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_81 = count == 32'h8 ? Station2_2_1 : Station3_2_1; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_82 = count == 32'h8 ? Station2_2_2 : Station3_2_2; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_83 = count == 32'h8 ? Station2_2_3 : Station3_2_3; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_84 = count == 32'h8 ? Station2_2_4 : Station3_2_4; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_85 = count == 32'h8 ? Station2_2_5 : Station3_2_5; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_86 = count == 32'h8 ? Station2_2_6 : Station3_2_6; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_87 = count == 32'h8 ? Station2_2_7 : Station3_2_7; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_88 = count == 32'h8 ? Station2_3_0 : Station3_3_0; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_89 = count == 32'h8 ? Station2_3_1 : Station3_3_1; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_90 = count == 32'h8 ? Station2_3_2 : Station3_3_2; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_91 = count == 32'h8 ? Station2_3_3 : Station3_3_3; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_92 = count == 32'h8 ? Station2_3_4 : Station3_3_4; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_93 = count == 32'h8 ? Station2_3_5 : Station3_3_5; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_94 = count == 32'h8 ? Station2_3_6 : Station3_3_6; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_95 = count == 32'h8 ? Station2_3_7 : Station3_3_7; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_96 = count == 32'h8 ? Station2_4_0 : Station3_4_0; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_97 = count == 32'h8 ? Station2_4_1 : Station3_4_1; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_98 = count == 32'h8 ? Station2_4_2 : Station3_4_2; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_99 = count == 32'h8 ? Station2_4_3 : Station3_4_3; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_100 = count == 32'h8 ? Station2_4_4 : Station3_4_4; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_101 = count == 32'h8 ? Station2_4_5 : Station3_4_5; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_102 = count == 32'h8 ? Station2_4_6 : Station3_4_6; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_103 = count == 32'h8 ? Station2_4_7 : Station3_4_7; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_104 = count == 32'h8 ? Station2_5_0 : Station3_5_0; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_105 = count == 32'h8 ? Station2_5_1 : Station3_5_1; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_106 = count == 32'h8 ? Station2_5_2 : Station3_5_2; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_107 = count == 32'h8 ? Station2_5_3 : Station3_5_3; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_108 = count == 32'h8 ? Station2_5_4 : Station3_5_4; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_109 = count == 32'h8 ? Station2_5_5 : Station3_5_5; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_110 = count == 32'h8 ? Station2_5_6 : Station3_5_6; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_111 = count == 32'h8 ? Station2_5_7 : Station3_5_7; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_112 = count == 32'h8 ? Station2_6_0 : Station3_6_0; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_113 = count == 32'h8 ? Station2_6_1 : Station3_6_1; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_114 = count == 32'h8 ? Station2_6_2 : Station3_6_2; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_115 = count == 32'h8 ? Station2_6_3 : Station3_6_3; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_116 = count == 32'h8 ? Station2_6_4 : Station3_6_4; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_117 = count == 32'h8 ? Station2_6_5 : Station3_6_5; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_118 = count == 32'h8 ? Station2_6_6 : Station3_6_6; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_119 = count == 32'h8 ? Station2_6_7 : Station3_6_7; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_120 = count == 32'h8 ? Station2_7_0 : Station3_7_0; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_121 = count == 32'h8 ? Station2_7_1 : Station3_7_1; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_122 = count == 32'h8 ? Station2_7_2 : Station3_7_2; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_123 = count == 32'h8 ? Station2_7_3 : Station3_7_3; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_124 = count == 32'h8 ? Station2_7_4 : Station3_7_4; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_125 = count == 32'h8 ? Station2_7_5 : Station3_7_5; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_126 = count == 32'h8 ? Station2_7_6 : Station3_7_6; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_127 = count == 32'h8 ? Station2_7_7 : Station3_7_7; // @[stationary_dpe.scala 49:24 50:15 27:26]
  wire [15:0] _GEN_128 = count == 32'h10 ? Station3_0_0 : Station4_0_0; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_129 = count == 32'h10 ? Station3_0_1 : Station4_0_1; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_130 = count == 32'h10 ? Station3_0_2 : Station4_0_2; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_131 = count == 32'h10 ? Station3_0_3 : Station4_0_3; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_132 = count == 32'h10 ? Station3_0_4 : Station4_0_4; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_133 = count == 32'h10 ? Station3_0_5 : Station4_0_5; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_134 = count == 32'h10 ? Station3_0_6 : Station4_0_6; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_135 = count == 32'h10 ? Station3_0_7 : Station4_0_7; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_136 = count == 32'h10 ? Station3_1_0 : Station4_1_0; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_137 = count == 32'h10 ? Station3_1_1 : Station4_1_1; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_138 = count == 32'h10 ? Station3_1_2 : Station4_1_2; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_139 = count == 32'h10 ? Station3_1_3 : Station4_1_3; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_140 = count == 32'h10 ? Station3_1_4 : Station4_1_4; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_141 = count == 32'h10 ? Station3_1_5 : Station4_1_5; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_142 = count == 32'h10 ? Station3_1_6 : Station4_1_6; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_143 = count == 32'h10 ? Station3_1_7 : Station4_1_7; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_144 = count == 32'h10 ? Station3_2_0 : Station4_2_0; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_145 = count == 32'h10 ? Station3_2_1 : Station4_2_1; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_146 = count == 32'h10 ? Station3_2_2 : Station4_2_2; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_147 = count == 32'h10 ? Station3_2_3 : Station4_2_3; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_148 = count == 32'h10 ? Station3_2_4 : Station4_2_4; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_149 = count == 32'h10 ? Station3_2_5 : Station4_2_5; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_150 = count == 32'h10 ? Station3_2_6 : Station4_2_6; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_151 = count == 32'h10 ? Station3_2_7 : Station4_2_7; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_152 = count == 32'h10 ? Station3_3_0 : Station4_3_0; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_153 = count == 32'h10 ? Station3_3_1 : Station4_3_1; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_154 = count == 32'h10 ? Station3_3_2 : Station4_3_2; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_155 = count == 32'h10 ? Station3_3_3 : Station4_3_3; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_156 = count == 32'h10 ? Station3_3_4 : Station4_3_4; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_157 = count == 32'h10 ? Station3_3_5 : Station4_3_5; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_158 = count == 32'h10 ? Station3_3_6 : Station4_3_6; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_159 = count == 32'h10 ? Station3_3_7 : Station4_3_7; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_160 = count == 32'h10 ? Station3_4_0 : Station4_4_0; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_161 = count == 32'h10 ? Station3_4_1 : Station4_4_1; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_162 = count == 32'h10 ? Station3_4_2 : Station4_4_2; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_163 = count == 32'h10 ? Station3_4_3 : Station4_4_3; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_164 = count == 32'h10 ? Station3_4_4 : Station4_4_4; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_165 = count == 32'h10 ? Station3_4_5 : Station4_4_5; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_166 = count == 32'h10 ? Station3_4_6 : Station4_4_6; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_167 = count == 32'h10 ? Station3_4_7 : Station4_4_7; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_168 = count == 32'h10 ? Station3_5_0 : Station4_5_0; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_169 = count == 32'h10 ? Station3_5_1 : Station4_5_1; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_170 = count == 32'h10 ? Station3_5_2 : Station4_5_2; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_171 = count == 32'h10 ? Station3_5_3 : Station4_5_3; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_172 = count == 32'h10 ? Station3_5_4 : Station4_5_4; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_173 = count == 32'h10 ? Station3_5_5 : Station4_5_5; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_174 = count == 32'h10 ? Station3_5_6 : Station4_5_6; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_175 = count == 32'h10 ? Station3_5_7 : Station4_5_7; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_176 = count == 32'h10 ? Station3_6_0 : Station4_6_0; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_177 = count == 32'h10 ? Station3_6_1 : Station4_6_1; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_178 = count == 32'h10 ? Station3_6_2 : Station4_6_2; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_179 = count == 32'h10 ? Station3_6_3 : Station4_6_3; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_180 = count == 32'h10 ? Station3_6_4 : Station4_6_4; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_181 = count == 32'h10 ? Station3_6_5 : Station4_6_5; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_182 = count == 32'h10 ? Station3_6_6 : Station4_6_6; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_183 = count == 32'h10 ? Station3_6_7 : Station4_6_7; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_184 = count == 32'h10 ? Station3_7_0 : Station4_7_0; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_185 = count == 32'h10 ? Station3_7_1 : Station4_7_1; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_186 = count == 32'h10 ? Station3_7_2 : Station4_7_2; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_187 = count == 32'h10 ? Station3_7_3 : Station4_7_3; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_188 = count == 32'h10 ? Station3_7_4 : Station4_7_4; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_189 = count == 32'h10 ? Station3_7_5 : Station4_7_5; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_190 = count == 32'h10 ? Station3_7_6 : Station4_7_6; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_191 = count == 32'h10 ? Station3_7_7 : Station4_7_7; // @[stationary_dpe.scala 54:27 55:15 28:27]
  wire [15:0] _GEN_192 = count == 32'h18 ? Station4_0_0 : Station5_0_0; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_193 = count == 32'h18 ? Station4_0_1 : Station5_0_1; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_194 = count == 32'h18 ? Station4_0_2 : Station5_0_2; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_195 = count == 32'h18 ? Station4_0_3 : Station5_0_3; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_196 = count == 32'h18 ? Station4_0_4 : Station5_0_4; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_197 = count == 32'h18 ? Station4_0_5 : Station5_0_5; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_198 = count == 32'h18 ? Station4_0_6 : Station5_0_6; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_199 = count == 32'h18 ? Station4_0_7 : Station5_0_7; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_200 = count == 32'h18 ? Station4_1_0 : Station5_1_0; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_201 = count == 32'h18 ? Station4_1_1 : Station5_1_1; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_202 = count == 32'h18 ? Station4_1_2 : Station5_1_2; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_203 = count == 32'h18 ? Station4_1_3 : Station5_1_3; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_204 = count == 32'h18 ? Station4_1_4 : Station5_1_4; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_205 = count == 32'h18 ? Station4_1_5 : Station5_1_5; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_206 = count == 32'h18 ? Station4_1_6 : Station5_1_6; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_207 = count == 32'h18 ? Station4_1_7 : Station5_1_7; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_208 = count == 32'h18 ? Station4_2_0 : Station5_2_0; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_209 = count == 32'h18 ? Station4_2_1 : Station5_2_1; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_210 = count == 32'h18 ? Station4_2_2 : Station5_2_2; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_211 = count == 32'h18 ? Station4_2_3 : Station5_2_3; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_212 = count == 32'h18 ? Station4_2_4 : Station5_2_4; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_213 = count == 32'h18 ? Station4_2_5 : Station5_2_5; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_214 = count == 32'h18 ? Station4_2_6 : Station5_2_6; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_215 = count == 32'h18 ? Station4_2_7 : Station5_2_7; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_216 = count == 32'h18 ? Station4_3_0 : Station5_3_0; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_217 = count == 32'h18 ? Station4_3_1 : Station5_3_1; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_218 = count == 32'h18 ? Station4_3_2 : Station5_3_2; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_219 = count == 32'h18 ? Station4_3_3 : Station5_3_3; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_220 = count == 32'h18 ? Station4_3_4 : Station5_3_4; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_221 = count == 32'h18 ? Station4_3_5 : Station5_3_5; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_222 = count == 32'h18 ? Station4_3_6 : Station5_3_6; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_223 = count == 32'h18 ? Station4_3_7 : Station5_3_7; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_224 = count == 32'h18 ? Station4_4_0 : Station5_4_0; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_225 = count == 32'h18 ? Station4_4_1 : Station5_4_1; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_226 = count == 32'h18 ? Station4_4_2 : Station5_4_2; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_227 = count == 32'h18 ? Station4_4_3 : Station5_4_3; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_228 = count == 32'h18 ? Station4_4_4 : Station5_4_4; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_229 = count == 32'h18 ? Station4_4_5 : Station5_4_5; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_230 = count == 32'h18 ? Station4_4_6 : Station5_4_6; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_231 = count == 32'h18 ? Station4_4_7 : Station5_4_7; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_232 = count == 32'h18 ? Station4_5_0 : Station5_5_0; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_233 = count == 32'h18 ? Station4_5_1 : Station5_5_1; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_234 = count == 32'h18 ? Station4_5_2 : Station5_5_2; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_235 = count == 32'h18 ? Station4_5_3 : Station5_5_3; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_236 = count == 32'h18 ? Station4_5_4 : Station5_5_4; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_237 = count == 32'h18 ? Station4_5_5 : Station5_5_5; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_238 = count == 32'h18 ? Station4_5_6 : Station5_5_6; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_239 = count == 32'h18 ? Station4_5_7 : Station5_5_7; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_240 = count == 32'h18 ? Station4_6_0 : Station5_6_0; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_241 = count == 32'h18 ? Station4_6_1 : Station5_6_1; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_242 = count == 32'h18 ? Station4_6_2 : Station5_6_2; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_243 = count == 32'h18 ? Station4_6_3 : Station5_6_3; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_244 = count == 32'h18 ? Station4_6_4 : Station5_6_4; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_245 = count == 32'h18 ? Station4_6_5 : Station5_6_5; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_246 = count == 32'h18 ? Station4_6_6 : Station5_6_6; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_247 = count == 32'h18 ? Station4_6_7 : Station5_6_7; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_248 = count == 32'h18 ? Station4_7_0 : Station5_7_0; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_249 = count == 32'h18 ? Station4_7_1 : Station5_7_1; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_250 = count == 32'h18 ? Station4_7_2 : Station5_7_2; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_251 = count == 32'h18 ? Station4_7_3 : Station5_7_3; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_252 = count == 32'h18 ? Station4_7_4 : Station5_7_4; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_253 = count == 32'h18 ? Station4_7_5 : Station5_7_5; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_254 = count == 32'h18 ? Station4_7_6 : Station5_7_6; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_255 = count == 32'h18 ? Station4_7_7 : Station5_7_7; // @[stationary_dpe.scala 58:27 59:15 29:28]
  wire [15:0] _GEN_256 = count == 32'h20 ? Station5_0_0 : Station6_0_0; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_257 = count == 32'h20 ? Station5_0_1 : Station6_0_1; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_258 = count == 32'h20 ? Station5_0_2 : Station6_0_2; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_259 = count == 32'h20 ? Station5_0_3 : Station6_0_3; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_260 = count == 32'h20 ? Station5_0_4 : Station6_0_4; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_261 = count == 32'h20 ? Station5_0_5 : Station6_0_5; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_262 = count == 32'h20 ? Station5_0_6 : Station6_0_6; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_263 = count == 32'h20 ? Station5_0_7 : Station6_0_7; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_264 = count == 32'h20 ? Station5_1_0 : Station6_1_0; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_265 = count == 32'h20 ? Station5_1_1 : Station6_1_1; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_266 = count == 32'h20 ? Station5_1_2 : Station6_1_2; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_267 = count == 32'h20 ? Station5_1_3 : Station6_1_3; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_268 = count == 32'h20 ? Station5_1_4 : Station6_1_4; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_269 = count == 32'h20 ? Station5_1_5 : Station6_1_5; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_270 = count == 32'h20 ? Station5_1_6 : Station6_1_6; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_271 = count == 32'h20 ? Station5_1_7 : Station6_1_7; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_272 = count == 32'h20 ? Station5_2_0 : Station6_2_0; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_273 = count == 32'h20 ? Station5_2_1 : Station6_2_1; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_274 = count == 32'h20 ? Station5_2_2 : Station6_2_2; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_275 = count == 32'h20 ? Station5_2_3 : Station6_2_3; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_276 = count == 32'h20 ? Station5_2_4 : Station6_2_4; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_277 = count == 32'h20 ? Station5_2_5 : Station6_2_5; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_278 = count == 32'h20 ? Station5_2_6 : Station6_2_6; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_279 = count == 32'h20 ? Station5_2_7 : Station6_2_7; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_280 = count == 32'h20 ? Station5_3_0 : Station6_3_0; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_281 = count == 32'h20 ? Station5_3_1 : Station6_3_1; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_282 = count == 32'h20 ? Station5_3_2 : Station6_3_2; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_283 = count == 32'h20 ? Station5_3_3 : Station6_3_3; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_284 = count == 32'h20 ? Station5_3_4 : Station6_3_4; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_285 = count == 32'h20 ? Station5_3_5 : Station6_3_5; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_286 = count == 32'h20 ? Station5_3_6 : Station6_3_6; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_287 = count == 32'h20 ? Station5_3_7 : Station6_3_7; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_288 = count == 32'h20 ? Station5_4_0 : Station6_4_0; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_289 = count == 32'h20 ? Station5_4_1 : Station6_4_1; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_290 = count == 32'h20 ? Station5_4_2 : Station6_4_2; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_291 = count == 32'h20 ? Station5_4_3 : Station6_4_3; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_292 = count == 32'h20 ? Station5_4_4 : Station6_4_4; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_293 = count == 32'h20 ? Station5_4_5 : Station6_4_5; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_294 = count == 32'h20 ? Station5_4_6 : Station6_4_6; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_295 = count == 32'h20 ? Station5_4_7 : Station6_4_7; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_296 = count == 32'h20 ? Station5_5_0 : Station6_5_0; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_297 = count == 32'h20 ? Station5_5_1 : Station6_5_1; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_298 = count == 32'h20 ? Station5_5_2 : Station6_5_2; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_299 = count == 32'h20 ? Station5_5_3 : Station6_5_3; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_300 = count == 32'h20 ? Station5_5_4 : Station6_5_4; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_301 = count == 32'h20 ? Station5_5_5 : Station6_5_5; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_302 = count == 32'h20 ? Station5_5_6 : Station6_5_6; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_303 = count == 32'h20 ? Station5_5_7 : Station6_5_7; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_304 = count == 32'h20 ? Station5_6_0 : Station6_6_0; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_305 = count == 32'h20 ? Station5_6_1 : Station6_6_1; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_306 = count == 32'h20 ? Station5_6_2 : Station6_6_2; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_307 = count == 32'h20 ? Station5_6_3 : Station6_6_3; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_308 = count == 32'h20 ? Station5_6_4 : Station6_6_4; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_309 = count == 32'h20 ? Station5_6_5 : Station6_6_5; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_310 = count == 32'h20 ? Station5_6_6 : Station6_6_6; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_311 = count == 32'h20 ? Station5_6_7 : Station6_6_7; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_312 = count == 32'h20 ? Station5_7_0 : Station6_7_0; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_313 = count == 32'h20 ? Station5_7_1 : Station6_7_1; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_314 = count == 32'h20 ? Station5_7_2 : Station6_7_2; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_315 = count == 32'h20 ? Station5_7_3 : Station6_7_3; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_316 = count == 32'h20 ? Station5_7_4 : Station6_7_4; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_317 = count == 32'h20 ? Station5_7_5 : Station6_7_5; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_318 = count == 32'h20 ? Station5_7_6 : Station6_7_6; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_319 = count == 32'h20 ? Station5_7_7 : Station6_7_7; // @[stationary_dpe.scala 62:27 63:15 30:29]
  wire [15:0] _GEN_320 = count == 32'h28 ? Station6_0_0 : Station7_0_0; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_321 = count == 32'h28 ? Station6_0_1 : Station7_0_1; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_322 = count == 32'h28 ? Station6_0_2 : Station7_0_2; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_323 = count == 32'h28 ? Station6_0_3 : Station7_0_3; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_324 = count == 32'h28 ? Station6_0_4 : Station7_0_4; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_325 = count == 32'h28 ? Station6_0_5 : Station7_0_5; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_326 = count == 32'h28 ? Station6_0_6 : Station7_0_6; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_327 = count == 32'h28 ? Station6_0_7 : Station7_0_7; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_328 = count == 32'h28 ? Station6_1_0 : Station7_1_0; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_329 = count == 32'h28 ? Station6_1_1 : Station7_1_1; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_330 = count == 32'h28 ? Station6_1_2 : Station7_1_2; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_331 = count == 32'h28 ? Station6_1_3 : Station7_1_3; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_332 = count == 32'h28 ? Station6_1_4 : Station7_1_4; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_333 = count == 32'h28 ? Station6_1_5 : Station7_1_5; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_334 = count == 32'h28 ? Station6_1_6 : Station7_1_6; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_335 = count == 32'h28 ? Station6_1_7 : Station7_1_7; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_336 = count == 32'h28 ? Station6_2_0 : Station7_2_0; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_337 = count == 32'h28 ? Station6_2_1 : Station7_2_1; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_338 = count == 32'h28 ? Station6_2_2 : Station7_2_2; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_339 = count == 32'h28 ? Station6_2_3 : Station7_2_3; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_340 = count == 32'h28 ? Station6_2_4 : Station7_2_4; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_341 = count == 32'h28 ? Station6_2_5 : Station7_2_5; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_342 = count == 32'h28 ? Station6_2_6 : Station7_2_6; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_343 = count == 32'h28 ? Station6_2_7 : Station7_2_7; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_344 = count == 32'h28 ? Station6_3_0 : Station7_3_0; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_345 = count == 32'h28 ? Station6_3_1 : Station7_3_1; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_346 = count == 32'h28 ? Station6_3_2 : Station7_3_2; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_347 = count == 32'h28 ? Station6_3_3 : Station7_3_3; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_348 = count == 32'h28 ? Station6_3_4 : Station7_3_4; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_349 = count == 32'h28 ? Station6_3_5 : Station7_3_5; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_350 = count == 32'h28 ? Station6_3_6 : Station7_3_6; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_351 = count == 32'h28 ? Station6_3_7 : Station7_3_7; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_352 = count == 32'h28 ? Station6_4_0 : Station7_4_0; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_353 = count == 32'h28 ? Station6_4_1 : Station7_4_1; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_354 = count == 32'h28 ? Station6_4_2 : Station7_4_2; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_355 = count == 32'h28 ? Station6_4_3 : Station7_4_3; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_356 = count == 32'h28 ? Station6_4_4 : Station7_4_4; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_357 = count == 32'h28 ? Station6_4_5 : Station7_4_5; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_358 = count == 32'h28 ? Station6_4_6 : Station7_4_6; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_359 = count == 32'h28 ? Station6_4_7 : Station7_4_7; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_360 = count == 32'h28 ? Station6_5_0 : Station7_5_0; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_361 = count == 32'h28 ? Station6_5_1 : Station7_5_1; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_362 = count == 32'h28 ? Station6_5_2 : Station7_5_2; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_363 = count == 32'h28 ? Station6_5_3 : Station7_5_3; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_364 = count == 32'h28 ? Station6_5_4 : Station7_5_4; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_365 = count == 32'h28 ? Station6_5_5 : Station7_5_5; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_366 = count == 32'h28 ? Station6_5_6 : Station7_5_6; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_367 = count == 32'h28 ? Station6_5_7 : Station7_5_7; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_368 = count == 32'h28 ? Station6_6_0 : Station7_6_0; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_369 = count == 32'h28 ? Station6_6_1 : Station7_6_1; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_370 = count == 32'h28 ? Station6_6_2 : Station7_6_2; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_371 = count == 32'h28 ? Station6_6_3 : Station7_6_3; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_372 = count == 32'h28 ? Station6_6_4 : Station7_6_4; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_373 = count == 32'h28 ? Station6_6_5 : Station7_6_5; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_374 = count == 32'h28 ? Station6_6_6 : Station7_6_6; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_375 = count == 32'h28 ? Station6_6_7 : Station7_6_7; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_376 = count == 32'h28 ? Station6_7_0 : Station7_7_0; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_377 = count == 32'h28 ? Station6_7_1 : Station7_7_1; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_378 = count == 32'h28 ? Station6_7_2 : Station7_7_2; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_379 = count == 32'h28 ? Station6_7_3 : Station7_7_3; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_380 = count == 32'h28 ? Station6_7_4 : Station7_7_4; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_381 = count == 32'h28 ? Station6_7_5 : Station7_7_5; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_382 = count == 32'h28 ? Station6_7_6 : Station7_7_6; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_383 = count == 32'h28 ? Station6_7_7 : Station7_7_7; // @[stationary_dpe.scala 66:27 67:15 31:30]
  wire [15:0] _GEN_384 = count == 32'h30 ? Station7_0_0 : Station8_0_0; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_385 = count == 32'h30 ? Station7_0_1 : Station8_0_1; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_386 = count == 32'h30 ? Station7_0_2 : Station8_0_2; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_387 = count == 32'h30 ? Station7_0_3 : Station8_0_3; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_388 = count == 32'h30 ? Station7_0_4 : Station8_0_4; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_389 = count == 32'h30 ? Station7_0_5 : Station8_0_5; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_390 = count == 32'h30 ? Station7_0_6 : Station8_0_6; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_391 = count == 32'h30 ? Station7_0_7 : Station8_0_7; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_392 = count == 32'h30 ? Station7_1_0 : Station8_1_0; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_393 = count == 32'h30 ? Station7_1_1 : Station8_1_1; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_394 = count == 32'h30 ? Station7_1_2 : Station8_1_2; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_395 = count == 32'h30 ? Station7_1_3 : Station8_1_3; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_396 = count == 32'h30 ? Station7_1_4 : Station8_1_4; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_397 = count == 32'h30 ? Station7_1_5 : Station8_1_5; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_398 = count == 32'h30 ? Station7_1_6 : Station8_1_6; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_399 = count == 32'h30 ? Station7_1_7 : Station8_1_7; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_400 = count == 32'h30 ? Station7_2_0 : Station8_2_0; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_401 = count == 32'h30 ? Station7_2_1 : Station8_2_1; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_402 = count == 32'h30 ? Station7_2_2 : Station8_2_2; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_403 = count == 32'h30 ? Station7_2_3 : Station8_2_3; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_404 = count == 32'h30 ? Station7_2_4 : Station8_2_4; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_405 = count == 32'h30 ? Station7_2_5 : Station8_2_5; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_406 = count == 32'h30 ? Station7_2_6 : Station8_2_6; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_407 = count == 32'h30 ? Station7_2_7 : Station8_2_7; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_408 = count == 32'h30 ? Station7_3_0 : Station8_3_0; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_409 = count == 32'h30 ? Station7_3_1 : Station8_3_1; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_410 = count == 32'h30 ? Station7_3_2 : Station8_3_2; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_411 = count == 32'h30 ? Station7_3_3 : Station8_3_3; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_412 = count == 32'h30 ? Station7_3_4 : Station8_3_4; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_413 = count == 32'h30 ? Station7_3_5 : Station8_3_5; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_414 = count == 32'h30 ? Station7_3_6 : Station8_3_6; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_415 = count == 32'h30 ? Station7_3_7 : Station8_3_7; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_416 = count == 32'h30 ? Station7_4_0 : Station8_4_0; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_417 = count == 32'h30 ? Station7_4_1 : Station8_4_1; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_418 = count == 32'h30 ? Station7_4_2 : Station8_4_2; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_419 = count == 32'h30 ? Station7_4_3 : Station8_4_3; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_420 = count == 32'h30 ? Station7_4_4 : Station8_4_4; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_421 = count == 32'h30 ? Station7_4_5 : Station8_4_5; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_422 = count == 32'h30 ? Station7_4_6 : Station8_4_6; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_423 = count == 32'h30 ? Station7_4_7 : Station8_4_7; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_424 = count == 32'h30 ? Station7_5_0 : Station8_5_0; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_425 = count == 32'h30 ? Station7_5_1 : Station8_5_1; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_426 = count == 32'h30 ? Station7_5_2 : Station8_5_2; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_427 = count == 32'h30 ? Station7_5_3 : Station8_5_3; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_428 = count == 32'h30 ? Station7_5_4 : Station8_5_4; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_429 = count == 32'h30 ? Station7_5_5 : Station8_5_5; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_430 = count == 32'h30 ? Station7_5_6 : Station8_5_6; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_431 = count == 32'h30 ? Station7_5_7 : Station8_5_7; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_432 = count == 32'h30 ? Station7_6_0 : Station8_6_0; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_433 = count == 32'h30 ? Station7_6_1 : Station8_6_1; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_434 = count == 32'h30 ? Station7_6_2 : Station8_6_2; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_435 = count == 32'h30 ? Station7_6_3 : Station8_6_3; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_436 = count == 32'h30 ? Station7_6_4 : Station8_6_4; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_437 = count == 32'h30 ? Station7_6_5 : Station8_6_5; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_438 = count == 32'h30 ? Station7_6_6 : Station8_6_6; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_439 = count == 32'h30 ? Station7_6_7 : Station8_6_7; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_440 = count == 32'h30 ? Station7_7_0 : Station8_7_0; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_441 = count == 32'h30 ? Station7_7_1 : Station8_7_1; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_442 = count == 32'h30 ? Station7_7_2 : Station8_7_2; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_443 = count == 32'h30 ? Station7_7_3 : Station8_7_3; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_444 = count == 32'h30 ? Station7_7_4 : Station8_7_4; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_445 = count == 32'h30 ? Station7_7_5 : Station8_7_5; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_446 = count == 32'h30 ? Station7_7_6 : Station8_7_6; // @[stationary_dpe.scala 70:27 71:15 32:31]
  wire [15:0] _GEN_447 = count == 32'h30 ? Station7_7_7 : Station8_7_7; // @[stationary_dpe.scala 70:27 71:15 32:31]
  reg [31:0] i; // @[stationary_dpe.scala 79:20]
  reg [31:0] j; // @[stationary_dpe.scala 80:20]
  wire  valid = count >= 32'h8; // @[stationary_dpe.scala 190:17]
  wire  _GEN_2264 = 3'h0 == i[2:0]; // @[stationary_dpe.scala 94:{43,43}]
  wire  _GEN_2265 = 3'h1 == j[2:0]; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_449 = 3'h0 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_0_1 : io_Stationary_matrix_0_0; // @[stationary_dpe.scala 94:{43,43}]
  wire  _GEN_2267 = 3'h2 == j[2:0]; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_450 = 3'h0 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_0_2 : _GEN_449; // @[stationary_dpe.scala 94:{43,43}]
  wire  _GEN_2269 = 3'h3 == j[2:0]; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_451 = 3'h0 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_0_3 : _GEN_450; // @[stationary_dpe.scala 94:{43,43}]
  wire  _GEN_2271 = 3'h4 == j[2:0]; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_452 = 3'h0 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_0_4 : _GEN_451; // @[stationary_dpe.scala 94:{43,43}]
  wire  _GEN_2273 = 3'h5 == j[2:0]; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_453 = 3'h0 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_0_5 : _GEN_452; // @[stationary_dpe.scala 94:{43,43}]
  wire  _GEN_2275 = 3'h6 == j[2:0]; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_454 = 3'h0 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_0_6 : _GEN_453; // @[stationary_dpe.scala 94:{43,43}]
  wire  _GEN_2277 = 3'h7 == j[2:0]; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_455 = 3'h0 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_0_7 : _GEN_454; // @[stationary_dpe.scala 94:{43,43}]
  wire  _GEN_2278 = 3'h1 == i[2:0]; // @[stationary_dpe.scala 94:{43,43}]
  wire  _GEN_2279 = 3'h0 == j[2:0]; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_456 = 3'h1 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_1_0 : _GEN_455; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_457 = 3'h1 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_1_1 : _GEN_456; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_458 = 3'h1 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_1_2 : _GEN_457; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_459 = 3'h1 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_1_3 : _GEN_458; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_460 = 3'h1 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_1_4 : _GEN_459; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_461 = 3'h1 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_1_5 : _GEN_460; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_462 = 3'h1 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_1_6 : _GEN_461; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_463 = 3'h1 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_1_7 : _GEN_462; // @[stationary_dpe.scala 94:{43,43}]
  wire  _GEN_2294 = 3'h2 == i[2:0]; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_464 = 3'h2 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_2_0 : _GEN_463; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_465 = 3'h2 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_2_1 : _GEN_464; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_466 = 3'h2 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_2_2 : _GEN_465; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_467 = 3'h2 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_2_3 : _GEN_466; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_468 = 3'h2 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_2_4 : _GEN_467; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_469 = 3'h2 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_2_5 : _GEN_468; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_470 = 3'h2 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_2_6 : _GEN_469; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_471 = 3'h2 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_2_7 : _GEN_470; // @[stationary_dpe.scala 94:{43,43}]
  wire  _GEN_2310 = 3'h3 == i[2:0]; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_472 = 3'h3 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_3_0 : _GEN_471; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_473 = 3'h3 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_3_1 : _GEN_472; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_474 = 3'h3 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_3_2 : _GEN_473; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_475 = 3'h3 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_3_3 : _GEN_474; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_476 = 3'h3 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_3_4 : _GEN_475; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_477 = 3'h3 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_3_5 : _GEN_476; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_478 = 3'h3 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_3_6 : _GEN_477; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_479 = 3'h3 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_3_7 : _GEN_478; // @[stationary_dpe.scala 94:{43,43}]
  wire  _GEN_2326 = 3'h4 == i[2:0]; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_480 = 3'h4 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_4_0 : _GEN_479; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_481 = 3'h4 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_4_1 : _GEN_480; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_482 = 3'h4 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_4_2 : _GEN_481; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_483 = 3'h4 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_4_3 : _GEN_482; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_484 = 3'h4 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_4_4 : _GEN_483; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_485 = 3'h4 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_4_5 : _GEN_484; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_486 = 3'h4 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_4_6 : _GEN_485; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_487 = 3'h4 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_4_7 : _GEN_486; // @[stationary_dpe.scala 94:{43,43}]
  wire  _GEN_2342 = 3'h5 == i[2:0]; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_488 = 3'h5 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_5_0 : _GEN_487; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_489 = 3'h5 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_5_1 : _GEN_488; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_490 = 3'h5 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_5_2 : _GEN_489; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_491 = 3'h5 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_5_3 : _GEN_490; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_492 = 3'h5 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_5_4 : _GEN_491; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_493 = 3'h5 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_5_5 : _GEN_492; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_494 = 3'h5 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_5_6 : _GEN_493; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_495 = 3'h5 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_5_7 : _GEN_494; // @[stationary_dpe.scala 94:{43,43}]
  wire  _GEN_2358 = 3'h6 == i[2:0]; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_496 = 3'h6 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_6_0 : _GEN_495; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_497 = 3'h6 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_6_1 : _GEN_496; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_498 = 3'h6 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_6_2 : _GEN_497; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_499 = 3'h6 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_6_3 : _GEN_498; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_500 = 3'h6 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_6_4 : _GEN_499; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_501 = 3'h6 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_6_5 : _GEN_500; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_502 = 3'h6 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_6_6 : _GEN_501; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_503 = 3'h6 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_6_7 : _GEN_502; // @[stationary_dpe.scala 94:{43,43}]
  wire  _GEN_2374 = 3'h7 == i[2:0]; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_504 = 3'h7 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_7_0 : _GEN_503; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_505 = 3'h7 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_7_1 : _GEN_504; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_506 = 3'h7 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_7_2 : _GEN_505; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_507 = 3'h7 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_7_3 : _GEN_506; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_508 = 3'h7 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_7_4 : _GEN_507; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_509 = 3'h7 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_7_5 : _GEN_508; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_510 = 3'h7 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_7_6 : _GEN_509; // @[stationary_dpe.scala 94:{43,43}]
  wire [15:0] _GEN_511 = 3'h7 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_7_7 : _GEN_510; // @[stationary_dpe.scala 94:{43,43}]
  wire [31:0] _count_T_1 = count + 32'h1; // @[stationary_dpe.scala 97:27]
  wire [31:0] _GEN_640 = _GEN_511 != 16'h0 ? _count_T_1 : count; // @[stationary_dpe.scala 94:51 97:18 23:27]
  wire [31:0] _GEN_705 = ~valid ? _GEN_640 : count; // @[stationary_dpe.scala 23:27 93:27]
  wire  valid1 = count >= 32'h10; // @[stationary_dpe.scala 194:18]
  wire [15:0] _GEN_707 = _GEN_2264 & _GEN_2265 ? Station2_0_1 : Station2_0_0; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_708 = _GEN_2264 & _GEN_2267 ? Station2_0_2 : _GEN_707; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_709 = _GEN_2264 & _GEN_2269 ? Station2_0_3 : _GEN_708; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_710 = _GEN_2264 & _GEN_2271 ? Station2_0_4 : _GEN_709; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_711 = _GEN_2264 & _GEN_2273 ? Station2_0_5 : _GEN_710; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_712 = _GEN_2264 & _GEN_2275 ? Station2_0_6 : _GEN_711; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_713 = _GEN_2264 & _GEN_2277 ? Station2_0_7 : _GEN_712; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_714 = _GEN_2278 & _GEN_2279 ? Station2_1_0 : _GEN_713; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_715 = _GEN_2278 & _GEN_2265 ? Station2_1_1 : _GEN_714; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_716 = _GEN_2278 & _GEN_2267 ? Station2_1_2 : _GEN_715; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_717 = _GEN_2278 & _GEN_2269 ? Station2_1_3 : _GEN_716; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_718 = _GEN_2278 & _GEN_2271 ? Station2_1_4 : _GEN_717; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_719 = _GEN_2278 & _GEN_2273 ? Station2_1_5 : _GEN_718; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_720 = _GEN_2278 & _GEN_2275 ? Station2_1_6 : _GEN_719; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_721 = _GEN_2278 & _GEN_2277 ? Station2_1_7 : _GEN_720; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_722 = _GEN_2294 & _GEN_2279 ? Station2_2_0 : _GEN_721; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_723 = _GEN_2294 & _GEN_2265 ? Station2_2_1 : _GEN_722; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_724 = _GEN_2294 & _GEN_2267 ? Station2_2_2 : _GEN_723; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_725 = _GEN_2294 & _GEN_2269 ? Station2_2_3 : _GEN_724; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_726 = _GEN_2294 & _GEN_2271 ? Station2_2_4 : _GEN_725; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_727 = _GEN_2294 & _GEN_2273 ? Station2_2_5 : _GEN_726; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_728 = _GEN_2294 & _GEN_2275 ? Station2_2_6 : _GEN_727; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_729 = _GEN_2294 & _GEN_2277 ? Station2_2_7 : _GEN_728; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_730 = _GEN_2310 & _GEN_2279 ? Station2_3_0 : _GEN_729; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_731 = _GEN_2310 & _GEN_2265 ? Station2_3_1 : _GEN_730; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_732 = _GEN_2310 & _GEN_2267 ? Station2_3_2 : _GEN_731; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_733 = _GEN_2310 & _GEN_2269 ? Station2_3_3 : _GEN_732; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_734 = _GEN_2310 & _GEN_2271 ? Station2_3_4 : _GEN_733; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_735 = _GEN_2310 & _GEN_2273 ? Station2_3_5 : _GEN_734; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_736 = _GEN_2310 & _GEN_2275 ? Station2_3_6 : _GEN_735; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_737 = _GEN_2310 & _GEN_2277 ? Station2_3_7 : _GEN_736; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_738 = _GEN_2326 & _GEN_2279 ? Station2_4_0 : _GEN_737; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_739 = _GEN_2326 & _GEN_2265 ? Station2_4_1 : _GEN_738; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_740 = _GEN_2326 & _GEN_2267 ? Station2_4_2 : _GEN_739; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_741 = _GEN_2326 & _GEN_2269 ? Station2_4_3 : _GEN_740; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_742 = _GEN_2326 & _GEN_2271 ? Station2_4_4 : _GEN_741; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_743 = _GEN_2326 & _GEN_2273 ? Station2_4_5 : _GEN_742; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_744 = _GEN_2326 & _GEN_2275 ? Station2_4_6 : _GEN_743; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_745 = _GEN_2326 & _GEN_2277 ? Station2_4_7 : _GEN_744; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_746 = _GEN_2342 & _GEN_2279 ? Station2_5_0 : _GEN_745; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_747 = _GEN_2342 & _GEN_2265 ? Station2_5_1 : _GEN_746; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_748 = _GEN_2342 & _GEN_2267 ? Station2_5_2 : _GEN_747; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_749 = _GEN_2342 & _GEN_2269 ? Station2_5_3 : _GEN_748; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_750 = _GEN_2342 & _GEN_2271 ? Station2_5_4 : _GEN_749; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_751 = _GEN_2342 & _GEN_2273 ? Station2_5_5 : _GEN_750; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_752 = _GEN_2342 & _GEN_2275 ? Station2_5_6 : _GEN_751; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_753 = _GEN_2342 & _GEN_2277 ? Station2_5_7 : _GEN_752; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_754 = _GEN_2358 & _GEN_2279 ? Station2_6_0 : _GEN_753; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_755 = _GEN_2358 & _GEN_2265 ? Station2_6_1 : _GEN_754; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_756 = _GEN_2358 & _GEN_2267 ? Station2_6_2 : _GEN_755; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_757 = _GEN_2358 & _GEN_2269 ? Station2_6_3 : _GEN_756; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_758 = _GEN_2358 & _GEN_2271 ? Station2_6_4 : _GEN_757; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_759 = _GEN_2358 & _GEN_2273 ? Station2_6_5 : _GEN_758; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_760 = _GEN_2358 & _GEN_2275 ? Station2_6_6 : _GEN_759; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_761 = _GEN_2358 & _GEN_2277 ? Station2_6_7 : _GEN_760; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_762 = _GEN_2374 & _GEN_2279 ? Station2_7_0 : _GEN_761; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_763 = _GEN_2374 & _GEN_2265 ? Station2_7_1 : _GEN_762; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_764 = _GEN_2374 & _GEN_2267 ? Station2_7_2 : _GEN_763; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_765 = _GEN_2374 & _GEN_2269 ? Station2_7_3 : _GEN_764; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_766 = _GEN_2374 & _GEN_2271 ? Station2_7_4 : _GEN_765; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_767 = _GEN_2374 & _GEN_2273 ? Station2_7_5 : _GEN_766; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_768 = _GEN_2374 & _GEN_2275 ? Station2_7_6 : _GEN_767; // @[stationary_dpe.scala 115:{31,31}]
  wire [15:0] _GEN_769 = _GEN_2374 & _GEN_2277 ? Station2_7_7 : _GEN_768; // @[stationary_dpe.scala 115:{31,31}]
  wire [31:0] _GEN_898 = _GEN_769 != 16'h0 ? _count_T_1 : _GEN_705; // @[stationary_dpe.scala 115:39 118:18]
  wire [31:0] _GEN_963 = ~valid1 ? _GEN_898 : _GEN_705; // @[stationary_dpe.scala 114:29]
  wire  valid2 = count >= 32'h18; // @[stationary_dpe.scala 198:17]
  wire [15:0] _GEN_965 = _GEN_2264 & _GEN_2265 ? Station3_0_1 : Station3_0_0; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_966 = _GEN_2264 & _GEN_2267 ? Station3_0_2 : _GEN_965; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_967 = _GEN_2264 & _GEN_2269 ? Station3_0_3 : _GEN_966; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_968 = _GEN_2264 & _GEN_2271 ? Station3_0_4 : _GEN_967; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_969 = _GEN_2264 & _GEN_2273 ? Station3_0_5 : _GEN_968; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_970 = _GEN_2264 & _GEN_2275 ? Station3_0_6 : _GEN_969; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_971 = _GEN_2264 & _GEN_2277 ? Station3_0_7 : _GEN_970; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_972 = _GEN_2278 & _GEN_2279 ? Station3_1_0 : _GEN_971; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_973 = _GEN_2278 & _GEN_2265 ? Station3_1_1 : _GEN_972; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_974 = _GEN_2278 & _GEN_2267 ? Station3_1_2 : _GEN_973; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_975 = _GEN_2278 & _GEN_2269 ? Station3_1_3 : _GEN_974; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_976 = _GEN_2278 & _GEN_2271 ? Station3_1_4 : _GEN_975; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_977 = _GEN_2278 & _GEN_2273 ? Station3_1_5 : _GEN_976; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_978 = _GEN_2278 & _GEN_2275 ? Station3_1_6 : _GEN_977; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_979 = _GEN_2278 & _GEN_2277 ? Station3_1_7 : _GEN_978; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_980 = _GEN_2294 & _GEN_2279 ? Station3_2_0 : _GEN_979; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_981 = _GEN_2294 & _GEN_2265 ? Station3_2_1 : _GEN_980; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_982 = _GEN_2294 & _GEN_2267 ? Station3_2_2 : _GEN_981; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_983 = _GEN_2294 & _GEN_2269 ? Station3_2_3 : _GEN_982; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_984 = _GEN_2294 & _GEN_2271 ? Station3_2_4 : _GEN_983; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_985 = _GEN_2294 & _GEN_2273 ? Station3_2_5 : _GEN_984; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_986 = _GEN_2294 & _GEN_2275 ? Station3_2_6 : _GEN_985; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_987 = _GEN_2294 & _GEN_2277 ? Station3_2_7 : _GEN_986; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_988 = _GEN_2310 & _GEN_2279 ? Station3_3_0 : _GEN_987; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_989 = _GEN_2310 & _GEN_2265 ? Station3_3_1 : _GEN_988; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_990 = _GEN_2310 & _GEN_2267 ? Station3_3_2 : _GEN_989; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_991 = _GEN_2310 & _GEN_2269 ? Station3_3_3 : _GEN_990; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_992 = _GEN_2310 & _GEN_2271 ? Station3_3_4 : _GEN_991; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_993 = _GEN_2310 & _GEN_2273 ? Station3_3_5 : _GEN_992; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_994 = _GEN_2310 & _GEN_2275 ? Station3_3_6 : _GEN_993; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_995 = _GEN_2310 & _GEN_2277 ? Station3_3_7 : _GEN_994; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_996 = _GEN_2326 & _GEN_2279 ? Station3_4_0 : _GEN_995; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_997 = _GEN_2326 & _GEN_2265 ? Station3_4_1 : _GEN_996; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_998 = _GEN_2326 & _GEN_2267 ? Station3_4_2 : _GEN_997; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_999 = _GEN_2326 & _GEN_2269 ? Station3_4_3 : _GEN_998; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_1000 = _GEN_2326 & _GEN_2271 ? Station3_4_4 : _GEN_999; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_1001 = _GEN_2326 & _GEN_2273 ? Station3_4_5 : _GEN_1000; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_1002 = _GEN_2326 & _GEN_2275 ? Station3_4_6 : _GEN_1001; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_1003 = _GEN_2326 & _GEN_2277 ? Station3_4_7 : _GEN_1002; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_1004 = _GEN_2342 & _GEN_2279 ? Station3_5_0 : _GEN_1003; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_1005 = _GEN_2342 & _GEN_2265 ? Station3_5_1 : _GEN_1004; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_1006 = _GEN_2342 & _GEN_2267 ? Station3_5_2 : _GEN_1005; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_1007 = _GEN_2342 & _GEN_2269 ? Station3_5_3 : _GEN_1006; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_1008 = _GEN_2342 & _GEN_2271 ? Station3_5_4 : _GEN_1007; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_1009 = _GEN_2342 & _GEN_2273 ? Station3_5_5 : _GEN_1008; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_1010 = _GEN_2342 & _GEN_2275 ? Station3_5_6 : _GEN_1009; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_1011 = _GEN_2342 & _GEN_2277 ? Station3_5_7 : _GEN_1010; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_1012 = _GEN_2358 & _GEN_2279 ? Station3_6_0 : _GEN_1011; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_1013 = _GEN_2358 & _GEN_2265 ? Station3_6_1 : _GEN_1012; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_1014 = _GEN_2358 & _GEN_2267 ? Station3_6_2 : _GEN_1013; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_1015 = _GEN_2358 & _GEN_2269 ? Station3_6_3 : _GEN_1014; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_1016 = _GEN_2358 & _GEN_2271 ? Station3_6_4 : _GEN_1015; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_1017 = _GEN_2358 & _GEN_2273 ? Station3_6_5 : _GEN_1016; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_1018 = _GEN_2358 & _GEN_2275 ? Station3_6_6 : _GEN_1017; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_1019 = _GEN_2358 & _GEN_2277 ? Station3_6_7 : _GEN_1018; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_1020 = _GEN_2374 & _GEN_2279 ? Station3_7_0 : _GEN_1019; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_1021 = _GEN_2374 & _GEN_2265 ? Station3_7_1 : _GEN_1020; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_1022 = _GEN_2374 & _GEN_2267 ? Station3_7_2 : _GEN_1021; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_1023 = _GEN_2374 & _GEN_2269 ? Station3_7_3 : _GEN_1022; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_1024 = _GEN_2374 & _GEN_2271 ? Station3_7_4 : _GEN_1023; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_1025 = _GEN_2374 & _GEN_2273 ? Station3_7_5 : _GEN_1024; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_1026 = _GEN_2374 & _GEN_2275 ? Station3_7_6 : _GEN_1025; // @[stationary_dpe.scala 127:{31,31}]
  wire [15:0] _GEN_1027 = _GEN_2374 & _GEN_2277 ? Station3_7_7 : _GEN_1026; // @[stationary_dpe.scala 127:{31,31}]
  wire [31:0] _GEN_1156 = _GEN_1027 != 16'h0 ? _count_T_1 : _GEN_963; // @[stationary_dpe.scala 127:39 130:18]
  wire [31:0] _GEN_1221 = ~valid2 ? _GEN_1156 : _GEN_963; // @[stationary_dpe.scala 126:29]
  wire  valid3 = count >= 32'h20; // @[stationary_dpe.scala 202:17]
  wire [15:0] _GEN_1223 = _GEN_2264 & _GEN_2265 ? Station4_0_1 : Station4_0_0; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1224 = _GEN_2264 & _GEN_2267 ? Station4_0_2 : _GEN_1223; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1225 = _GEN_2264 & _GEN_2269 ? Station4_0_3 : _GEN_1224; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1226 = _GEN_2264 & _GEN_2271 ? Station4_0_4 : _GEN_1225; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1227 = _GEN_2264 & _GEN_2273 ? Station4_0_5 : _GEN_1226; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1228 = _GEN_2264 & _GEN_2275 ? Station4_0_6 : _GEN_1227; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1229 = _GEN_2264 & _GEN_2277 ? Station4_0_7 : _GEN_1228; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1230 = _GEN_2278 & _GEN_2279 ? Station4_1_0 : _GEN_1229; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1231 = _GEN_2278 & _GEN_2265 ? Station4_1_1 : _GEN_1230; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1232 = _GEN_2278 & _GEN_2267 ? Station4_1_2 : _GEN_1231; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1233 = _GEN_2278 & _GEN_2269 ? Station4_1_3 : _GEN_1232; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1234 = _GEN_2278 & _GEN_2271 ? Station4_1_4 : _GEN_1233; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1235 = _GEN_2278 & _GEN_2273 ? Station4_1_5 : _GEN_1234; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1236 = _GEN_2278 & _GEN_2275 ? Station4_1_6 : _GEN_1235; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1237 = _GEN_2278 & _GEN_2277 ? Station4_1_7 : _GEN_1236; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1238 = _GEN_2294 & _GEN_2279 ? Station4_2_0 : _GEN_1237; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1239 = _GEN_2294 & _GEN_2265 ? Station4_2_1 : _GEN_1238; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1240 = _GEN_2294 & _GEN_2267 ? Station4_2_2 : _GEN_1239; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1241 = _GEN_2294 & _GEN_2269 ? Station4_2_3 : _GEN_1240; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1242 = _GEN_2294 & _GEN_2271 ? Station4_2_4 : _GEN_1241; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1243 = _GEN_2294 & _GEN_2273 ? Station4_2_5 : _GEN_1242; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1244 = _GEN_2294 & _GEN_2275 ? Station4_2_6 : _GEN_1243; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1245 = _GEN_2294 & _GEN_2277 ? Station4_2_7 : _GEN_1244; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1246 = _GEN_2310 & _GEN_2279 ? Station4_3_0 : _GEN_1245; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1247 = _GEN_2310 & _GEN_2265 ? Station4_3_1 : _GEN_1246; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1248 = _GEN_2310 & _GEN_2267 ? Station4_3_2 : _GEN_1247; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1249 = _GEN_2310 & _GEN_2269 ? Station4_3_3 : _GEN_1248; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1250 = _GEN_2310 & _GEN_2271 ? Station4_3_4 : _GEN_1249; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1251 = _GEN_2310 & _GEN_2273 ? Station4_3_5 : _GEN_1250; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1252 = _GEN_2310 & _GEN_2275 ? Station4_3_6 : _GEN_1251; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1253 = _GEN_2310 & _GEN_2277 ? Station4_3_7 : _GEN_1252; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1254 = _GEN_2326 & _GEN_2279 ? Station4_4_0 : _GEN_1253; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1255 = _GEN_2326 & _GEN_2265 ? Station4_4_1 : _GEN_1254; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1256 = _GEN_2326 & _GEN_2267 ? Station4_4_2 : _GEN_1255; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1257 = _GEN_2326 & _GEN_2269 ? Station4_4_3 : _GEN_1256; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1258 = _GEN_2326 & _GEN_2271 ? Station4_4_4 : _GEN_1257; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1259 = _GEN_2326 & _GEN_2273 ? Station4_4_5 : _GEN_1258; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1260 = _GEN_2326 & _GEN_2275 ? Station4_4_6 : _GEN_1259; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1261 = _GEN_2326 & _GEN_2277 ? Station4_4_7 : _GEN_1260; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1262 = _GEN_2342 & _GEN_2279 ? Station4_5_0 : _GEN_1261; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1263 = _GEN_2342 & _GEN_2265 ? Station4_5_1 : _GEN_1262; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1264 = _GEN_2342 & _GEN_2267 ? Station4_5_2 : _GEN_1263; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1265 = _GEN_2342 & _GEN_2269 ? Station4_5_3 : _GEN_1264; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1266 = _GEN_2342 & _GEN_2271 ? Station4_5_4 : _GEN_1265; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1267 = _GEN_2342 & _GEN_2273 ? Station4_5_5 : _GEN_1266; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1268 = _GEN_2342 & _GEN_2275 ? Station4_5_6 : _GEN_1267; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1269 = _GEN_2342 & _GEN_2277 ? Station4_5_7 : _GEN_1268; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1270 = _GEN_2358 & _GEN_2279 ? Station4_6_0 : _GEN_1269; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1271 = _GEN_2358 & _GEN_2265 ? Station4_6_1 : _GEN_1270; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1272 = _GEN_2358 & _GEN_2267 ? Station4_6_2 : _GEN_1271; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1273 = _GEN_2358 & _GEN_2269 ? Station4_6_3 : _GEN_1272; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1274 = _GEN_2358 & _GEN_2271 ? Station4_6_4 : _GEN_1273; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1275 = _GEN_2358 & _GEN_2273 ? Station4_6_5 : _GEN_1274; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1276 = _GEN_2358 & _GEN_2275 ? Station4_6_6 : _GEN_1275; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1277 = _GEN_2358 & _GEN_2277 ? Station4_6_7 : _GEN_1276; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1278 = _GEN_2374 & _GEN_2279 ? Station4_7_0 : _GEN_1277; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1279 = _GEN_2374 & _GEN_2265 ? Station4_7_1 : _GEN_1278; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1280 = _GEN_2374 & _GEN_2267 ? Station4_7_2 : _GEN_1279; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1281 = _GEN_2374 & _GEN_2269 ? Station4_7_3 : _GEN_1280; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1282 = _GEN_2374 & _GEN_2271 ? Station4_7_4 : _GEN_1281; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1283 = _GEN_2374 & _GEN_2273 ? Station4_7_5 : _GEN_1282; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1284 = _GEN_2374 & _GEN_2275 ? Station4_7_6 : _GEN_1283; // @[stationary_dpe.scala 139:{31,31}]
  wire [15:0] _GEN_1285 = _GEN_2374 & _GEN_2277 ? Station4_7_7 : _GEN_1284; // @[stationary_dpe.scala 139:{31,31}]
  wire [31:0] _GEN_1414 = _GEN_1285 != 16'h0 ? _count_T_1 : _GEN_1221; // @[stationary_dpe.scala 139:39 142:18]
  wire [31:0] _GEN_1479 = ~valid3 ? _GEN_1414 : _GEN_1221; // @[stationary_dpe.scala 138:28]
  wire  valid4 = count >= 32'h28; // @[stationary_dpe.scala 206:17]
  wire [15:0] _GEN_1481 = _GEN_2264 & _GEN_2265 ? Station5_0_1 : Station5_0_0; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1482 = _GEN_2264 & _GEN_2267 ? Station5_0_2 : _GEN_1481; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1483 = _GEN_2264 & _GEN_2269 ? Station5_0_3 : _GEN_1482; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1484 = _GEN_2264 & _GEN_2271 ? Station5_0_4 : _GEN_1483; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1485 = _GEN_2264 & _GEN_2273 ? Station5_0_5 : _GEN_1484; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1486 = _GEN_2264 & _GEN_2275 ? Station5_0_6 : _GEN_1485; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1487 = _GEN_2264 & _GEN_2277 ? Station5_0_7 : _GEN_1486; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1488 = _GEN_2278 & _GEN_2279 ? Station5_1_0 : _GEN_1487; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1489 = _GEN_2278 & _GEN_2265 ? Station5_1_1 : _GEN_1488; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1490 = _GEN_2278 & _GEN_2267 ? Station5_1_2 : _GEN_1489; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1491 = _GEN_2278 & _GEN_2269 ? Station5_1_3 : _GEN_1490; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1492 = _GEN_2278 & _GEN_2271 ? Station5_1_4 : _GEN_1491; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1493 = _GEN_2278 & _GEN_2273 ? Station5_1_5 : _GEN_1492; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1494 = _GEN_2278 & _GEN_2275 ? Station5_1_6 : _GEN_1493; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1495 = _GEN_2278 & _GEN_2277 ? Station5_1_7 : _GEN_1494; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1496 = _GEN_2294 & _GEN_2279 ? Station5_2_0 : _GEN_1495; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1497 = _GEN_2294 & _GEN_2265 ? Station5_2_1 : _GEN_1496; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1498 = _GEN_2294 & _GEN_2267 ? Station5_2_2 : _GEN_1497; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1499 = _GEN_2294 & _GEN_2269 ? Station5_2_3 : _GEN_1498; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1500 = _GEN_2294 & _GEN_2271 ? Station5_2_4 : _GEN_1499; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1501 = _GEN_2294 & _GEN_2273 ? Station5_2_5 : _GEN_1500; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1502 = _GEN_2294 & _GEN_2275 ? Station5_2_6 : _GEN_1501; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1503 = _GEN_2294 & _GEN_2277 ? Station5_2_7 : _GEN_1502; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1504 = _GEN_2310 & _GEN_2279 ? Station5_3_0 : _GEN_1503; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1505 = _GEN_2310 & _GEN_2265 ? Station5_3_1 : _GEN_1504; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1506 = _GEN_2310 & _GEN_2267 ? Station5_3_2 : _GEN_1505; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1507 = _GEN_2310 & _GEN_2269 ? Station5_3_3 : _GEN_1506; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1508 = _GEN_2310 & _GEN_2271 ? Station5_3_4 : _GEN_1507; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1509 = _GEN_2310 & _GEN_2273 ? Station5_3_5 : _GEN_1508; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1510 = _GEN_2310 & _GEN_2275 ? Station5_3_6 : _GEN_1509; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1511 = _GEN_2310 & _GEN_2277 ? Station5_3_7 : _GEN_1510; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1512 = _GEN_2326 & _GEN_2279 ? Station5_4_0 : _GEN_1511; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1513 = _GEN_2326 & _GEN_2265 ? Station5_4_1 : _GEN_1512; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1514 = _GEN_2326 & _GEN_2267 ? Station5_4_2 : _GEN_1513; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1515 = _GEN_2326 & _GEN_2269 ? Station5_4_3 : _GEN_1514; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1516 = _GEN_2326 & _GEN_2271 ? Station5_4_4 : _GEN_1515; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1517 = _GEN_2326 & _GEN_2273 ? Station5_4_5 : _GEN_1516; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1518 = _GEN_2326 & _GEN_2275 ? Station5_4_6 : _GEN_1517; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1519 = _GEN_2326 & _GEN_2277 ? Station5_4_7 : _GEN_1518; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1520 = _GEN_2342 & _GEN_2279 ? Station5_5_0 : _GEN_1519; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1521 = _GEN_2342 & _GEN_2265 ? Station5_5_1 : _GEN_1520; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1522 = _GEN_2342 & _GEN_2267 ? Station5_5_2 : _GEN_1521; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1523 = _GEN_2342 & _GEN_2269 ? Station5_5_3 : _GEN_1522; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1524 = _GEN_2342 & _GEN_2271 ? Station5_5_4 : _GEN_1523; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1525 = _GEN_2342 & _GEN_2273 ? Station5_5_5 : _GEN_1524; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1526 = _GEN_2342 & _GEN_2275 ? Station5_5_6 : _GEN_1525; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1527 = _GEN_2342 & _GEN_2277 ? Station5_5_7 : _GEN_1526; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1528 = _GEN_2358 & _GEN_2279 ? Station5_6_0 : _GEN_1527; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1529 = _GEN_2358 & _GEN_2265 ? Station5_6_1 : _GEN_1528; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1530 = _GEN_2358 & _GEN_2267 ? Station5_6_2 : _GEN_1529; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1531 = _GEN_2358 & _GEN_2269 ? Station5_6_3 : _GEN_1530; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1532 = _GEN_2358 & _GEN_2271 ? Station5_6_4 : _GEN_1531; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1533 = _GEN_2358 & _GEN_2273 ? Station5_6_5 : _GEN_1532; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1534 = _GEN_2358 & _GEN_2275 ? Station5_6_6 : _GEN_1533; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1535 = _GEN_2358 & _GEN_2277 ? Station5_6_7 : _GEN_1534; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1536 = _GEN_2374 & _GEN_2279 ? Station5_7_0 : _GEN_1535; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1537 = _GEN_2374 & _GEN_2265 ? Station5_7_1 : _GEN_1536; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1538 = _GEN_2374 & _GEN_2267 ? Station5_7_2 : _GEN_1537; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1539 = _GEN_2374 & _GEN_2269 ? Station5_7_3 : _GEN_1538; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1540 = _GEN_2374 & _GEN_2271 ? Station5_7_4 : _GEN_1539; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1541 = _GEN_2374 & _GEN_2273 ? Station5_7_5 : _GEN_1540; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1542 = _GEN_2374 & _GEN_2275 ? Station5_7_6 : _GEN_1541; // @[stationary_dpe.scala 151:{31,31}]
  wire [15:0] _GEN_1543 = _GEN_2374 & _GEN_2277 ? Station5_7_7 : _GEN_1542; // @[stationary_dpe.scala 151:{31,31}]
  wire [31:0] _GEN_1672 = _GEN_1543 != 16'h0 ? _count_T_1 : _GEN_1479; // @[stationary_dpe.scala 151:39 154:18]
  wire [31:0] _GEN_1737 = ~valid4 ? _GEN_1672 : _GEN_1479; // @[stationary_dpe.scala 150:28]
  wire  valid5 = count >= 32'h30; // @[stationary_dpe.scala 210:17]
  wire [15:0] _GEN_1739 = _GEN_2264 & _GEN_2265 ? Station6_0_1 : Station6_0_0; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1740 = _GEN_2264 & _GEN_2267 ? Station6_0_2 : _GEN_1739; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1741 = _GEN_2264 & _GEN_2269 ? Station6_0_3 : _GEN_1740; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1742 = _GEN_2264 & _GEN_2271 ? Station6_0_4 : _GEN_1741; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1743 = _GEN_2264 & _GEN_2273 ? Station6_0_5 : _GEN_1742; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1744 = _GEN_2264 & _GEN_2275 ? Station6_0_6 : _GEN_1743; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1745 = _GEN_2264 & _GEN_2277 ? Station6_0_7 : _GEN_1744; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1746 = _GEN_2278 & _GEN_2279 ? Station6_1_0 : _GEN_1745; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1747 = _GEN_2278 & _GEN_2265 ? Station6_1_1 : _GEN_1746; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1748 = _GEN_2278 & _GEN_2267 ? Station6_1_2 : _GEN_1747; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1749 = _GEN_2278 & _GEN_2269 ? Station6_1_3 : _GEN_1748; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1750 = _GEN_2278 & _GEN_2271 ? Station6_1_4 : _GEN_1749; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1751 = _GEN_2278 & _GEN_2273 ? Station6_1_5 : _GEN_1750; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1752 = _GEN_2278 & _GEN_2275 ? Station6_1_6 : _GEN_1751; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1753 = _GEN_2278 & _GEN_2277 ? Station6_1_7 : _GEN_1752; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1754 = _GEN_2294 & _GEN_2279 ? Station6_2_0 : _GEN_1753; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1755 = _GEN_2294 & _GEN_2265 ? Station6_2_1 : _GEN_1754; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1756 = _GEN_2294 & _GEN_2267 ? Station6_2_2 : _GEN_1755; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1757 = _GEN_2294 & _GEN_2269 ? Station6_2_3 : _GEN_1756; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1758 = _GEN_2294 & _GEN_2271 ? Station6_2_4 : _GEN_1757; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1759 = _GEN_2294 & _GEN_2273 ? Station6_2_5 : _GEN_1758; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1760 = _GEN_2294 & _GEN_2275 ? Station6_2_6 : _GEN_1759; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1761 = _GEN_2294 & _GEN_2277 ? Station6_2_7 : _GEN_1760; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1762 = _GEN_2310 & _GEN_2279 ? Station6_3_0 : _GEN_1761; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1763 = _GEN_2310 & _GEN_2265 ? Station6_3_1 : _GEN_1762; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1764 = _GEN_2310 & _GEN_2267 ? Station6_3_2 : _GEN_1763; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1765 = _GEN_2310 & _GEN_2269 ? Station6_3_3 : _GEN_1764; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1766 = _GEN_2310 & _GEN_2271 ? Station6_3_4 : _GEN_1765; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1767 = _GEN_2310 & _GEN_2273 ? Station6_3_5 : _GEN_1766; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1768 = _GEN_2310 & _GEN_2275 ? Station6_3_6 : _GEN_1767; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1769 = _GEN_2310 & _GEN_2277 ? Station6_3_7 : _GEN_1768; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1770 = _GEN_2326 & _GEN_2279 ? Station6_4_0 : _GEN_1769; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1771 = _GEN_2326 & _GEN_2265 ? Station6_4_1 : _GEN_1770; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1772 = _GEN_2326 & _GEN_2267 ? Station6_4_2 : _GEN_1771; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1773 = _GEN_2326 & _GEN_2269 ? Station6_4_3 : _GEN_1772; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1774 = _GEN_2326 & _GEN_2271 ? Station6_4_4 : _GEN_1773; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1775 = _GEN_2326 & _GEN_2273 ? Station6_4_5 : _GEN_1774; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1776 = _GEN_2326 & _GEN_2275 ? Station6_4_6 : _GEN_1775; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1777 = _GEN_2326 & _GEN_2277 ? Station6_4_7 : _GEN_1776; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1778 = _GEN_2342 & _GEN_2279 ? Station6_5_0 : _GEN_1777; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1779 = _GEN_2342 & _GEN_2265 ? Station6_5_1 : _GEN_1778; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1780 = _GEN_2342 & _GEN_2267 ? Station6_5_2 : _GEN_1779; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1781 = _GEN_2342 & _GEN_2269 ? Station6_5_3 : _GEN_1780; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1782 = _GEN_2342 & _GEN_2271 ? Station6_5_4 : _GEN_1781; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1783 = _GEN_2342 & _GEN_2273 ? Station6_5_5 : _GEN_1782; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1784 = _GEN_2342 & _GEN_2275 ? Station6_5_6 : _GEN_1783; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1785 = _GEN_2342 & _GEN_2277 ? Station6_5_7 : _GEN_1784; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1786 = _GEN_2358 & _GEN_2279 ? Station6_6_0 : _GEN_1785; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1787 = _GEN_2358 & _GEN_2265 ? Station6_6_1 : _GEN_1786; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1788 = _GEN_2358 & _GEN_2267 ? Station6_6_2 : _GEN_1787; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1789 = _GEN_2358 & _GEN_2269 ? Station6_6_3 : _GEN_1788; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1790 = _GEN_2358 & _GEN_2271 ? Station6_6_4 : _GEN_1789; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1791 = _GEN_2358 & _GEN_2273 ? Station6_6_5 : _GEN_1790; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1792 = _GEN_2358 & _GEN_2275 ? Station6_6_6 : _GEN_1791; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1793 = _GEN_2358 & _GEN_2277 ? Station6_6_7 : _GEN_1792; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1794 = _GEN_2374 & _GEN_2279 ? Station6_7_0 : _GEN_1793; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1795 = _GEN_2374 & _GEN_2265 ? Station6_7_1 : _GEN_1794; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1796 = _GEN_2374 & _GEN_2267 ? Station6_7_2 : _GEN_1795; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1797 = _GEN_2374 & _GEN_2269 ? Station6_7_3 : _GEN_1796; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1798 = _GEN_2374 & _GEN_2271 ? Station6_7_4 : _GEN_1797; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1799 = _GEN_2374 & _GEN_2273 ? Station6_7_5 : _GEN_1798; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1800 = _GEN_2374 & _GEN_2275 ? Station6_7_6 : _GEN_1799; // @[stationary_dpe.scala 163:{31,31}]
  wire [15:0] _GEN_1801 = _GEN_2374 & _GEN_2277 ? Station6_7_7 : _GEN_1800; // @[stationary_dpe.scala 163:{31,31}]
  wire [31:0] _GEN_1930 = _GEN_1801 != 16'h0 ? _count_T_1 : _GEN_1737; // @[stationary_dpe.scala 163:39 166:18]
  wire [31:0] _GEN_1995 = ~valid5 ? _GEN_1930 : _GEN_1737; // @[stationary_dpe.scala 162:28]
  wire  valid6 = count >= 32'h38; // @[stationary_dpe.scala 215:17]
  wire [15:0] _GEN_1997 = _GEN_2264 & _GEN_2265 ? Station7_0_1 : Station7_0_0; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_1998 = _GEN_2264 & _GEN_2267 ? Station7_0_2 : _GEN_1997; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_1999 = _GEN_2264 & _GEN_2269 ? Station7_0_3 : _GEN_1998; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2000 = _GEN_2264 & _GEN_2271 ? Station7_0_4 : _GEN_1999; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2001 = _GEN_2264 & _GEN_2273 ? Station7_0_5 : _GEN_2000; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2002 = _GEN_2264 & _GEN_2275 ? Station7_0_6 : _GEN_2001; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2003 = _GEN_2264 & _GEN_2277 ? Station7_0_7 : _GEN_2002; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2004 = _GEN_2278 & _GEN_2279 ? Station7_1_0 : _GEN_2003; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2005 = _GEN_2278 & _GEN_2265 ? Station7_1_1 : _GEN_2004; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2006 = _GEN_2278 & _GEN_2267 ? Station7_1_2 : _GEN_2005; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2007 = _GEN_2278 & _GEN_2269 ? Station7_1_3 : _GEN_2006; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2008 = _GEN_2278 & _GEN_2271 ? Station7_1_4 : _GEN_2007; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2009 = _GEN_2278 & _GEN_2273 ? Station7_1_5 : _GEN_2008; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2010 = _GEN_2278 & _GEN_2275 ? Station7_1_6 : _GEN_2009; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2011 = _GEN_2278 & _GEN_2277 ? Station7_1_7 : _GEN_2010; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2012 = _GEN_2294 & _GEN_2279 ? Station7_2_0 : _GEN_2011; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2013 = _GEN_2294 & _GEN_2265 ? Station7_2_1 : _GEN_2012; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2014 = _GEN_2294 & _GEN_2267 ? Station7_2_2 : _GEN_2013; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2015 = _GEN_2294 & _GEN_2269 ? Station7_2_3 : _GEN_2014; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2016 = _GEN_2294 & _GEN_2271 ? Station7_2_4 : _GEN_2015; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2017 = _GEN_2294 & _GEN_2273 ? Station7_2_5 : _GEN_2016; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2018 = _GEN_2294 & _GEN_2275 ? Station7_2_6 : _GEN_2017; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2019 = _GEN_2294 & _GEN_2277 ? Station7_2_7 : _GEN_2018; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2020 = _GEN_2310 & _GEN_2279 ? Station7_3_0 : _GEN_2019; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2021 = _GEN_2310 & _GEN_2265 ? Station7_3_1 : _GEN_2020; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2022 = _GEN_2310 & _GEN_2267 ? Station7_3_2 : _GEN_2021; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2023 = _GEN_2310 & _GEN_2269 ? Station7_3_3 : _GEN_2022; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2024 = _GEN_2310 & _GEN_2271 ? Station7_3_4 : _GEN_2023; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2025 = _GEN_2310 & _GEN_2273 ? Station7_3_5 : _GEN_2024; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2026 = _GEN_2310 & _GEN_2275 ? Station7_3_6 : _GEN_2025; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2027 = _GEN_2310 & _GEN_2277 ? Station7_3_7 : _GEN_2026; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2028 = _GEN_2326 & _GEN_2279 ? Station7_4_0 : _GEN_2027; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2029 = _GEN_2326 & _GEN_2265 ? Station7_4_1 : _GEN_2028; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2030 = _GEN_2326 & _GEN_2267 ? Station7_4_2 : _GEN_2029; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2031 = _GEN_2326 & _GEN_2269 ? Station7_4_3 : _GEN_2030; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2032 = _GEN_2326 & _GEN_2271 ? Station7_4_4 : _GEN_2031; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2033 = _GEN_2326 & _GEN_2273 ? Station7_4_5 : _GEN_2032; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2034 = _GEN_2326 & _GEN_2275 ? Station7_4_6 : _GEN_2033; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2035 = _GEN_2326 & _GEN_2277 ? Station7_4_7 : _GEN_2034; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2036 = _GEN_2342 & _GEN_2279 ? Station7_5_0 : _GEN_2035; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2037 = _GEN_2342 & _GEN_2265 ? Station7_5_1 : _GEN_2036; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2038 = _GEN_2342 & _GEN_2267 ? Station7_5_2 : _GEN_2037; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2039 = _GEN_2342 & _GEN_2269 ? Station7_5_3 : _GEN_2038; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2040 = _GEN_2342 & _GEN_2271 ? Station7_5_4 : _GEN_2039; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2041 = _GEN_2342 & _GEN_2273 ? Station7_5_5 : _GEN_2040; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2042 = _GEN_2342 & _GEN_2275 ? Station7_5_6 : _GEN_2041; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2043 = _GEN_2342 & _GEN_2277 ? Station7_5_7 : _GEN_2042; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2044 = _GEN_2358 & _GEN_2279 ? Station7_6_0 : _GEN_2043; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2045 = _GEN_2358 & _GEN_2265 ? Station7_6_1 : _GEN_2044; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2046 = _GEN_2358 & _GEN_2267 ? Station7_6_2 : _GEN_2045; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2047 = _GEN_2358 & _GEN_2269 ? Station7_6_3 : _GEN_2046; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2048 = _GEN_2358 & _GEN_2271 ? Station7_6_4 : _GEN_2047; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2049 = _GEN_2358 & _GEN_2273 ? Station7_6_5 : _GEN_2048; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2050 = _GEN_2358 & _GEN_2275 ? Station7_6_6 : _GEN_2049; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2051 = _GEN_2358 & _GEN_2277 ? Station7_6_7 : _GEN_2050; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2052 = _GEN_2374 & _GEN_2279 ? Station7_7_0 : _GEN_2051; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2053 = _GEN_2374 & _GEN_2265 ? Station7_7_1 : _GEN_2052; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2054 = _GEN_2374 & _GEN_2267 ? Station7_7_2 : _GEN_2053; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2055 = _GEN_2374 & _GEN_2269 ? Station7_7_3 : _GEN_2054; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2056 = _GEN_2374 & _GEN_2271 ? Station7_7_4 : _GEN_2055; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2057 = _GEN_2374 & _GEN_2273 ? Station7_7_5 : _GEN_2056; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2058 = _GEN_2374 & _GEN_2275 ? Station7_7_6 : _GEN_2057; // @[stationary_dpe.scala 175:{31,31}]
  wire [15:0] _GEN_2059 = _GEN_2374 & _GEN_2277 ? Station7_7_7 : _GEN_2058; // @[stationary_dpe.scala 175:{31,31}]
  wire  _T_57 = j == 32'h7; // @[stationary_dpe.scala 222:46]
  wire [31:0] _i_T_1 = i + 32'h1; // @[stationary_dpe.scala 223:16]
  wire [31:0] _j_T_1 = j + 32'h1; // @[stationary_dpe.scala 227:16]
  assign io_o_Stationary_matrix1_0_0 = io_Stationary_matrix_0_0; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_0_1 = io_Stationary_matrix_0_1; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_0_2 = io_Stationary_matrix_0_2; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_0_3 = io_Stationary_matrix_0_3; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_0_4 = io_Stationary_matrix_0_4; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_0_5 = io_Stationary_matrix_0_5; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_0_6 = io_Stationary_matrix_0_6; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_0_7 = io_Stationary_matrix_0_7; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_1_0 = io_Stationary_matrix_1_0; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_1_1 = io_Stationary_matrix_1_1; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_1_2 = io_Stationary_matrix_1_2; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_1_3 = io_Stationary_matrix_1_3; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_1_4 = io_Stationary_matrix_1_4; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_1_5 = io_Stationary_matrix_1_5; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_1_6 = io_Stationary_matrix_1_6; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_1_7 = io_Stationary_matrix_1_7; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_2_0 = io_Stationary_matrix_2_0; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_2_1 = io_Stationary_matrix_2_1; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_2_2 = io_Stationary_matrix_2_2; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_2_3 = io_Stationary_matrix_2_3; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_2_4 = io_Stationary_matrix_2_4; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_2_5 = io_Stationary_matrix_2_5; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_2_6 = io_Stationary_matrix_2_6; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_2_7 = io_Stationary_matrix_2_7; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_3_0 = io_Stationary_matrix_3_0; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_3_1 = io_Stationary_matrix_3_1; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_3_2 = io_Stationary_matrix_3_2; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_3_3 = io_Stationary_matrix_3_3; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_3_4 = io_Stationary_matrix_3_4; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_3_5 = io_Stationary_matrix_3_5; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_3_6 = io_Stationary_matrix_3_6; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_3_7 = io_Stationary_matrix_3_7; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_4_0 = io_Stationary_matrix_4_0; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_4_1 = io_Stationary_matrix_4_1; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_4_2 = io_Stationary_matrix_4_2; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_4_3 = io_Stationary_matrix_4_3; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_4_4 = io_Stationary_matrix_4_4; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_4_5 = io_Stationary_matrix_4_5; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_4_6 = io_Stationary_matrix_4_6; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_4_7 = io_Stationary_matrix_4_7; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_5_0 = io_Stationary_matrix_5_0; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_5_1 = io_Stationary_matrix_5_1; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_5_2 = io_Stationary_matrix_5_2; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_5_3 = io_Stationary_matrix_5_3; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_5_4 = io_Stationary_matrix_5_4; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_5_5 = io_Stationary_matrix_5_5; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_5_6 = io_Stationary_matrix_5_6; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_5_7 = io_Stationary_matrix_5_7; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_6_0 = io_Stationary_matrix_6_0; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_6_1 = io_Stationary_matrix_6_1; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_6_2 = io_Stationary_matrix_6_2; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_6_3 = io_Stationary_matrix_6_3; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_6_4 = io_Stationary_matrix_6_4; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_6_5 = io_Stationary_matrix_6_5; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_6_6 = io_Stationary_matrix_6_6; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_6_7 = io_Stationary_matrix_6_7; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_7_0 = io_Stationary_matrix_7_0; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_7_1 = io_Stationary_matrix_7_1; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_7_2 = io_Stationary_matrix_7_2; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_7_3 = io_Stationary_matrix_7_3; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_7_4 = io_Stationary_matrix_7_4; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_7_5 = io_Stationary_matrix_7_5; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_7_6 = io_Stationary_matrix_7_6; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix1_7_7 = io_Stationary_matrix_7_7; // @[stationary_dpe.scala 24:29]
  assign io_o_Stationary_matrix2_0_0 = Station2_0_0; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_0_1 = Station2_0_1; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_0_2 = Station2_0_2; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_0_3 = Station2_0_3; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_0_4 = Station2_0_4; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_0_5 = Station2_0_5; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_0_6 = Station2_0_6; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_0_7 = Station2_0_7; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_1_0 = Station2_1_0; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_1_1 = Station2_1_1; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_1_2 = Station2_1_2; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_1_3 = Station2_1_3; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_1_4 = Station2_1_4; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_1_5 = Station2_1_5; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_1_6 = Station2_1_6; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_1_7 = Station2_1_7; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_2_0 = Station2_2_0; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_2_1 = Station2_2_1; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_2_2 = Station2_2_2; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_2_3 = Station2_2_3; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_2_4 = Station2_2_4; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_2_5 = Station2_2_5; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_2_6 = Station2_2_6; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_2_7 = Station2_2_7; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_3_0 = Station2_3_0; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_3_1 = Station2_3_1; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_3_2 = Station2_3_2; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_3_3 = Station2_3_3; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_3_4 = Station2_3_4; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_3_5 = Station2_3_5; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_3_6 = Station2_3_6; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_3_7 = Station2_3_7; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_4_0 = Station2_4_0; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_4_1 = Station2_4_1; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_4_2 = Station2_4_2; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_4_3 = Station2_4_3; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_4_4 = Station2_4_4; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_4_5 = Station2_4_5; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_4_6 = Station2_4_6; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_4_7 = Station2_4_7; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_5_0 = Station2_5_0; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_5_1 = Station2_5_1; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_5_2 = Station2_5_2; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_5_3 = Station2_5_3; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_5_4 = Station2_5_4; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_5_5 = Station2_5_5; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_5_6 = Station2_5_6; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_5_7 = Station2_5_7; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_6_0 = Station2_6_0; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_6_1 = Station2_6_1; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_6_2 = Station2_6_2; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_6_3 = Station2_6_3; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_6_4 = Station2_6_4; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_6_5 = Station2_6_5; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_6_6 = Station2_6_6; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_6_7 = Station2_6_7; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_7_0 = Station2_7_0; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_7_1 = Station2_7_1; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_7_2 = Station2_7_2; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_7_3 = Station2_7_3; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_7_4 = Station2_7_4; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_7_5 = Station2_7_5; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_7_6 = Station2_7_6; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix2_7_7 = Station2_7_7; // @[stationary_dpe.scala 106:29]
  assign io_o_Stationary_matrix3_0_0 = Station3_0_0; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_0_1 = Station3_0_1; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_0_2 = Station3_0_2; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_0_3 = Station3_0_3; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_0_4 = Station3_0_4; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_0_5 = Station3_0_5; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_0_6 = Station3_0_6; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_0_7 = Station3_0_7; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_1_0 = Station3_1_0; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_1_1 = Station3_1_1; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_1_2 = Station3_1_2; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_1_3 = Station3_1_3; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_1_4 = Station3_1_4; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_1_5 = Station3_1_5; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_1_6 = Station3_1_6; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_1_7 = Station3_1_7; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_2_0 = Station3_2_0; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_2_1 = Station3_2_1; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_2_2 = Station3_2_2; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_2_3 = Station3_2_3; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_2_4 = Station3_2_4; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_2_5 = Station3_2_5; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_2_6 = Station3_2_6; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_2_7 = Station3_2_7; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_3_0 = Station3_3_0; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_3_1 = Station3_3_1; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_3_2 = Station3_3_2; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_3_3 = Station3_3_3; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_3_4 = Station3_3_4; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_3_5 = Station3_3_5; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_3_6 = Station3_3_6; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_3_7 = Station3_3_7; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_4_0 = Station3_4_0; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_4_1 = Station3_4_1; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_4_2 = Station3_4_2; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_4_3 = Station3_4_3; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_4_4 = Station3_4_4; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_4_5 = Station3_4_5; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_4_6 = Station3_4_6; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_4_7 = Station3_4_7; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_5_0 = Station3_5_0; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_5_1 = Station3_5_1; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_5_2 = Station3_5_2; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_5_3 = Station3_5_3; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_5_4 = Station3_5_4; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_5_5 = Station3_5_5; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_5_6 = Station3_5_6; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_5_7 = Station3_5_7; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_6_0 = Station3_6_0; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_6_1 = Station3_6_1; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_6_2 = Station3_6_2; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_6_3 = Station3_6_3; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_6_4 = Station3_6_4; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_6_5 = Station3_6_5; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_6_6 = Station3_6_6; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_6_7 = Station3_6_7; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_7_0 = Station3_7_0; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_7_1 = Station3_7_1; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_7_2 = Station3_7_2; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_7_3 = Station3_7_3; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_7_4 = Station3_7_4; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_7_5 = Station3_7_5; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_7_6 = Station3_7_6; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix3_7_7 = Station3_7_7; // @[stationary_dpe.scala 124:29]
  assign io_o_Stationary_matrix4_0_0 = Station4_0_0; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_0_1 = Station4_0_1; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_0_2 = Station4_0_2; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_0_3 = Station4_0_3; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_0_4 = Station4_0_4; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_0_5 = Station4_0_5; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_0_6 = Station4_0_6; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_0_7 = Station4_0_7; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_1_0 = Station4_1_0; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_1_1 = Station4_1_1; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_1_2 = Station4_1_2; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_1_3 = Station4_1_3; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_1_4 = Station4_1_4; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_1_5 = Station4_1_5; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_1_6 = Station4_1_6; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_1_7 = Station4_1_7; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_2_0 = Station4_2_0; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_2_1 = Station4_2_1; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_2_2 = Station4_2_2; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_2_3 = Station4_2_3; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_2_4 = Station4_2_4; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_2_5 = Station4_2_5; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_2_6 = Station4_2_6; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_2_7 = Station4_2_7; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_3_0 = Station4_3_0; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_3_1 = Station4_3_1; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_3_2 = Station4_3_2; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_3_3 = Station4_3_3; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_3_4 = Station4_3_4; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_3_5 = Station4_3_5; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_3_6 = Station4_3_6; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_3_7 = Station4_3_7; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_4_0 = Station4_4_0; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_4_1 = Station4_4_1; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_4_2 = Station4_4_2; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_4_3 = Station4_4_3; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_4_4 = Station4_4_4; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_4_5 = Station4_4_5; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_4_6 = Station4_4_6; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_4_7 = Station4_4_7; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_5_0 = Station4_5_0; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_5_1 = Station4_5_1; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_5_2 = Station4_5_2; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_5_3 = Station4_5_3; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_5_4 = Station4_5_4; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_5_5 = Station4_5_5; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_5_6 = Station4_5_6; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_5_7 = Station4_5_7; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_6_0 = Station4_6_0; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_6_1 = Station4_6_1; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_6_2 = Station4_6_2; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_6_3 = Station4_6_3; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_6_4 = Station4_6_4; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_6_5 = Station4_6_5; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_6_6 = Station4_6_6; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_6_7 = Station4_6_7; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_7_0 = Station4_7_0; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_7_1 = Station4_7_1; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_7_2 = Station4_7_2; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_7_3 = Station4_7_3; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_7_4 = Station4_7_4; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_7_5 = Station4_7_5; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_7_6 = Station4_7_6; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix4_7_7 = Station4_7_7; // @[stationary_dpe.scala 136:29]
  assign io_o_Stationary_matrix5_0_0 = Station5_0_0; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_0_1 = Station5_0_1; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_0_2 = Station5_0_2; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_0_3 = Station5_0_3; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_0_4 = Station5_0_4; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_0_5 = Station5_0_5; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_0_6 = Station5_0_6; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_0_7 = Station5_0_7; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_1_0 = Station5_1_0; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_1_1 = Station5_1_1; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_1_2 = Station5_1_2; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_1_3 = Station5_1_3; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_1_4 = Station5_1_4; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_1_5 = Station5_1_5; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_1_6 = Station5_1_6; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_1_7 = Station5_1_7; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_2_0 = Station5_2_0; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_2_1 = Station5_2_1; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_2_2 = Station5_2_2; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_2_3 = Station5_2_3; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_2_4 = Station5_2_4; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_2_5 = Station5_2_5; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_2_6 = Station5_2_6; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_2_7 = Station5_2_7; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_3_0 = Station5_3_0; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_3_1 = Station5_3_1; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_3_2 = Station5_3_2; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_3_3 = Station5_3_3; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_3_4 = Station5_3_4; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_3_5 = Station5_3_5; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_3_6 = Station5_3_6; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_3_7 = Station5_3_7; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_4_0 = Station5_4_0; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_4_1 = Station5_4_1; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_4_2 = Station5_4_2; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_4_3 = Station5_4_3; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_4_4 = Station5_4_4; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_4_5 = Station5_4_5; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_4_6 = Station5_4_6; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_4_7 = Station5_4_7; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_5_0 = Station5_5_0; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_5_1 = Station5_5_1; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_5_2 = Station5_5_2; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_5_3 = Station5_5_3; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_5_4 = Station5_5_4; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_5_5 = Station5_5_5; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_5_6 = Station5_5_6; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_5_7 = Station5_5_7; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_6_0 = Station5_6_0; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_6_1 = Station5_6_1; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_6_2 = Station5_6_2; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_6_3 = Station5_6_3; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_6_4 = Station5_6_4; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_6_5 = Station5_6_5; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_6_6 = Station5_6_6; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_6_7 = Station5_6_7; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_7_0 = Station5_7_0; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_7_1 = Station5_7_1; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_7_2 = Station5_7_2; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_7_3 = Station5_7_3; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_7_4 = Station5_7_4; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_7_5 = Station5_7_5; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_7_6 = Station5_7_6; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix5_7_7 = Station5_7_7; // @[stationary_dpe.scala 148:29]
  assign io_o_Stationary_matrix6_0_0 = Station6_0_0; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_0_1 = Station6_0_1; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_0_2 = Station6_0_2; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_0_3 = Station6_0_3; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_0_4 = Station6_0_4; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_0_5 = Station6_0_5; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_0_6 = Station6_0_6; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_0_7 = Station6_0_7; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_1_0 = Station6_1_0; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_1_1 = Station6_1_1; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_1_2 = Station6_1_2; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_1_3 = Station6_1_3; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_1_4 = Station6_1_4; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_1_5 = Station6_1_5; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_1_6 = Station6_1_6; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_1_7 = Station6_1_7; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_2_0 = Station6_2_0; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_2_1 = Station6_2_1; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_2_2 = Station6_2_2; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_2_3 = Station6_2_3; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_2_4 = Station6_2_4; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_2_5 = Station6_2_5; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_2_6 = Station6_2_6; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_2_7 = Station6_2_7; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_3_0 = Station6_3_0; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_3_1 = Station6_3_1; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_3_2 = Station6_3_2; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_3_3 = Station6_3_3; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_3_4 = Station6_3_4; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_3_5 = Station6_3_5; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_3_6 = Station6_3_6; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_3_7 = Station6_3_7; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_4_0 = Station6_4_0; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_4_1 = Station6_4_1; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_4_2 = Station6_4_2; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_4_3 = Station6_4_3; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_4_4 = Station6_4_4; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_4_5 = Station6_4_5; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_4_6 = Station6_4_6; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_4_7 = Station6_4_7; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_5_0 = Station6_5_0; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_5_1 = Station6_5_1; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_5_2 = Station6_5_2; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_5_3 = Station6_5_3; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_5_4 = Station6_5_4; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_5_5 = Station6_5_5; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_5_6 = Station6_5_6; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_5_7 = Station6_5_7; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_6_0 = Station6_6_0; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_6_1 = Station6_6_1; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_6_2 = Station6_6_2; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_6_3 = Station6_6_3; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_6_4 = Station6_6_4; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_6_5 = Station6_6_5; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_6_6 = Station6_6_6; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_6_7 = Station6_6_7; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_7_0 = Station6_7_0; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_7_1 = Station6_7_1; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_7_2 = Station6_7_2; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_7_3 = Station6_7_3; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_7_4 = Station6_7_4; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_7_5 = Station6_7_5; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_7_6 = Station6_7_6; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix6_7_7 = Station6_7_7; // @[stationary_dpe.scala 160:29]
  assign io_o_Stationary_matrix7_0_0 = Station7_0_0; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_0_1 = Station7_0_1; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_0_2 = Station7_0_2; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_0_3 = Station7_0_3; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_0_4 = Station7_0_4; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_0_5 = Station7_0_5; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_0_6 = Station7_0_6; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_0_7 = Station7_0_7; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_1_0 = Station7_1_0; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_1_1 = Station7_1_1; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_1_2 = Station7_1_2; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_1_3 = Station7_1_3; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_1_4 = Station7_1_4; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_1_5 = Station7_1_5; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_1_6 = Station7_1_6; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_1_7 = Station7_1_7; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_2_0 = Station7_2_0; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_2_1 = Station7_2_1; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_2_2 = Station7_2_2; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_2_3 = Station7_2_3; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_2_4 = Station7_2_4; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_2_5 = Station7_2_5; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_2_6 = Station7_2_6; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_2_7 = Station7_2_7; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_3_0 = Station7_3_0; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_3_1 = Station7_3_1; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_3_2 = Station7_3_2; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_3_3 = Station7_3_3; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_3_4 = Station7_3_4; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_3_5 = Station7_3_5; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_3_6 = Station7_3_6; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_3_7 = Station7_3_7; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_4_0 = Station7_4_0; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_4_1 = Station7_4_1; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_4_2 = Station7_4_2; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_4_3 = Station7_4_3; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_4_4 = Station7_4_4; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_4_5 = Station7_4_5; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_4_6 = Station7_4_6; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_4_7 = Station7_4_7; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_5_0 = Station7_5_0; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_5_1 = Station7_5_1; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_5_2 = Station7_5_2; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_5_3 = Station7_5_3; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_5_4 = Station7_5_4; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_5_5 = Station7_5_5; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_5_6 = Station7_5_6; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_5_7 = Station7_5_7; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_6_0 = Station7_6_0; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_6_1 = Station7_6_1; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_6_2 = Station7_6_2; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_6_3 = Station7_6_3; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_6_4 = Station7_6_4; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_6_5 = Station7_6_5; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_6_6 = Station7_6_6; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_6_7 = Station7_6_7; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_7_0 = Station7_7_0; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_7_1 = Station7_7_1; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_7_2 = Station7_7_2; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_7_3 = Station7_7_3; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_7_4 = Station7_7_4; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_7_5 = Station7_7_5; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_7_6 = Station7_7_6; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix7_7_7 = Station7_7_7; // @[stationary_dpe.scala 172:29]
  assign io_o_Stationary_matrix8_0_0 = Station8_0_0; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_0_1 = Station8_0_1; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_0_2 = Station8_0_2; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_0_3 = Station8_0_3; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_0_4 = Station8_0_4; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_0_5 = Station8_0_5; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_0_6 = Station8_0_6; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_0_7 = Station8_0_7; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_1_0 = Station8_1_0; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_1_1 = Station8_1_1; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_1_2 = Station8_1_2; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_1_3 = Station8_1_3; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_1_4 = Station8_1_4; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_1_5 = Station8_1_5; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_1_6 = Station8_1_6; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_1_7 = Station8_1_7; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_2_0 = Station8_2_0; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_2_1 = Station8_2_1; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_2_2 = Station8_2_2; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_2_3 = Station8_2_3; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_2_4 = Station8_2_4; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_2_5 = Station8_2_5; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_2_6 = Station8_2_6; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_2_7 = Station8_2_7; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_3_0 = Station8_3_0; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_3_1 = Station8_3_1; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_3_2 = Station8_3_2; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_3_3 = Station8_3_3; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_3_4 = Station8_3_4; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_3_5 = Station8_3_5; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_3_6 = Station8_3_6; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_3_7 = Station8_3_7; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_4_0 = Station8_4_0; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_4_1 = Station8_4_1; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_4_2 = Station8_4_2; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_4_3 = Station8_4_3; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_4_4 = Station8_4_4; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_4_5 = Station8_4_5; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_4_6 = Station8_4_6; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_4_7 = Station8_4_7; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_5_0 = Station8_5_0; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_5_1 = Station8_5_1; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_5_2 = Station8_5_2; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_5_3 = Station8_5_3; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_5_4 = Station8_5_4; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_5_5 = Station8_5_5; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_5_6 = Station8_5_6; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_5_7 = Station8_5_7; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_6_0 = Station8_6_0; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_6_1 = Station8_6_1; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_6_2 = Station8_6_2; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_6_3 = Station8_6_3; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_6_4 = Station8_6_4; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_6_5 = Station8_6_5; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_6_6 = Station8_6_6; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_6_7 = Station8_6_7; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_7_0 = Station8_7_0; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_7_1 = Station8_7_1; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_7_2 = Station8_7_2; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_7_3 = Station8_7_3; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_7_4 = Station8_7_4; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_7_5 = Station8_7_5; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_7_6 = Station8_7_6; // @[stationary_dpe.scala 184:29]
  assign io_o_Stationary_matrix8_7_7 = Station8_7_7; // @[stationary_dpe.scala 184:29]
  always @(posedge clock) begin
    if (reset) begin // @[stationary_dpe.scala 23:27]
      count <= 32'h0; // @[stationary_dpe.scala 23:27]
    end else if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        count <= _count_T_1; // @[stationary_dpe.scala 178:18]
      end else begin
        count <= _GEN_1995;
      end
    end else begin
      count <= _GEN_1995;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2264 & _GEN_2279) begin // @[stationary_dpe.scala 95:32]
          Station2_0_0 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_0_0 <= _GEN_0;
        end
      end else begin
        Station2_0_0 <= _GEN_0;
      end
    end else begin
      Station2_0_0 <= _GEN_0;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2264 & _GEN_2265) begin // @[stationary_dpe.scala 95:32]
          Station2_0_1 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_0_1 <= _GEN_1;
        end
      end else begin
        Station2_0_1 <= _GEN_1;
      end
    end else begin
      Station2_0_1 <= _GEN_1;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2264 & _GEN_2267) begin // @[stationary_dpe.scala 95:32]
          Station2_0_2 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_0_2 <= _GEN_2;
        end
      end else begin
        Station2_0_2 <= _GEN_2;
      end
    end else begin
      Station2_0_2 <= _GEN_2;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2264 & _GEN_2269) begin // @[stationary_dpe.scala 95:32]
          Station2_0_3 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_0_3 <= _GEN_3;
        end
      end else begin
        Station2_0_3 <= _GEN_3;
      end
    end else begin
      Station2_0_3 <= _GEN_3;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2264 & _GEN_2271) begin // @[stationary_dpe.scala 95:32]
          Station2_0_4 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_0_4 <= _GEN_4;
        end
      end else begin
        Station2_0_4 <= _GEN_4;
      end
    end else begin
      Station2_0_4 <= _GEN_4;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2264 & _GEN_2273) begin // @[stationary_dpe.scala 95:32]
          Station2_0_5 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_0_5 <= _GEN_5;
        end
      end else begin
        Station2_0_5 <= _GEN_5;
      end
    end else begin
      Station2_0_5 <= _GEN_5;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2264 & _GEN_2275) begin // @[stationary_dpe.scala 95:32]
          Station2_0_6 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_0_6 <= _GEN_6;
        end
      end else begin
        Station2_0_6 <= _GEN_6;
      end
    end else begin
      Station2_0_6 <= _GEN_6;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2264 & _GEN_2277) begin // @[stationary_dpe.scala 95:32]
          Station2_0_7 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_0_7 <= _GEN_7;
        end
      end else begin
        Station2_0_7 <= _GEN_7;
      end
    end else begin
      Station2_0_7 <= _GEN_7;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2278 & _GEN_2279) begin // @[stationary_dpe.scala 95:32]
          Station2_1_0 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_1_0 <= _GEN_8;
        end
      end else begin
        Station2_1_0 <= _GEN_8;
      end
    end else begin
      Station2_1_0 <= _GEN_8;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2278 & _GEN_2265) begin // @[stationary_dpe.scala 95:32]
          Station2_1_1 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_1_1 <= _GEN_9;
        end
      end else begin
        Station2_1_1 <= _GEN_9;
      end
    end else begin
      Station2_1_1 <= _GEN_9;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2278 & _GEN_2267) begin // @[stationary_dpe.scala 95:32]
          Station2_1_2 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_1_2 <= _GEN_10;
        end
      end else begin
        Station2_1_2 <= _GEN_10;
      end
    end else begin
      Station2_1_2 <= _GEN_10;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2278 & _GEN_2269) begin // @[stationary_dpe.scala 95:32]
          Station2_1_3 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_1_3 <= _GEN_11;
        end
      end else begin
        Station2_1_3 <= _GEN_11;
      end
    end else begin
      Station2_1_3 <= _GEN_11;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2278 & _GEN_2271) begin // @[stationary_dpe.scala 95:32]
          Station2_1_4 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_1_4 <= _GEN_12;
        end
      end else begin
        Station2_1_4 <= _GEN_12;
      end
    end else begin
      Station2_1_4 <= _GEN_12;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2278 & _GEN_2273) begin // @[stationary_dpe.scala 95:32]
          Station2_1_5 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_1_5 <= _GEN_13;
        end
      end else begin
        Station2_1_5 <= _GEN_13;
      end
    end else begin
      Station2_1_5 <= _GEN_13;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2278 & _GEN_2275) begin // @[stationary_dpe.scala 95:32]
          Station2_1_6 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_1_6 <= _GEN_14;
        end
      end else begin
        Station2_1_6 <= _GEN_14;
      end
    end else begin
      Station2_1_6 <= _GEN_14;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2278 & _GEN_2277) begin // @[stationary_dpe.scala 95:32]
          Station2_1_7 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_1_7 <= _GEN_15;
        end
      end else begin
        Station2_1_7 <= _GEN_15;
      end
    end else begin
      Station2_1_7 <= _GEN_15;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2294 & _GEN_2279) begin // @[stationary_dpe.scala 95:32]
          Station2_2_0 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_2_0 <= _GEN_16;
        end
      end else begin
        Station2_2_0 <= _GEN_16;
      end
    end else begin
      Station2_2_0 <= _GEN_16;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2294 & _GEN_2265) begin // @[stationary_dpe.scala 95:32]
          Station2_2_1 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_2_1 <= _GEN_17;
        end
      end else begin
        Station2_2_1 <= _GEN_17;
      end
    end else begin
      Station2_2_1 <= _GEN_17;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2294 & _GEN_2267) begin // @[stationary_dpe.scala 95:32]
          Station2_2_2 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_2_2 <= _GEN_18;
        end
      end else begin
        Station2_2_2 <= _GEN_18;
      end
    end else begin
      Station2_2_2 <= _GEN_18;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2294 & _GEN_2269) begin // @[stationary_dpe.scala 95:32]
          Station2_2_3 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_2_3 <= _GEN_19;
        end
      end else begin
        Station2_2_3 <= _GEN_19;
      end
    end else begin
      Station2_2_3 <= _GEN_19;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2294 & _GEN_2271) begin // @[stationary_dpe.scala 95:32]
          Station2_2_4 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_2_4 <= _GEN_20;
        end
      end else begin
        Station2_2_4 <= _GEN_20;
      end
    end else begin
      Station2_2_4 <= _GEN_20;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2294 & _GEN_2273) begin // @[stationary_dpe.scala 95:32]
          Station2_2_5 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_2_5 <= _GEN_21;
        end
      end else begin
        Station2_2_5 <= _GEN_21;
      end
    end else begin
      Station2_2_5 <= _GEN_21;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2294 & _GEN_2275) begin // @[stationary_dpe.scala 95:32]
          Station2_2_6 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_2_6 <= _GEN_22;
        end
      end else begin
        Station2_2_6 <= _GEN_22;
      end
    end else begin
      Station2_2_6 <= _GEN_22;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2294 & _GEN_2277) begin // @[stationary_dpe.scala 95:32]
          Station2_2_7 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_2_7 <= _GEN_23;
        end
      end else begin
        Station2_2_7 <= _GEN_23;
      end
    end else begin
      Station2_2_7 <= _GEN_23;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2310 & _GEN_2279) begin // @[stationary_dpe.scala 95:32]
          Station2_3_0 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_3_0 <= _GEN_24;
        end
      end else begin
        Station2_3_0 <= _GEN_24;
      end
    end else begin
      Station2_3_0 <= _GEN_24;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2310 & _GEN_2265) begin // @[stationary_dpe.scala 95:32]
          Station2_3_1 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_3_1 <= _GEN_25;
        end
      end else begin
        Station2_3_1 <= _GEN_25;
      end
    end else begin
      Station2_3_1 <= _GEN_25;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2310 & _GEN_2267) begin // @[stationary_dpe.scala 95:32]
          Station2_3_2 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_3_2 <= _GEN_26;
        end
      end else begin
        Station2_3_2 <= _GEN_26;
      end
    end else begin
      Station2_3_2 <= _GEN_26;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2310 & _GEN_2269) begin // @[stationary_dpe.scala 95:32]
          Station2_3_3 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_3_3 <= _GEN_27;
        end
      end else begin
        Station2_3_3 <= _GEN_27;
      end
    end else begin
      Station2_3_3 <= _GEN_27;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2310 & _GEN_2271) begin // @[stationary_dpe.scala 95:32]
          Station2_3_4 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_3_4 <= _GEN_28;
        end
      end else begin
        Station2_3_4 <= _GEN_28;
      end
    end else begin
      Station2_3_4 <= _GEN_28;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2310 & _GEN_2273) begin // @[stationary_dpe.scala 95:32]
          Station2_3_5 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_3_5 <= _GEN_29;
        end
      end else begin
        Station2_3_5 <= _GEN_29;
      end
    end else begin
      Station2_3_5 <= _GEN_29;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2310 & _GEN_2275) begin // @[stationary_dpe.scala 95:32]
          Station2_3_6 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_3_6 <= _GEN_30;
        end
      end else begin
        Station2_3_6 <= _GEN_30;
      end
    end else begin
      Station2_3_6 <= _GEN_30;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2310 & _GEN_2277) begin // @[stationary_dpe.scala 95:32]
          Station2_3_7 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_3_7 <= _GEN_31;
        end
      end else begin
        Station2_3_7 <= _GEN_31;
      end
    end else begin
      Station2_3_7 <= _GEN_31;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2326 & _GEN_2279) begin // @[stationary_dpe.scala 95:32]
          Station2_4_0 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_4_0 <= _GEN_32;
        end
      end else begin
        Station2_4_0 <= _GEN_32;
      end
    end else begin
      Station2_4_0 <= _GEN_32;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2326 & _GEN_2265) begin // @[stationary_dpe.scala 95:32]
          Station2_4_1 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_4_1 <= _GEN_33;
        end
      end else begin
        Station2_4_1 <= _GEN_33;
      end
    end else begin
      Station2_4_1 <= _GEN_33;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2326 & _GEN_2267) begin // @[stationary_dpe.scala 95:32]
          Station2_4_2 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_4_2 <= _GEN_34;
        end
      end else begin
        Station2_4_2 <= _GEN_34;
      end
    end else begin
      Station2_4_2 <= _GEN_34;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2326 & _GEN_2269) begin // @[stationary_dpe.scala 95:32]
          Station2_4_3 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_4_3 <= _GEN_35;
        end
      end else begin
        Station2_4_3 <= _GEN_35;
      end
    end else begin
      Station2_4_3 <= _GEN_35;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2326 & _GEN_2271) begin // @[stationary_dpe.scala 95:32]
          Station2_4_4 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_4_4 <= _GEN_36;
        end
      end else begin
        Station2_4_4 <= _GEN_36;
      end
    end else begin
      Station2_4_4 <= _GEN_36;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2326 & _GEN_2273) begin // @[stationary_dpe.scala 95:32]
          Station2_4_5 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_4_5 <= _GEN_37;
        end
      end else begin
        Station2_4_5 <= _GEN_37;
      end
    end else begin
      Station2_4_5 <= _GEN_37;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2326 & _GEN_2275) begin // @[stationary_dpe.scala 95:32]
          Station2_4_6 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_4_6 <= _GEN_38;
        end
      end else begin
        Station2_4_6 <= _GEN_38;
      end
    end else begin
      Station2_4_6 <= _GEN_38;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2326 & _GEN_2277) begin // @[stationary_dpe.scala 95:32]
          Station2_4_7 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_4_7 <= _GEN_39;
        end
      end else begin
        Station2_4_7 <= _GEN_39;
      end
    end else begin
      Station2_4_7 <= _GEN_39;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2342 & _GEN_2279) begin // @[stationary_dpe.scala 95:32]
          Station2_5_0 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_5_0 <= _GEN_40;
        end
      end else begin
        Station2_5_0 <= _GEN_40;
      end
    end else begin
      Station2_5_0 <= _GEN_40;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2342 & _GEN_2265) begin // @[stationary_dpe.scala 95:32]
          Station2_5_1 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_5_1 <= _GEN_41;
        end
      end else begin
        Station2_5_1 <= _GEN_41;
      end
    end else begin
      Station2_5_1 <= _GEN_41;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2342 & _GEN_2267) begin // @[stationary_dpe.scala 95:32]
          Station2_5_2 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_5_2 <= _GEN_42;
        end
      end else begin
        Station2_5_2 <= _GEN_42;
      end
    end else begin
      Station2_5_2 <= _GEN_42;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2342 & _GEN_2269) begin // @[stationary_dpe.scala 95:32]
          Station2_5_3 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_5_3 <= _GEN_43;
        end
      end else begin
        Station2_5_3 <= _GEN_43;
      end
    end else begin
      Station2_5_3 <= _GEN_43;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2342 & _GEN_2271) begin // @[stationary_dpe.scala 95:32]
          Station2_5_4 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_5_4 <= _GEN_44;
        end
      end else begin
        Station2_5_4 <= _GEN_44;
      end
    end else begin
      Station2_5_4 <= _GEN_44;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2342 & _GEN_2273) begin // @[stationary_dpe.scala 95:32]
          Station2_5_5 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_5_5 <= _GEN_45;
        end
      end else begin
        Station2_5_5 <= _GEN_45;
      end
    end else begin
      Station2_5_5 <= _GEN_45;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2342 & _GEN_2275) begin // @[stationary_dpe.scala 95:32]
          Station2_5_6 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_5_6 <= _GEN_46;
        end
      end else begin
        Station2_5_6 <= _GEN_46;
      end
    end else begin
      Station2_5_6 <= _GEN_46;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2342 & _GEN_2277) begin // @[stationary_dpe.scala 95:32]
          Station2_5_7 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_5_7 <= _GEN_47;
        end
      end else begin
        Station2_5_7 <= _GEN_47;
      end
    end else begin
      Station2_5_7 <= _GEN_47;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2358 & _GEN_2279) begin // @[stationary_dpe.scala 95:32]
          Station2_6_0 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_6_0 <= _GEN_48;
        end
      end else begin
        Station2_6_0 <= _GEN_48;
      end
    end else begin
      Station2_6_0 <= _GEN_48;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2358 & _GEN_2265) begin // @[stationary_dpe.scala 95:32]
          Station2_6_1 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_6_1 <= _GEN_49;
        end
      end else begin
        Station2_6_1 <= _GEN_49;
      end
    end else begin
      Station2_6_1 <= _GEN_49;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2358 & _GEN_2267) begin // @[stationary_dpe.scala 95:32]
          Station2_6_2 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_6_2 <= _GEN_50;
        end
      end else begin
        Station2_6_2 <= _GEN_50;
      end
    end else begin
      Station2_6_2 <= _GEN_50;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2358 & _GEN_2269) begin // @[stationary_dpe.scala 95:32]
          Station2_6_3 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_6_3 <= _GEN_51;
        end
      end else begin
        Station2_6_3 <= _GEN_51;
      end
    end else begin
      Station2_6_3 <= _GEN_51;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2358 & _GEN_2271) begin // @[stationary_dpe.scala 95:32]
          Station2_6_4 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_6_4 <= _GEN_52;
        end
      end else begin
        Station2_6_4 <= _GEN_52;
      end
    end else begin
      Station2_6_4 <= _GEN_52;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2358 & _GEN_2273) begin // @[stationary_dpe.scala 95:32]
          Station2_6_5 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_6_5 <= _GEN_53;
        end
      end else begin
        Station2_6_5 <= _GEN_53;
      end
    end else begin
      Station2_6_5 <= _GEN_53;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2358 & _GEN_2275) begin // @[stationary_dpe.scala 95:32]
          Station2_6_6 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_6_6 <= _GEN_54;
        end
      end else begin
        Station2_6_6 <= _GEN_54;
      end
    end else begin
      Station2_6_6 <= _GEN_54;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2358 & _GEN_2277) begin // @[stationary_dpe.scala 95:32]
          Station2_6_7 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_6_7 <= _GEN_55;
        end
      end else begin
        Station2_6_7 <= _GEN_55;
      end
    end else begin
      Station2_6_7 <= _GEN_55;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2374 & _GEN_2279) begin // @[stationary_dpe.scala 95:32]
          Station2_7_0 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_7_0 <= _GEN_56;
        end
      end else begin
        Station2_7_0 <= _GEN_56;
      end
    end else begin
      Station2_7_0 <= _GEN_56;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2374 & _GEN_2265) begin // @[stationary_dpe.scala 95:32]
          Station2_7_1 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_7_1 <= _GEN_57;
        end
      end else begin
        Station2_7_1 <= _GEN_57;
      end
    end else begin
      Station2_7_1 <= _GEN_57;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2374 & _GEN_2267) begin // @[stationary_dpe.scala 95:32]
          Station2_7_2 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_7_2 <= _GEN_58;
        end
      end else begin
        Station2_7_2 <= _GEN_58;
      end
    end else begin
      Station2_7_2 <= _GEN_58;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2374 & _GEN_2269) begin // @[stationary_dpe.scala 95:32]
          Station2_7_3 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_7_3 <= _GEN_59;
        end
      end else begin
        Station2_7_3 <= _GEN_59;
      end
    end else begin
      Station2_7_3 <= _GEN_59;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2374 & _GEN_2271) begin // @[stationary_dpe.scala 95:32]
          Station2_7_4 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_7_4 <= _GEN_60;
        end
      end else begin
        Station2_7_4 <= _GEN_60;
      end
    end else begin
      Station2_7_4 <= _GEN_60;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2374 & _GEN_2273) begin // @[stationary_dpe.scala 95:32]
          Station2_7_5 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_7_5 <= _GEN_61;
        end
      end else begin
        Station2_7_5 <= _GEN_61;
      end
    end else begin
      Station2_7_5 <= _GEN_61;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2374 & _GEN_2275) begin // @[stationary_dpe.scala 95:32]
          Station2_7_6 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_7_6 <= _GEN_62;
        end
      end else begin
        Station2_7_6 <= _GEN_62;
      end
    end else begin
      Station2_7_6 <= _GEN_62;
    end
    if (~valid) begin // @[stationary_dpe.scala 93:27]
      if (_GEN_511 != 16'h0) begin // @[stationary_dpe.scala 94:51]
        if (_GEN_2374 & _GEN_2277) begin // @[stationary_dpe.scala 95:32]
          Station2_7_7 <= 16'h0; // @[stationary_dpe.scala 95:32]
        end else begin
          Station2_7_7 <= _GEN_63;
        end
      end else begin
        Station2_7_7 <= _GEN_63;
      end
    end else begin
      Station2_7_7 <= _GEN_63;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2264 & _GEN_2279) begin // @[stationary_dpe.scala 116:32]
          Station3_0_0 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_0_0 <= _GEN_64;
        end
      end else begin
        Station3_0_0 <= _GEN_64;
      end
    end else begin
      Station3_0_0 <= _GEN_64;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2264 & _GEN_2265) begin // @[stationary_dpe.scala 116:32]
          Station3_0_1 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_0_1 <= _GEN_65;
        end
      end else begin
        Station3_0_1 <= _GEN_65;
      end
    end else begin
      Station3_0_1 <= _GEN_65;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2264 & _GEN_2267) begin // @[stationary_dpe.scala 116:32]
          Station3_0_2 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_0_2 <= _GEN_66;
        end
      end else begin
        Station3_0_2 <= _GEN_66;
      end
    end else begin
      Station3_0_2 <= _GEN_66;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2264 & _GEN_2269) begin // @[stationary_dpe.scala 116:32]
          Station3_0_3 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_0_3 <= _GEN_67;
        end
      end else begin
        Station3_0_3 <= _GEN_67;
      end
    end else begin
      Station3_0_3 <= _GEN_67;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2264 & _GEN_2271) begin // @[stationary_dpe.scala 116:32]
          Station3_0_4 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_0_4 <= _GEN_68;
        end
      end else begin
        Station3_0_4 <= _GEN_68;
      end
    end else begin
      Station3_0_4 <= _GEN_68;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2264 & _GEN_2273) begin // @[stationary_dpe.scala 116:32]
          Station3_0_5 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_0_5 <= _GEN_69;
        end
      end else begin
        Station3_0_5 <= _GEN_69;
      end
    end else begin
      Station3_0_5 <= _GEN_69;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2264 & _GEN_2275) begin // @[stationary_dpe.scala 116:32]
          Station3_0_6 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_0_6 <= _GEN_70;
        end
      end else begin
        Station3_0_6 <= _GEN_70;
      end
    end else begin
      Station3_0_6 <= _GEN_70;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2264 & _GEN_2277) begin // @[stationary_dpe.scala 116:32]
          Station3_0_7 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_0_7 <= _GEN_71;
        end
      end else begin
        Station3_0_7 <= _GEN_71;
      end
    end else begin
      Station3_0_7 <= _GEN_71;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2278 & _GEN_2279) begin // @[stationary_dpe.scala 116:32]
          Station3_1_0 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_1_0 <= _GEN_72;
        end
      end else begin
        Station3_1_0 <= _GEN_72;
      end
    end else begin
      Station3_1_0 <= _GEN_72;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2278 & _GEN_2265) begin // @[stationary_dpe.scala 116:32]
          Station3_1_1 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_1_1 <= _GEN_73;
        end
      end else begin
        Station3_1_1 <= _GEN_73;
      end
    end else begin
      Station3_1_1 <= _GEN_73;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2278 & _GEN_2267) begin // @[stationary_dpe.scala 116:32]
          Station3_1_2 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_1_2 <= _GEN_74;
        end
      end else begin
        Station3_1_2 <= _GEN_74;
      end
    end else begin
      Station3_1_2 <= _GEN_74;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2278 & _GEN_2269) begin // @[stationary_dpe.scala 116:32]
          Station3_1_3 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_1_3 <= _GEN_75;
        end
      end else begin
        Station3_1_3 <= _GEN_75;
      end
    end else begin
      Station3_1_3 <= _GEN_75;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2278 & _GEN_2271) begin // @[stationary_dpe.scala 116:32]
          Station3_1_4 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_1_4 <= _GEN_76;
        end
      end else begin
        Station3_1_4 <= _GEN_76;
      end
    end else begin
      Station3_1_4 <= _GEN_76;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2278 & _GEN_2273) begin // @[stationary_dpe.scala 116:32]
          Station3_1_5 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_1_5 <= _GEN_77;
        end
      end else begin
        Station3_1_5 <= _GEN_77;
      end
    end else begin
      Station3_1_5 <= _GEN_77;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2278 & _GEN_2275) begin // @[stationary_dpe.scala 116:32]
          Station3_1_6 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_1_6 <= _GEN_78;
        end
      end else begin
        Station3_1_6 <= _GEN_78;
      end
    end else begin
      Station3_1_6 <= _GEN_78;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2278 & _GEN_2277) begin // @[stationary_dpe.scala 116:32]
          Station3_1_7 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_1_7 <= _GEN_79;
        end
      end else begin
        Station3_1_7 <= _GEN_79;
      end
    end else begin
      Station3_1_7 <= _GEN_79;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2294 & _GEN_2279) begin // @[stationary_dpe.scala 116:32]
          Station3_2_0 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_2_0 <= _GEN_80;
        end
      end else begin
        Station3_2_0 <= _GEN_80;
      end
    end else begin
      Station3_2_0 <= _GEN_80;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2294 & _GEN_2265) begin // @[stationary_dpe.scala 116:32]
          Station3_2_1 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_2_1 <= _GEN_81;
        end
      end else begin
        Station3_2_1 <= _GEN_81;
      end
    end else begin
      Station3_2_1 <= _GEN_81;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2294 & _GEN_2267) begin // @[stationary_dpe.scala 116:32]
          Station3_2_2 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_2_2 <= _GEN_82;
        end
      end else begin
        Station3_2_2 <= _GEN_82;
      end
    end else begin
      Station3_2_2 <= _GEN_82;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2294 & _GEN_2269) begin // @[stationary_dpe.scala 116:32]
          Station3_2_3 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_2_3 <= _GEN_83;
        end
      end else begin
        Station3_2_3 <= _GEN_83;
      end
    end else begin
      Station3_2_3 <= _GEN_83;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2294 & _GEN_2271) begin // @[stationary_dpe.scala 116:32]
          Station3_2_4 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_2_4 <= _GEN_84;
        end
      end else begin
        Station3_2_4 <= _GEN_84;
      end
    end else begin
      Station3_2_4 <= _GEN_84;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2294 & _GEN_2273) begin // @[stationary_dpe.scala 116:32]
          Station3_2_5 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_2_5 <= _GEN_85;
        end
      end else begin
        Station3_2_5 <= _GEN_85;
      end
    end else begin
      Station3_2_5 <= _GEN_85;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2294 & _GEN_2275) begin // @[stationary_dpe.scala 116:32]
          Station3_2_6 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_2_6 <= _GEN_86;
        end
      end else begin
        Station3_2_6 <= _GEN_86;
      end
    end else begin
      Station3_2_6 <= _GEN_86;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2294 & _GEN_2277) begin // @[stationary_dpe.scala 116:32]
          Station3_2_7 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_2_7 <= _GEN_87;
        end
      end else begin
        Station3_2_7 <= _GEN_87;
      end
    end else begin
      Station3_2_7 <= _GEN_87;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2310 & _GEN_2279) begin // @[stationary_dpe.scala 116:32]
          Station3_3_0 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_3_0 <= _GEN_88;
        end
      end else begin
        Station3_3_0 <= _GEN_88;
      end
    end else begin
      Station3_3_0 <= _GEN_88;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2310 & _GEN_2265) begin // @[stationary_dpe.scala 116:32]
          Station3_3_1 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_3_1 <= _GEN_89;
        end
      end else begin
        Station3_3_1 <= _GEN_89;
      end
    end else begin
      Station3_3_1 <= _GEN_89;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2310 & _GEN_2267) begin // @[stationary_dpe.scala 116:32]
          Station3_3_2 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_3_2 <= _GEN_90;
        end
      end else begin
        Station3_3_2 <= _GEN_90;
      end
    end else begin
      Station3_3_2 <= _GEN_90;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2310 & _GEN_2269) begin // @[stationary_dpe.scala 116:32]
          Station3_3_3 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_3_3 <= _GEN_91;
        end
      end else begin
        Station3_3_3 <= _GEN_91;
      end
    end else begin
      Station3_3_3 <= _GEN_91;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2310 & _GEN_2271) begin // @[stationary_dpe.scala 116:32]
          Station3_3_4 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_3_4 <= _GEN_92;
        end
      end else begin
        Station3_3_4 <= _GEN_92;
      end
    end else begin
      Station3_3_4 <= _GEN_92;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2310 & _GEN_2273) begin // @[stationary_dpe.scala 116:32]
          Station3_3_5 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_3_5 <= _GEN_93;
        end
      end else begin
        Station3_3_5 <= _GEN_93;
      end
    end else begin
      Station3_3_5 <= _GEN_93;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2310 & _GEN_2275) begin // @[stationary_dpe.scala 116:32]
          Station3_3_6 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_3_6 <= _GEN_94;
        end
      end else begin
        Station3_3_6 <= _GEN_94;
      end
    end else begin
      Station3_3_6 <= _GEN_94;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2310 & _GEN_2277) begin // @[stationary_dpe.scala 116:32]
          Station3_3_7 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_3_7 <= _GEN_95;
        end
      end else begin
        Station3_3_7 <= _GEN_95;
      end
    end else begin
      Station3_3_7 <= _GEN_95;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2326 & _GEN_2279) begin // @[stationary_dpe.scala 116:32]
          Station3_4_0 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_4_0 <= _GEN_96;
        end
      end else begin
        Station3_4_0 <= _GEN_96;
      end
    end else begin
      Station3_4_0 <= _GEN_96;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2326 & _GEN_2265) begin // @[stationary_dpe.scala 116:32]
          Station3_4_1 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_4_1 <= _GEN_97;
        end
      end else begin
        Station3_4_1 <= _GEN_97;
      end
    end else begin
      Station3_4_1 <= _GEN_97;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2326 & _GEN_2267) begin // @[stationary_dpe.scala 116:32]
          Station3_4_2 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_4_2 <= _GEN_98;
        end
      end else begin
        Station3_4_2 <= _GEN_98;
      end
    end else begin
      Station3_4_2 <= _GEN_98;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2326 & _GEN_2269) begin // @[stationary_dpe.scala 116:32]
          Station3_4_3 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_4_3 <= _GEN_99;
        end
      end else begin
        Station3_4_3 <= _GEN_99;
      end
    end else begin
      Station3_4_3 <= _GEN_99;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2326 & _GEN_2271) begin // @[stationary_dpe.scala 116:32]
          Station3_4_4 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_4_4 <= _GEN_100;
        end
      end else begin
        Station3_4_4 <= _GEN_100;
      end
    end else begin
      Station3_4_4 <= _GEN_100;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2326 & _GEN_2273) begin // @[stationary_dpe.scala 116:32]
          Station3_4_5 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_4_5 <= _GEN_101;
        end
      end else begin
        Station3_4_5 <= _GEN_101;
      end
    end else begin
      Station3_4_5 <= _GEN_101;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2326 & _GEN_2275) begin // @[stationary_dpe.scala 116:32]
          Station3_4_6 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_4_6 <= _GEN_102;
        end
      end else begin
        Station3_4_6 <= _GEN_102;
      end
    end else begin
      Station3_4_6 <= _GEN_102;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2326 & _GEN_2277) begin // @[stationary_dpe.scala 116:32]
          Station3_4_7 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_4_7 <= _GEN_103;
        end
      end else begin
        Station3_4_7 <= _GEN_103;
      end
    end else begin
      Station3_4_7 <= _GEN_103;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2342 & _GEN_2279) begin // @[stationary_dpe.scala 116:32]
          Station3_5_0 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_5_0 <= _GEN_104;
        end
      end else begin
        Station3_5_0 <= _GEN_104;
      end
    end else begin
      Station3_5_0 <= _GEN_104;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2342 & _GEN_2265) begin // @[stationary_dpe.scala 116:32]
          Station3_5_1 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_5_1 <= _GEN_105;
        end
      end else begin
        Station3_5_1 <= _GEN_105;
      end
    end else begin
      Station3_5_1 <= _GEN_105;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2342 & _GEN_2267) begin // @[stationary_dpe.scala 116:32]
          Station3_5_2 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_5_2 <= _GEN_106;
        end
      end else begin
        Station3_5_2 <= _GEN_106;
      end
    end else begin
      Station3_5_2 <= _GEN_106;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2342 & _GEN_2269) begin // @[stationary_dpe.scala 116:32]
          Station3_5_3 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_5_3 <= _GEN_107;
        end
      end else begin
        Station3_5_3 <= _GEN_107;
      end
    end else begin
      Station3_5_3 <= _GEN_107;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2342 & _GEN_2271) begin // @[stationary_dpe.scala 116:32]
          Station3_5_4 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_5_4 <= _GEN_108;
        end
      end else begin
        Station3_5_4 <= _GEN_108;
      end
    end else begin
      Station3_5_4 <= _GEN_108;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2342 & _GEN_2273) begin // @[stationary_dpe.scala 116:32]
          Station3_5_5 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_5_5 <= _GEN_109;
        end
      end else begin
        Station3_5_5 <= _GEN_109;
      end
    end else begin
      Station3_5_5 <= _GEN_109;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2342 & _GEN_2275) begin // @[stationary_dpe.scala 116:32]
          Station3_5_6 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_5_6 <= _GEN_110;
        end
      end else begin
        Station3_5_6 <= _GEN_110;
      end
    end else begin
      Station3_5_6 <= _GEN_110;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2342 & _GEN_2277) begin // @[stationary_dpe.scala 116:32]
          Station3_5_7 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_5_7 <= _GEN_111;
        end
      end else begin
        Station3_5_7 <= _GEN_111;
      end
    end else begin
      Station3_5_7 <= _GEN_111;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2358 & _GEN_2279) begin // @[stationary_dpe.scala 116:32]
          Station3_6_0 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_6_0 <= _GEN_112;
        end
      end else begin
        Station3_6_0 <= _GEN_112;
      end
    end else begin
      Station3_6_0 <= _GEN_112;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2358 & _GEN_2265) begin // @[stationary_dpe.scala 116:32]
          Station3_6_1 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_6_1 <= _GEN_113;
        end
      end else begin
        Station3_6_1 <= _GEN_113;
      end
    end else begin
      Station3_6_1 <= _GEN_113;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2358 & _GEN_2267) begin // @[stationary_dpe.scala 116:32]
          Station3_6_2 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_6_2 <= _GEN_114;
        end
      end else begin
        Station3_6_2 <= _GEN_114;
      end
    end else begin
      Station3_6_2 <= _GEN_114;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2358 & _GEN_2269) begin // @[stationary_dpe.scala 116:32]
          Station3_6_3 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_6_3 <= _GEN_115;
        end
      end else begin
        Station3_6_3 <= _GEN_115;
      end
    end else begin
      Station3_6_3 <= _GEN_115;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2358 & _GEN_2271) begin // @[stationary_dpe.scala 116:32]
          Station3_6_4 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_6_4 <= _GEN_116;
        end
      end else begin
        Station3_6_4 <= _GEN_116;
      end
    end else begin
      Station3_6_4 <= _GEN_116;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2358 & _GEN_2273) begin // @[stationary_dpe.scala 116:32]
          Station3_6_5 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_6_5 <= _GEN_117;
        end
      end else begin
        Station3_6_5 <= _GEN_117;
      end
    end else begin
      Station3_6_5 <= _GEN_117;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2358 & _GEN_2275) begin // @[stationary_dpe.scala 116:32]
          Station3_6_6 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_6_6 <= _GEN_118;
        end
      end else begin
        Station3_6_6 <= _GEN_118;
      end
    end else begin
      Station3_6_6 <= _GEN_118;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2358 & _GEN_2277) begin // @[stationary_dpe.scala 116:32]
          Station3_6_7 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_6_7 <= _GEN_119;
        end
      end else begin
        Station3_6_7 <= _GEN_119;
      end
    end else begin
      Station3_6_7 <= _GEN_119;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2374 & _GEN_2279) begin // @[stationary_dpe.scala 116:32]
          Station3_7_0 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_7_0 <= _GEN_120;
        end
      end else begin
        Station3_7_0 <= _GEN_120;
      end
    end else begin
      Station3_7_0 <= _GEN_120;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2374 & _GEN_2265) begin // @[stationary_dpe.scala 116:32]
          Station3_7_1 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_7_1 <= _GEN_121;
        end
      end else begin
        Station3_7_1 <= _GEN_121;
      end
    end else begin
      Station3_7_1 <= _GEN_121;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2374 & _GEN_2267) begin // @[stationary_dpe.scala 116:32]
          Station3_7_2 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_7_2 <= _GEN_122;
        end
      end else begin
        Station3_7_2 <= _GEN_122;
      end
    end else begin
      Station3_7_2 <= _GEN_122;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2374 & _GEN_2269) begin // @[stationary_dpe.scala 116:32]
          Station3_7_3 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_7_3 <= _GEN_123;
        end
      end else begin
        Station3_7_3 <= _GEN_123;
      end
    end else begin
      Station3_7_3 <= _GEN_123;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2374 & _GEN_2271) begin // @[stationary_dpe.scala 116:32]
          Station3_7_4 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_7_4 <= _GEN_124;
        end
      end else begin
        Station3_7_4 <= _GEN_124;
      end
    end else begin
      Station3_7_4 <= _GEN_124;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2374 & _GEN_2273) begin // @[stationary_dpe.scala 116:32]
          Station3_7_5 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_7_5 <= _GEN_125;
        end
      end else begin
        Station3_7_5 <= _GEN_125;
      end
    end else begin
      Station3_7_5 <= _GEN_125;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2374 & _GEN_2275) begin // @[stationary_dpe.scala 116:32]
          Station3_7_6 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_7_6 <= _GEN_126;
        end
      end else begin
        Station3_7_6 <= _GEN_126;
      end
    end else begin
      Station3_7_6 <= _GEN_126;
    end
    if (~valid1) begin // @[stationary_dpe.scala 114:29]
      if (_GEN_769 != 16'h0) begin // @[stationary_dpe.scala 115:39]
        if (_GEN_2374 & _GEN_2277) begin // @[stationary_dpe.scala 116:32]
          Station3_7_7 <= 16'h0; // @[stationary_dpe.scala 116:32]
        end else begin
          Station3_7_7 <= _GEN_127;
        end
      end else begin
        Station3_7_7 <= _GEN_127;
      end
    end else begin
      Station3_7_7 <= _GEN_127;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2264 & _GEN_2279) begin // @[stationary_dpe.scala 128:32]
          Station4_0_0 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_0_0 <= _GEN_128;
        end
      end else begin
        Station4_0_0 <= _GEN_128;
      end
    end else begin
      Station4_0_0 <= _GEN_128;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2264 & _GEN_2265) begin // @[stationary_dpe.scala 128:32]
          Station4_0_1 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_0_1 <= _GEN_129;
        end
      end else begin
        Station4_0_1 <= _GEN_129;
      end
    end else begin
      Station4_0_1 <= _GEN_129;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2264 & _GEN_2267) begin // @[stationary_dpe.scala 128:32]
          Station4_0_2 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_0_2 <= _GEN_130;
        end
      end else begin
        Station4_0_2 <= _GEN_130;
      end
    end else begin
      Station4_0_2 <= _GEN_130;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2264 & _GEN_2269) begin // @[stationary_dpe.scala 128:32]
          Station4_0_3 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_0_3 <= _GEN_131;
        end
      end else begin
        Station4_0_3 <= _GEN_131;
      end
    end else begin
      Station4_0_3 <= _GEN_131;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2264 & _GEN_2271) begin // @[stationary_dpe.scala 128:32]
          Station4_0_4 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_0_4 <= _GEN_132;
        end
      end else begin
        Station4_0_4 <= _GEN_132;
      end
    end else begin
      Station4_0_4 <= _GEN_132;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2264 & _GEN_2273) begin // @[stationary_dpe.scala 128:32]
          Station4_0_5 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_0_5 <= _GEN_133;
        end
      end else begin
        Station4_0_5 <= _GEN_133;
      end
    end else begin
      Station4_0_5 <= _GEN_133;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2264 & _GEN_2275) begin // @[stationary_dpe.scala 128:32]
          Station4_0_6 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_0_6 <= _GEN_134;
        end
      end else begin
        Station4_0_6 <= _GEN_134;
      end
    end else begin
      Station4_0_6 <= _GEN_134;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2264 & _GEN_2277) begin // @[stationary_dpe.scala 128:32]
          Station4_0_7 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_0_7 <= _GEN_135;
        end
      end else begin
        Station4_0_7 <= _GEN_135;
      end
    end else begin
      Station4_0_7 <= _GEN_135;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2278 & _GEN_2279) begin // @[stationary_dpe.scala 128:32]
          Station4_1_0 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_1_0 <= _GEN_136;
        end
      end else begin
        Station4_1_0 <= _GEN_136;
      end
    end else begin
      Station4_1_0 <= _GEN_136;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2278 & _GEN_2265) begin // @[stationary_dpe.scala 128:32]
          Station4_1_1 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_1_1 <= _GEN_137;
        end
      end else begin
        Station4_1_1 <= _GEN_137;
      end
    end else begin
      Station4_1_1 <= _GEN_137;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2278 & _GEN_2267) begin // @[stationary_dpe.scala 128:32]
          Station4_1_2 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_1_2 <= _GEN_138;
        end
      end else begin
        Station4_1_2 <= _GEN_138;
      end
    end else begin
      Station4_1_2 <= _GEN_138;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2278 & _GEN_2269) begin // @[stationary_dpe.scala 128:32]
          Station4_1_3 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_1_3 <= _GEN_139;
        end
      end else begin
        Station4_1_3 <= _GEN_139;
      end
    end else begin
      Station4_1_3 <= _GEN_139;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2278 & _GEN_2271) begin // @[stationary_dpe.scala 128:32]
          Station4_1_4 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_1_4 <= _GEN_140;
        end
      end else begin
        Station4_1_4 <= _GEN_140;
      end
    end else begin
      Station4_1_4 <= _GEN_140;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2278 & _GEN_2273) begin // @[stationary_dpe.scala 128:32]
          Station4_1_5 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_1_5 <= _GEN_141;
        end
      end else begin
        Station4_1_5 <= _GEN_141;
      end
    end else begin
      Station4_1_5 <= _GEN_141;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2278 & _GEN_2275) begin // @[stationary_dpe.scala 128:32]
          Station4_1_6 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_1_6 <= _GEN_142;
        end
      end else begin
        Station4_1_6 <= _GEN_142;
      end
    end else begin
      Station4_1_6 <= _GEN_142;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2278 & _GEN_2277) begin // @[stationary_dpe.scala 128:32]
          Station4_1_7 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_1_7 <= _GEN_143;
        end
      end else begin
        Station4_1_7 <= _GEN_143;
      end
    end else begin
      Station4_1_7 <= _GEN_143;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2294 & _GEN_2279) begin // @[stationary_dpe.scala 128:32]
          Station4_2_0 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_2_0 <= _GEN_144;
        end
      end else begin
        Station4_2_0 <= _GEN_144;
      end
    end else begin
      Station4_2_0 <= _GEN_144;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2294 & _GEN_2265) begin // @[stationary_dpe.scala 128:32]
          Station4_2_1 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_2_1 <= _GEN_145;
        end
      end else begin
        Station4_2_1 <= _GEN_145;
      end
    end else begin
      Station4_2_1 <= _GEN_145;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2294 & _GEN_2267) begin // @[stationary_dpe.scala 128:32]
          Station4_2_2 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_2_2 <= _GEN_146;
        end
      end else begin
        Station4_2_2 <= _GEN_146;
      end
    end else begin
      Station4_2_2 <= _GEN_146;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2294 & _GEN_2269) begin // @[stationary_dpe.scala 128:32]
          Station4_2_3 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_2_3 <= _GEN_147;
        end
      end else begin
        Station4_2_3 <= _GEN_147;
      end
    end else begin
      Station4_2_3 <= _GEN_147;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2294 & _GEN_2271) begin // @[stationary_dpe.scala 128:32]
          Station4_2_4 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_2_4 <= _GEN_148;
        end
      end else begin
        Station4_2_4 <= _GEN_148;
      end
    end else begin
      Station4_2_4 <= _GEN_148;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2294 & _GEN_2273) begin // @[stationary_dpe.scala 128:32]
          Station4_2_5 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_2_5 <= _GEN_149;
        end
      end else begin
        Station4_2_5 <= _GEN_149;
      end
    end else begin
      Station4_2_5 <= _GEN_149;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2294 & _GEN_2275) begin // @[stationary_dpe.scala 128:32]
          Station4_2_6 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_2_6 <= _GEN_150;
        end
      end else begin
        Station4_2_6 <= _GEN_150;
      end
    end else begin
      Station4_2_6 <= _GEN_150;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2294 & _GEN_2277) begin // @[stationary_dpe.scala 128:32]
          Station4_2_7 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_2_7 <= _GEN_151;
        end
      end else begin
        Station4_2_7 <= _GEN_151;
      end
    end else begin
      Station4_2_7 <= _GEN_151;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2310 & _GEN_2279) begin // @[stationary_dpe.scala 128:32]
          Station4_3_0 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_3_0 <= _GEN_152;
        end
      end else begin
        Station4_3_0 <= _GEN_152;
      end
    end else begin
      Station4_3_0 <= _GEN_152;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2310 & _GEN_2265) begin // @[stationary_dpe.scala 128:32]
          Station4_3_1 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_3_1 <= _GEN_153;
        end
      end else begin
        Station4_3_1 <= _GEN_153;
      end
    end else begin
      Station4_3_1 <= _GEN_153;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2310 & _GEN_2267) begin // @[stationary_dpe.scala 128:32]
          Station4_3_2 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_3_2 <= _GEN_154;
        end
      end else begin
        Station4_3_2 <= _GEN_154;
      end
    end else begin
      Station4_3_2 <= _GEN_154;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2310 & _GEN_2269) begin // @[stationary_dpe.scala 128:32]
          Station4_3_3 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_3_3 <= _GEN_155;
        end
      end else begin
        Station4_3_3 <= _GEN_155;
      end
    end else begin
      Station4_3_3 <= _GEN_155;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2310 & _GEN_2271) begin // @[stationary_dpe.scala 128:32]
          Station4_3_4 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_3_4 <= _GEN_156;
        end
      end else begin
        Station4_3_4 <= _GEN_156;
      end
    end else begin
      Station4_3_4 <= _GEN_156;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2310 & _GEN_2273) begin // @[stationary_dpe.scala 128:32]
          Station4_3_5 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_3_5 <= _GEN_157;
        end
      end else begin
        Station4_3_5 <= _GEN_157;
      end
    end else begin
      Station4_3_5 <= _GEN_157;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2310 & _GEN_2275) begin // @[stationary_dpe.scala 128:32]
          Station4_3_6 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_3_6 <= _GEN_158;
        end
      end else begin
        Station4_3_6 <= _GEN_158;
      end
    end else begin
      Station4_3_6 <= _GEN_158;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2310 & _GEN_2277) begin // @[stationary_dpe.scala 128:32]
          Station4_3_7 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_3_7 <= _GEN_159;
        end
      end else begin
        Station4_3_7 <= _GEN_159;
      end
    end else begin
      Station4_3_7 <= _GEN_159;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2326 & _GEN_2279) begin // @[stationary_dpe.scala 128:32]
          Station4_4_0 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_4_0 <= _GEN_160;
        end
      end else begin
        Station4_4_0 <= _GEN_160;
      end
    end else begin
      Station4_4_0 <= _GEN_160;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2326 & _GEN_2265) begin // @[stationary_dpe.scala 128:32]
          Station4_4_1 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_4_1 <= _GEN_161;
        end
      end else begin
        Station4_4_1 <= _GEN_161;
      end
    end else begin
      Station4_4_1 <= _GEN_161;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2326 & _GEN_2267) begin // @[stationary_dpe.scala 128:32]
          Station4_4_2 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_4_2 <= _GEN_162;
        end
      end else begin
        Station4_4_2 <= _GEN_162;
      end
    end else begin
      Station4_4_2 <= _GEN_162;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2326 & _GEN_2269) begin // @[stationary_dpe.scala 128:32]
          Station4_4_3 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_4_3 <= _GEN_163;
        end
      end else begin
        Station4_4_3 <= _GEN_163;
      end
    end else begin
      Station4_4_3 <= _GEN_163;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2326 & _GEN_2271) begin // @[stationary_dpe.scala 128:32]
          Station4_4_4 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_4_4 <= _GEN_164;
        end
      end else begin
        Station4_4_4 <= _GEN_164;
      end
    end else begin
      Station4_4_4 <= _GEN_164;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2326 & _GEN_2273) begin // @[stationary_dpe.scala 128:32]
          Station4_4_5 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_4_5 <= _GEN_165;
        end
      end else begin
        Station4_4_5 <= _GEN_165;
      end
    end else begin
      Station4_4_5 <= _GEN_165;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2326 & _GEN_2275) begin // @[stationary_dpe.scala 128:32]
          Station4_4_6 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_4_6 <= _GEN_166;
        end
      end else begin
        Station4_4_6 <= _GEN_166;
      end
    end else begin
      Station4_4_6 <= _GEN_166;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2326 & _GEN_2277) begin // @[stationary_dpe.scala 128:32]
          Station4_4_7 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_4_7 <= _GEN_167;
        end
      end else begin
        Station4_4_7 <= _GEN_167;
      end
    end else begin
      Station4_4_7 <= _GEN_167;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2342 & _GEN_2279) begin // @[stationary_dpe.scala 128:32]
          Station4_5_0 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_5_0 <= _GEN_168;
        end
      end else begin
        Station4_5_0 <= _GEN_168;
      end
    end else begin
      Station4_5_0 <= _GEN_168;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2342 & _GEN_2265) begin // @[stationary_dpe.scala 128:32]
          Station4_5_1 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_5_1 <= _GEN_169;
        end
      end else begin
        Station4_5_1 <= _GEN_169;
      end
    end else begin
      Station4_5_1 <= _GEN_169;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2342 & _GEN_2267) begin // @[stationary_dpe.scala 128:32]
          Station4_5_2 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_5_2 <= _GEN_170;
        end
      end else begin
        Station4_5_2 <= _GEN_170;
      end
    end else begin
      Station4_5_2 <= _GEN_170;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2342 & _GEN_2269) begin // @[stationary_dpe.scala 128:32]
          Station4_5_3 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_5_3 <= _GEN_171;
        end
      end else begin
        Station4_5_3 <= _GEN_171;
      end
    end else begin
      Station4_5_3 <= _GEN_171;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2342 & _GEN_2271) begin // @[stationary_dpe.scala 128:32]
          Station4_5_4 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_5_4 <= _GEN_172;
        end
      end else begin
        Station4_5_4 <= _GEN_172;
      end
    end else begin
      Station4_5_4 <= _GEN_172;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2342 & _GEN_2273) begin // @[stationary_dpe.scala 128:32]
          Station4_5_5 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_5_5 <= _GEN_173;
        end
      end else begin
        Station4_5_5 <= _GEN_173;
      end
    end else begin
      Station4_5_5 <= _GEN_173;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2342 & _GEN_2275) begin // @[stationary_dpe.scala 128:32]
          Station4_5_6 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_5_6 <= _GEN_174;
        end
      end else begin
        Station4_5_6 <= _GEN_174;
      end
    end else begin
      Station4_5_6 <= _GEN_174;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2342 & _GEN_2277) begin // @[stationary_dpe.scala 128:32]
          Station4_5_7 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_5_7 <= _GEN_175;
        end
      end else begin
        Station4_5_7 <= _GEN_175;
      end
    end else begin
      Station4_5_7 <= _GEN_175;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2358 & _GEN_2279) begin // @[stationary_dpe.scala 128:32]
          Station4_6_0 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_6_0 <= _GEN_176;
        end
      end else begin
        Station4_6_0 <= _GEN_176;
      end
    end else begin
      Station4_6_0 <= _GEN_176;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2358 & _GEN_2265) begin // @[stationary_dpe.scala 128:32]
          Station4_6_1 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_6_1 <= _GEN_177;
        end
      end else begin
        Station4_6_1 <= _GEN_177;
      end
    end else begin
      Station4_6_1 <= _GEN_177;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2358 & _GEN_2267) begin // @[stationary_dpe.scala 128:32]
          Station4_6_2 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_6_2 <= _GEN_178;
        end
      end else begin
        Station4_6_2 <= _GEN_178;
      end
    end else begin
      Station4_6_2 <= _GEN_178;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2358 & _GEN_2269) begin // @[stationary_dpe.scala 128:32]
          Station4_6_3 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_6_3 <= _GEN_179;
        end
      end else begin
        Station4_6_3 <= _GEN_179;
      end
    end else begin
      Station4_6_3 <= _GEN_179;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2358 & _GEN_2271) begin // @[stationary_dpe.scala 128:32]
          Station4_6_4 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_6_4 <= _GEN_180;
        end
      end else begin
        Station4_6_4 <= _GEN_180;
      end
    end else begin
      Station4_6_4 <= _GEN_180;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2358 & _GEN_2273) begin // @[stationary_dpe.scala 128:32]
          Station4_6_5 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_6_5 <= _GEN_181;
        end
      end else begin
        Station4_6_5 <= _GEN_181;
      end
    end else begin
      Station4_6_5 <= _GEN_181;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2358 & _GEN_2275) begin // @[stationary_dpe.scala 128:32]
          Station4_6_6 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_6_6 <= _GEN_182;
        end
      end else begin
        Station4_6_6 <= _GEN_182;
      end
    end else begin
      Station4_6_6 <= _GEN_182;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2358 & _GEN_2277) begin // @[stationary_dpe.scala 128:32]
          Station4_6_7 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_6_7 <= _GEN_183;
        end
      end else begin
        Station4_6_7 <= _GEN_183;
      end
    end else begin
      Station4_6_7 <= _GEN_183;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2374 & _GEN_2279) begin // @[stationary_dpe.scala 128:32]
          Station4_7_0 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_7_0 <= _GEN_184;
        end
      end else begin
        Station4_7_0 <= _GEN_184;
      end
    end else begin
      Station4_7_0 <= _GEN_184;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2374 & _GEN_2265) begin // @[stationary_dpe.scala 128:32]
          Station4_7_1 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_7_1 <= _GEN_185;
        end
      end else begin
        Station4_7_1 <= _GEN_185;
      end
    end else begin
      Station4_7_1 <= _GEN_185;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2374 & _GEN_2267) begin // @[stationary_dpe.scala 128:32]
          Station4_7_2 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_7_2 <= _GEN_186;
        end
      end else begin
        Station4_7_2 <= _GEN_186;
      end
    end else begin
      Station4_7_2 <= _GEN_186;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2374 & _GEN_2269) begin // @[stationary_dpe.scala 128:32]
          Station4_7_3 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_7_3 <= _GEN_187;
        end
      end else begin
        Station4_7_3 <= _GEN_187;
      end
    end else begin
      Station4_7_3 <= _GEN_187;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2374 & _GEN_2271) begin // @[stationary_dpe.scala 128:32]
          Station4_7_4 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_7_4 <= _GEN_188;
        end
      end else begin
        Station4_7_4 <= _GEN_188;
      end
    end else begin
      Station4_7_4 <= _GEN_188;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2374 & _GEN_2273) begin // @[stationary_dpe.scala 128:32]
          Station4_7_5 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_7_5 <= _GEN_189;
        end
      end else begin
        Station4_7_5 <= _GEN_189;
      end
    end else begin
      Station4_7_5 <= _GEN_189;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2374 & _GEN_2275) begin // @[stationary_dpe.scala 128:32]
          Station4_7_6 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_7_6 <= _GEN_190;
        end
      end else begin
        Station4_7_6 <= _GEN_190;
      end
    end else begin
      Station4_7_6 <= _GEN_190;
    end
    if (~valid2) begin // @[stationary_dpe.scala 126:29]
      if (_GEN_1027 != 16'h0) begin // @[stationary_dpe.scala 127:39]
        if (_GEN_2374 & _GEN_2277) begin // @[stationary_dpe.scala 128:32]
          Station4_7_7 <= 16'h0; // @[stationary_dpe.scala 128:32]
        end else begin
          Station4_7_7 <= _GEN_191;
        end
      end else begin
        Station4_7_7 <= _GEN_191;
      end
    end else begin
      Station4_7_7 <= _GEN_191;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2264 & _GEN_2279) begin // @[stationary_dpe.scala 140:32]
          Station5_0_0 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_0_0 <= _GEN_192;
        end
      end else begin
        Station5_0_0 <= _GEN_192;
      end
    end else begin
      Station5_0_0 <= _GEN_192;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2264 & _GEN_2265) begin // @[stationary_dpe.scala 140:32]
          Station5_0_1 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_0_1 <= _GEN_193;
        end
      end else begin
        Station5_0_1 <= _GEN_193;
      end
    end else begin
      Station5_0_1 <= _GEN_193;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2264 & _GEN_2267) begin // @[stationary_dpe.scala 140:32]
          Station5_0_2 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_0_2 <= _GEN_194;
        end
      end else begin
        Station5_0_2 <= _GEN_194;
      end
    end else begin
      Station5_0_2 <= _GEN_194;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2264 & _GEN_2269) begin // @[stationary_dpe.scala 140:32]
          Station5_0_3 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_0_3 <= _GEN_195;
        end
      end else begin
        Station5_0_3 <= _GEN_195;
      end
    end else begin
      Station5_0_3 <= _GEN_195;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2264 & _GEN_2271) begin // @[stationary_dpe.scala 140:32]
          Station5_0_4 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_0_4 <= _GEN_196;
        end
      end else begin
        Station5_0_4 <= _GEN_196;
      end
    end else begin
      Station5_0_4 <= _GEN_196;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2264 & _GEN_2273) begin // @[stationary_dpe.scala 140:32]
          Station5_0_5 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_0_5 <= _GEN_197;
        end
      end else begin
        Station5_0_5 <= _GEN_197;
      end
    end else begin
      Station5_0_5 <= _GEN_197;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2264 & _GEN_2275) begin // @[stationary_dpe.scala 140:32]
          Station5_0_6 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_0_6 <= _GEN_198;
        end
      end else begin
        Station5_0_6 <= _GEN_198;
      end
    end else begin
      Station5_0_6 <= _GEN_198;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2264 & _GEN_2277) begin // @[stationary_dpe.scala 140:32]
          Station5_0_7 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_0_7 <= _GEN_199;
        end
      end else begin
        Station5_0_7 <= _GEN_199;
      end
    end else begin
      Station5_0_7 <= _GEN_199;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2278 & _GEN_2279) begin // @[stationary_dpe.scala 140:32]
          Station5_1_0 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_1_0 <= _GEN_200;
        end
      end else begin
        Station5_1_0 <= _GEN_200;
      end
    end else begin
      Station5_1_0 <= _GEN_200;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2278 & _GEN_2265) begin // @[stationary_dpe.scala 140:32]
          Station5_1_1 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_1_1 <= _GEN_201;
        end
      end else begin
        Station5_1_1 <= _GEN_201;
      end
    end else begin
      Station5_1_1 <= _GEN_201;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2278 & _GEN_2267) begin // @[stationary_dpe.scala 140:32]
          Station5_1_2 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_1_2 <= _GEN_202;
        end
      end else begin
        Station5_1_2 <= _GEN_202;
      end
    end else begin
      Station5_1_2 <= _GEN_202;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2278 & _GEN_2269) begin // @[stationary_dpe.scala 140:32]
          Station5_1_3 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_1_3 <= _GEN_203;
        end
      end else begin
        Station5_1_3 <= _GEN_203;
      end
    end else begin
      Station5_1_3 <= _GEN_203;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2278 & _GEN_2271) begin // @[stationary_dpe.scala 140:32]
          Station5_1_4 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_1_4 <= _GEN_204;
        end
      end else begin
        Station5_1_4 <= _GEN_204;
      end
    end else begin
      Station5_1_4 <= _GEN_204;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2278 & _GEN_2273) begin // @[stationary_dpe.scala 140:32]
          Station5_1_5 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_1_5 <= _GEN_205;
        end
      end else begin
        Station5_1_5 <= _GEN_205;
      end
    end else begin
      Station5_1_5 <= _GEN_205;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2278 & _GEN_2275) begin // @[stationary_dpe.scala 140:32]
          Station5_1_6 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_1_6 <= _GEN_206;
        end
      end else begin
        Station5_1_6 <= _GEN_206;
      end
    end else begin
      Station5_1_6 <= _GEN_206;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2278 & _GEN_2277) begin // @[stationary_dpe.scala 140:32]
          Station5_1_7 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_1_7 <= _GEN_207;
        end
      end else begin
        Station5_1_7 <= _GEN_207;
      end
    end else begin
      Station5_1_7 <= _GEN_207;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2294 & _GEN_2279) begin // @[stationary_dpe.scala 140:32]
          Station5_2_0 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_2_0 <= _GEN_208;
        end
      end else begin
        Station5_2_0 <= _GEN_208;
      end
    end else begin
      Station5_2_0 <= _GEN_208;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2294 & _GEN_2265) begin // @[stationary_dpe.scala 140:32]
          Station5_2_1 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_2_1 <= _GEN_209;
        end
      end else begin
        Station5_2_1 <= _GEN_209;
      end
    end else begin
      Station5_2_1 <= _GEN_209;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2294 & _GEN_2267) begin // @[stationary_dpe.scala 140:32]
          Station5_2_2 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_2_2 <= _GEN_210;
        end
      end else begin
        Station5_2_2 <= _GEN_210;
      end
    end else begin
      Station5_2_2 <= _GEN_210;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2294 & _GEN_2269) begin // @[stationary_dpe.scala 140:32]
          Station5_2_3 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_2_3 <= _GEN_211;
        end
      end else begin
        Station5_2_3 <= _GEN_211;
      end
    end else begin
      Station5_2_3 <= _GEN_211;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2294 & _GEN_2271) begin // @[stationary_dpe.scala 140:32]
          Station5_2_4 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_2_4 <= _GEN_212;
        end
      end else begin
        Station5_2_4 <= _GEN_212;
      end
    end else begin
      Station5_2_4 <= _GEN_212;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2294 & _GEN_2273) begin // @[stationary_dpe.scala 140:32]
          Station5_2_5 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_2_5 <= _GEN_213;
        end
      end else begin
        Station5_2_5 <= _GEN_213;
      end
    end else begin
      Station5_2_5 <= _GEN_213;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2294 & _GEN_2275) begin // @[stationary_dpe.scala 140:32]
          Station5_2_6 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_2_6 <= _GEN_214;
        end
      end else begin
        Station5_2_6 <= _GEN_214;
      end
    end else begin
      Station5_2_6 <= _GEN_214;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2294 & _GEN_2277) begin // @[stationary_dpe.scala 140:32]
          Station5_2_7 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_2_7 <= _GEN_215;
        end
      end else begin
        Station5_2_7 <= _GEN_215;
      end
    end else begin
      Station5_2_7 <= _GEN_215;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2310 & _GEN_2279) begin // @[stationary_dpe.scala 140:32]
          Station5_3_0 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_3_0 <= _GEN_216;
        end
      end else begin
        Station5_3_0 <= _GEN_216;
      end
    end else begin
      Station5_3_0 <= _GEN_216;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2310 & _GEN_2265) begin // @[stationary_dpe.scala 140:32]
          Station5_3_1 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_3_1 <= _GEN_217;
        end
      end else begin
        Station5_3_1 <= _GEN_217;
      end
    end else begin
      Station5_3_1 <= _GEN_217;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2310 & _GEN_2267) begin // @[stationary_dpe.scala 140:32]
          Station5_3_2 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_3_2 <= _GEN_218;
        end
      end else begin
        Station5_3_2 <= _GEN_218;
      end
    end else begin
      Station5_3_2 <= _GEN_218;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2310 & _GEN_2269) begin // @[stationary_dpe.scala 140:32]
          Station5_3_3 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_3_3 <= _GEN_219;
        end
      end else begin
        Station5_3_3 <= _GEN_219;
      end
    end else begin
      Station5_3_3 <= _GEN_219;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2310 & _GEN_2271) begin // @[stationary_dpe.scala 140:32]
          Station5_3_4 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_3_4 <= _GEN_220;
        end
      end else begin
        Station5_3_4 <= _GEN_220;
      end
    end else begin
      Station5_3_4 <= _GEN_220;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2310 & _GEN_2273) begin // @[stationary_dpe.scala 140:32]
          Station5_3_5 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_3_5 <= _GEN_221;
        end
      end else begin
        Station5_3_5 <= _GEN_221;
      end
    end else begin
      Station5_3_5 <= _GEN_221;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2310 & _GEN_2275) begin // @[stationary_dpe.scala 140:32]
          Station5_3_6 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_3_6 <= _GEN_222;
        end
      end else begin
        Station5_3_6 <= _GEN_222;
      end
    end else begin
      Station5_3_6 <= _GEN_222;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2310 & _GEN_2277) begin // @[stationary_dpe.scala 140:32]
          Station5_3_7 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_3_7 <= _GEN_223;
        end
      end else begin
        Station5_3_7 <= _GEN_223;
      end
    end else begin
      Station5_3_7 <= _GEN_223;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2326 & _GEN_2279) begin // @[stationary_dpe.scala 140:32]
          Station5_4_0 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_4_0 <= _GEN_224;
        end
      end else begin
        Station5_4_0 <= _GEN_224;
      end
    end else begin
      Station5_4_0 <= _GEN_224;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2326 & _GEN_2265) begin // @[stationary_dpe.scala 140:32]
          Station5_4_1 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_4_1 <= _GEN_225;
        end
      end else begin
        Station5_4_1 <= _GEN_225;
      end
    end else begin
      Station5_4_1 <= _GEN_225;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2326 & _GEN_2267) begin // @[stationary_dpe.scala 140:32]
          Station5_4_2 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_4_2 <= _GEN_226;
        end
      end else begin
        Station5_4_2 <= _GEN_226;
      end
    end else begin
      Station5_4_2 <= _GEN_226;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2326 & _GEN_2269) begin // @[stationary_dpe.scala 140:32]
          Station5_4_3 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_4_3 <= _GEN_227;
        end
      end else begin
        Station5_4_3 <= _GEN_227;
      end
    end else begin
      Station5_4_3 <= _GEN_227;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2326 & _GEN_2271) begin // @[stationary_dpe.scala 140:32]
          Station5_4_4 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_4_4 <= _GEN_228;
        end
      end else begin
        Station5_4_4 <= _GEN_228;
      end
    end else begin
      Station5_4_4 <= _GEN_228;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2326 & _GEN_2273) begin // @[stationary_dpe.scala 140:32]
          Station5_4_5 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_4_5 <= _GEN_229;
        end
      end else begin
        Station5_4_5 <= _GEN_229;
      end
    end else begin
      Station5_4_5 <= _GEN_229;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2326 & _GEN_2275) begin // @[stationary_dpe.scala 140:32]
          Station5_4_6 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_4_6 <= _GEN_230;
        end
      end else begin
        Station5_4_6 <= _GEN_230;
      end
    end else begin
      Station5_4_6 <= _GEN_230;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2326 & _GEN_2277) begin // @[stationary_dpe.scala 140:32]
          Station5_4_7 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_4_7 <= _GEN_231;
        end
      end else begin
        Station5_4_7 <= _GEN_231;
      end
    end else begin
      Station5_4_7 <= _GEN_231;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2342 & _GEN_2279) begin // @[stationary_dpe.scala 140:32]
          Station5_5_0 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_5_0 <= _GEN_232;
        end
      end else begin
        Station5_5_0 <= _GEN_232;
      end
    end else begin
      Station5_5_0 <= _GEN_232;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2342 & _GEN_2265) begin // @[stationary_dpe.scala 140:32]
          Station5_5_1 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_5_1 <= _GEN_233;
        end
      end else begin
        Station5_5_1 <= _GEN_233;
      end
    end else begin
      Station5_5_1 <= _GEN_233;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2342 & _GEN_2267) begin // @[stationary_dpe.scala 140:32]
          Station5_5_2 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_5_2 <= _GEN_234;
        end
      end else begin
        Station5_5_2 <= _GEN_234;
      end
    end else begin
      Station5_5_2 <= _GEN_234;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2342 & _GEN_2269) begin // @[stationary_dpe.scala 140:32]
          Station5_5_3 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_5_3 <= _GEN_235;
        end
      end else begin
        Station5_5_3 <= _GEN_235;
      end
    end else begin
      Station5_5_3 <= _GEN_235;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2342 & _GEN_2271) begin // @[stationary_dpe.scala 140:32]
          Station5_5_4 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_5_4 <= _GEN_236;
        end
      end else begin
        Station5_5_4 <= _GEN_236;
      end
    end else begin
      Station5_5_4 <= _GEN_236;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2342 & _GEN_2273) begin // @[stationary_dpe.scala 140:32]
          Station5_5_5 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_5_5 <= _GEN_237;
        end
      end else begin
        Station5_5_5 <= _GEN_237;
      end
    end else begin
      Station5_5_5 <= _GEN_237;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2342 & _GEN_2275) begin // @[stationary_dpe.scala 140:32]
          Station5_5_6 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_5_6 <= _GEN_238;
        end
      end else begin
        Station5_5_6 <= _GEN_238;
      end
    end else begin
      Station5_5_6 <= _GEN_238;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2342 & _GEN_2277) begin // @[stationary_dpe.scala 140:32]
          Station5_5_7 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_5_7 <= _GEN_239;
        end
      end else begin
        Station5_5_7 <= _GEN_239;
      end
    end else begin
      Station5_5_7 <= _GEN_239;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2358 & _GEN_2279) begin // @[stationary_dpe.scala 140:32]
          Station5_6_0 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_6_0 <= _GEN_240;
        end
      end else begin
        Station5_6_0 <= _GEN_240;
      end
    end else begin
      Station5_6_0 <= _GEN_240;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2358 & _GEN_2265) begin // @[stationary_dpe.scala 140:32]
          Station5_6_1 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_6_1 <= _GEN_241;
        end
      end else begin
        Station5_6_1 <= _GEN_241;
      end
    end else begin
      Station5_6_1 <= _GEN_241;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2358 & _GEN_2267) begin // @[stationary_dpe.scala 140:32]
          Station5_6_2 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_6_2 <= _GEN_242;
        end
      end else begin
        Station5_6_2 <= _GEN_242;
      end
    end else begin
      Station5_6_2 <= _GEN_242;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2358 & _GEN_2269) begin // @[stationary_dpe.scala 140:32]
          Station5_6_3 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_6_3 <= _GEN_243;
        end
      end else begin
        Station5_6_3 <= _GEN_243;
      end
    end else begin
      Station5_6_3 <= _GEN_243;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2358 & _GEN_2271) begin // @[stationary_dpe.scala 140:32]
          Station5_6_4 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_6_4 <= _GEN_244;
        end
      end else begin
        Station5_6_4 <= _GEN_244;
      end
    end else begin
      Station5_6_4 <= _GEN_244;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2358 & _GEN_2273) begin // @[stationary_dpe.scala 140:32]
          Station5_6_5 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_6_5 <= _GEN_245;
        end
      end else begin
        Station5_6_5 <= _GEN_245;
      end
    end else begin
      Station5_6_5 <= _GEN_245;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2358 & _GEN_2275) begin // @[stationary_dpe.scala 140:32]
          Station5_6_6 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_6_6 <= _GEN_246;
        end
      end else begin
        Station5_6_6 <= _GEN_246;
      end
    end else begin
      Station5_6_6 <= _GEN_246;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2358 & _GEN_2277) begin // @[stationary_dpe.scala 140:32]
          Station5_6_7 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_6_7 <= _GEN_247;
        end
      end else begin
        Station5_6_7 <= _GEN_247;
      end
    end else begin
      Station5_6_7 <= _GEN_247;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2374 & _GEN_2279) begin // @[stationary_dpe.scala 140:32]
          Station5_7_0 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_7_0 <= _GEN_248;
        end
      end else begin
        Station5_7_0 <= _GEN_248;
      end
    end else begin
      Station5_7_0 <= _GEN_248;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2374 & _GEN_2265) begin // @[stationary_dpe.scala 140:32]
          Station5_7_1 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_7_1 <= _GEN_249;
        end
      end else begin
        Station5_7_1 <= _GEN_249;
      end
    end else begin
      Station5_7_1 <= _GEN_249;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2374 & _GEN_2267) begin // @[stationary_dpe.scala 140:32]
          Station5_7_2 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_7_2 <= _GEN_250;
        end
      end else begin
        Station5_7_2 <= _GEN_250;
      end
    end else begin
      Station5_7_2 <= _GEN_250;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2374 & _GEN_2269) begin // @[stationary_dpe.scala 140:32]
          Station5_7_3 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_7_3 <= _GEN_251;
        end
      end else begin
        Station5_7_3 <= _GEN_251;
      end
    end else begin
      Station5_7_3 <= _GEN_251;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2374 & _GEN_2271) begin // @[stationary_dpe.scala 140:32]
          Station5_7_4 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_7_4 <= _GEN_252;
        end
      end else begin
        Station5_7_4 <= _GEN_252;
      end
    end else begin
      Station5_7_4 <= _GEN_252;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2374 & _GEN_2273) begin // @[stationary_dpe.scala 140:32]
          Station5_7_5 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_7_5 <= _GEN_253;
        end
      end else begin
        Station5_7_5 <= _GEN_253;
      end
    end else begin
      Station5_7_5 <= _GEN_253;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2374 & _GEN_2275) begin // @[stationary_dpe.scala 140:32]
          Station5_7_6 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_7_6 <= _GEN_254;
        end
      end else begin
        Station5_7_6 <= _GEN_254;
      end
    end else begin
      Station5_7_6 <= _GEN_254;
    end
    if (~valid3) begin // @[stationary_dpe.scala 138:28]
      if (_GEN_1285 != 16'h0) begin // @[stationary_dpe.scala 139:39]
        if (_GEN_2374 & _GEN_2277) begin // @[stationary_dpe.scala 140:32]
          Station5_7_7 <= 16'h0; // @[stationary_dpe.scala 140:32]
        end else begin
          Station5_7_7 <= _GEN_255;
        end
      end else begin
        Station5_7_7 <= _GEN_255;
      end
    end else begin
      Station5_7_7 <= _GEN_255;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2264 & _GEN_2279) begin // @[stationary_dpe.scala 152:32]
          Station6_0_0 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_0_0 <= _GEN_256;
        end
      end else begin
        Station6_0_0 <= _GEN_256;
      end
    end else begin
      Station6_0_0 <= _GEN_256;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2264 & _GEN_2265) begin // @[stationary_dpe.scala 152:32]
          Station6_0_1 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_0_1 <= _GEN_257;
        end
      end else begin
        Station6_0_1 <= _GEN_257;
      end
    end else begin
      Station6_0_1 <= _GEN_257;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2264 & _GEN_2267) begin // @[stationary_dpe.scala 152:32]
          Station6_0_2 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_0_2 <= _GEN_258;
        end
      end else begin
        Station6_0_2 <= _GEN_258;
      end
    end else begin
      Station6_0_2 <= _GEN_258;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2264 & _GEN_2269) begin // @[stationary_dpe.scala 152:32]
          Station6_0_3 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_0_3 <= _GEN_259;
        end
      end else begin
        Station6_0_3 <= _GEN_259;
      end
    end else begin
      Station6_0_3 <= _GEN_259;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2264 & _GEN_2271) begin // @[stationary_dpe.scala 152:32]
          Station6_0_4 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_0_4 <= _GEN_260;
        end
      end else begin
        Station6_0_4 <= _GEN_260;
      end
    end else begin
      Station6_0_4 <= _GEN_260;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2264 & _GEN_2273) begin // @[stationary_dpe.scala 152:32]
          Station6_0_5 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_0_5 <= _GEN_261;
        end
      end else begin
        Station6_0_5 <= _GEN_261;
      end
    end else begin
      Station6_0_5 <= _GEN_261;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2264 & _GEN_2275) begin // @[stationary_dpe.scala 152:32]
          Station6_0_6 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_0_6 <= _GEN_262;
        end
      end else begin
        Station6_0_6 <= _GEN_262;
      end
    end else begin
      Station6_0_6 <= _GEN_262;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2264 & _GEN_2277) begin // @[stationary_dpe.scala 152:32]
          Station6_0_7 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_0_7 <= _GEN_263;
        end
      end else begin
        Station6_0_7 <= _GEN_263;
      end
    end else begin
      Station6_0_7 <= _GEN_263;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2278 & _GEN_2279) begin // @[stationary_dpe.scala 152:32]
          Station6_1_0 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_1_0 <= _GEN_264;
        end
      end else begin
        Station6_1_0 <= _GEN_264;
      end
    end else begin
      Station6_1_0 <= _GEN_264;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2278 & _GEN_2265) begin // @[stationary_dpe.scala 152:32]
          Station6_1_1 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_1_1 <= _GEN_265;
        end
      end else begin
        Station6_1_1 <= _GEN_265;
      end
    end else begin
      Station6_1_1 <= _GEN_265;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2278 & _GEN_2267) begin // @[stationary_dpe.scala 152:32]
          Station6_1_2 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_1_2 <= _GEN_266;
        end
      end else begin
        Station6_1_2 <= _GEN_266;
      end
    end else begin
      Station6_1_2 <= _GEN_266;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2278 & _GEN_2269) begin // @[stationary_dpe.scala 152:32]
          Station6_1_3 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_1_3 <= _GEN_267;
        end
      end else begin
        Station6_1_3 <= _GEN_267;
      end
    end else begin
      Station6_1_3 <= _GEN_267;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2278 & _GEN_2271) begin // @[stationary_dpe.scala 152:32]
          Station6_1_4 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_1_4 <= _GEN_268;
        end
      end else begin
        Station6_1_4 <= _GEN_268;
      end
    end else begin
      Station6_1_4 <= _GEN_268;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2278 & _GEN_2273) begin // @[stationary_dpe.scala 152:32]
          Station6_1_5 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_1_5 <= _GEN_269;
        end
      end else begin
        Station6_1_5 <= _GEN_269;
      end
    end else begin
      Station6_1_5 <= _GEN_269;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2278 & _GEN_2275) begin // @[stationary_dpe.scala 152:32]
          Station6_1_6 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_1_6 <= _GEN_270;
        end
      end else begin
        Station6_1_6 <= _GEN_270;
      end
    end else begin
      Station6_1_6 <= _GEN_270;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2278 & _GEN_2277) begin // @[stationary_dpe.scala 152:32]
          Station6_1_7 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_1_7 <= _GEN_271;
        end
      end else begin
        Station6_1_7 <= _GEN_271;
      end
    end else begin
      Station6_1_7 <= _GEN_271;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2294 & _GEN_2279) begin // @[stationary_dpe.scala 152:32]
          Station6_2_0 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_2_0 <= _GEN_272;
        end
      end else begin
        Station6_2_0 <= _GEN_272;
      end
    end else begin
      Station6_2_0 <= _GEN_272;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2294 & _GEN_2265) begin // @[stationary_dpe.scala 152:32]
          Station6_2_1 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_2_1 <= _GEN_273;
        end
      end else begin
        Station6_2_1 <= _GEN_273;
      end
    end else begin
      Station6_2_1 <= _GEN_273;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2294 & _GEN_2267) begin // @[stationary_dpe.scala 152:32]
          Station6_2_2 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_2_2 <= _GEN_274;
        end
      end else begin
        Station6_2_2 <= _GEN_274;
      end
    end else begin
      Station6_2_2 <= _GEN_274;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2294 & _GEN_2269) begin // @[stationary_dpe.scala 152:32]
          Station6_2_3 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_2_3 <= _GEN_275;
        end
      end else begin
        Station6_2_3 <= _GEN_275;
      end
    end else begin
      Station6_2_3 <= _GEN_275;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2294 & _GEN_2271) begin // @[stationary_dpe.scala 152:32]
          Station6_2_4 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_2_4 <= _GEN_276;
        end
      end else begin
        Station6_2_4 <= _GEN_276;
      end
    end else begin
      Station6_2_4 <= _GEN_276;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2294 & _GEN_2273) begin // @[stationary_dpe.scala 152:32]
          Station6_2_5 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_2_5 <= _GEN_277;
        end
      end else begin
        Station6_2_5 <= _GEN_277;
      end
    end else begin
      Station6_2_5 <= _GEN_277;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2294 & _GEN_2275) begin // @[stationary_dpe.scala 152:32]
          Station6_2_6 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_2_6 <= _GEN_278;
        end
      end else begin
        Station6_2_6 <= _GEN_278;
      end
    end else begin
      Station6_2_6 <= _GEN_278;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2294 & _GEN_2277) begin // @[stationary_dpe.scala 152:32]
          Station6_2_7 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_2_7 <= _GEN_279;
        end
      end else begin
        Station6_2_7 <= _GEN_279;
      end
    end else begin
      Station6_2_7 <= _GEN_279;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2310 & _GEN_2279) begin // @[stationary_dpe.scala 152:32]
          Station6_3_0 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_3_0 <= _GEN_280;
        end
      end else begin
        Station6_3_0 <= _GEN_280;
      end
    end else begin
      Station6_3_0 <= _GEN_280;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2310 & _GEN_2265) begin // @[stationary_dpe.scala 152:32]
          Station6_3_1 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_3_1 <= _GEN_281;
        end
      end else begin
        Station6_3_1 <= _GEN_281;
      end
    end else begin
      Station6_3_1 <= _GEN_281;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2310 & _GEN_2267) begin // @[stationary_dpe.scala 152:32]
          Station6_3_2 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_3_2 <= _GEN_282;
        end
      end else begin
        Station6_3_2 <= _GEN_282;
      end
    end else begin
      Station6_3_2 <= _GEN_282;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2310 & _GEN_2269) begin // @[stationary_dpe.scala 152:32]
          Station6_3_3 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_3_3 <= _GEN_283;
        end
      end else begin
        Station6_3_3 <= _GEN_283;
      end
    end else begin
      Station6_3_3 <= _GEN_283;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2310 & _GEN_2271) begin // @[stationary_dpe.scala 152:32]
          Station6_3_4 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_3_4 <= _GEN_284;
        end
      end else begin
        Station6_3_4 <= _GEN_284;
      end
    end else begin
      Station6_3_4 <= _GEN_284;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2310 & _GEN_2273) begin // @[stationary_dpe.scala 152:32]
          Station6_3_5 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_3_5 <= _GEN_285;
        end
      end else begin
        Station6_3_5 <= _GEN_285;
      end
    end else begin
      Station6_3_5 <= _GEN_285;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2310 & _GEN_2275) begin // @[stationary_dpe.scala 152:32]
          Station6_3_6 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_3_6 <= _GEN_286;
        end
      end else begin
        Station6_3_6 <= _GEN_286;
      end
    end else begin
      Station6_3_6 <= _GEN_286;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2310 & _GEN_2277) begin // @[stationary_dpe.scala 152:32]
          Station6_3_7 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_3_7 <= _GEN_287;
        end
      end else begin
        Station6_3_7 <= _GEN_287;
      end
    end else begin
      Station6_3_7 <= _GEN_287;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2326 & _GEN_2279) begin // @[stationary_dpe.scala 152:32]
          Station6_4_0 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_4_0 <= _GEN_288;
        end
      end else begin
        Station6_4_0 <= _GEN_288;
      end
    end else begin
      Station6_4_0 <= _GEN_288;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2326 & _GEN_2265) begin // @[stationary_dpe.scala 152:32]
          Station6_4_1 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_4_1 <= _GEN_289;
        end
      end else begin
        Station6_4_1 <= _GEN_289;
      end
    end else begin
      Station6_4_1 <= _GEN_289;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2326 & _GEN_2267) begin // @[stationary_dpe.scala 152:32]
          Station6_4_2 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_4_2 <= _GEN_290;
        end
      end else begin
        Station6_4_2 <= _GEN_290;
      end
    end else begin
      Station6_4_2 <= _GEN_290;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2326 & _GEN_2269) begin // @[stationary_dpe.scala 152:32]
          Station6_4_3 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_4_3 <= _GEN_291;
        end
      end else begin
        Station6_4_3 <= _GEN_291;
      end
    end else begin
      Station6_4_3 <= _GEN_291;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2326 & _GEN_2271) begin // @[stationary_dpe.scala 152:32]
          Station6_4_4 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_4_4 <= _GEN_292;
        end
      end else begin
        Station6_4_4 <= _GEN_292;
      end
    end else begin
      Station6_4_4 <= _GEN_292;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2326 & _GEN_2273) begin // @[stationary_dpe.scala 152:32]
          Station6_4_5 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_4_5 <= _GEN_293;
        end
      end else begin
        Station6_4_5 <= _GEN_293;
      end
    end else begin
      Station6_4_5 <= _GEN_293;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2326 & _GEN_2275) begin // @[stationary_dpe.scala 152:32]
          Station6_4_6 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_4_6 <= _GEN_294;
        end
      end else begin
        Station6_4_6 <= _GEN_294;
      end
    end else begin
      Station6_4_6 <= _GEN_294;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2326 & _GEN_2277) begin // @[stationary_dpe.scala 152:32]
          Station6_4_7 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_4_7 <= _GEN_295;
        end
      end else begin
        Station6_4_7 <= _GEN_295;
      end
    end else begin
      Station6_4_7 <= _GEN_295;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2342 & _GEN_2279) begin // @[stationary_dpe.scala 152:32]
          Station6_5_0 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_5_0 <= _GEN_296;
        end
      end else begin
        Station6_5_0 <= _GEN_296;
      end
    end else begin
      Station6_5_0 <= _GEN_296;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2342 & _GEN_2265) begin // @[stationary_dpe.scala 152:32]
          Station6_5_1 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_5_1 <= _GEN_297;
        end
      end else begin
        Station6_5_1 <= _GEN_297;
      end
    end else begin
      Station6_5_1 <= _GEN_297;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2342 & _GEN_2267) begin // @[stationary_dpe.scala 152:32]
          Station6_5_2 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_5_2 <= _GEN_298;
        end
      end else begin
        Station6_5_2 <= _GEN_298;
      end
    end else begin
      Station6_5_2 <= _GEN_298;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2342 & _GEN_2269) begin // @[stationary_dpe.scala 152:32]
          Station6_5_3 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_5_3 <= _GEN_299;
        end
      end else begin
        Station6_5_3 <= _GEN_299;
      end
    end else begin
      Station6_5_3 <= _GEN_299;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2342 & _GEN_2271) begin // @[stationary_dpe.scala 152:32]
          Station6_5_4 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_5_4 <= _GEN_300;
        end
      end else begin
        Station6_5_4 <= _GEN_300;
      end
    end else begin
      Station6_5_4 <= _GEN_300;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2342 & _GEN_2273) begin // @[stationary_dpe.scala 152:32]
          Station6_5_5 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_5_5 <= _GEN_301;
        end
      end else begin
        Station6_5_5 <= _GEN_301;
      end
    end else begin
      Station6_5_5 <= _GEN_301;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2342 & _GEN_2275) begin // @[stationary_dpe.scala 152:32]
          Station6_5_6 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_5_6 <= _GEN_302;
        end
      end else begin
        Station6_5_6 <= _GEN_302;
      end
    end else begin
      Station6_5_6 <= _GEN_302;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2342 & _GEN_2277) begin // @[stationary_dpe.scala 152:32]
          Station6_5_7 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_5_7 <= _GEN_303;
        end
      end else begin
        Station6_5_7 <= _GEN_303;
      end
    end else begin
      Station6_5_7 <= _GEN_303;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2358 & _GEN_2279) begin // @[stationary_dpe.scala 152:32]
          Station6_6_0 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_6_0 <= _GEN_304;
        end
      end else begin
        Station6_6_0 <= _GEN_304;
      end
    end else begin
      Station6_6_0 <= _GEN_304;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2358 & _GEN_2265) begin // @[stationary_dpe.scala 152:32]
          Station6_6_1 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_6_1 <= _GEN_305;
        end
      end else begin
        Station6_6_1 <= _GEN_305;
      end
    end else begin
      Station6_6_1 <= _GEN_305;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2358 & _GEN_2267) begin // @[stationary_dpe.scala 152:32]
          Station6_6_2 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_6_2 <= _GEN_306;
        end
      end else begin
        Station6_6_2 <= _GEN_306;
      end
    end else begin
      Station6_6_2 <= _GEN_306;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2358 & _GEN_2269) begin // @[stationary_dpe.scala 152:32]
          Station6_6_3 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_6_3 <= _GEN_307;
        end
      end else begin
        Station6_6_3 <= _GEN_307;
      end
    end else begin
      Station6_6_3 <= _GEN_307;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2358 & _GEN_2271) begin // @[stationary_dpe.scala 152:32]
          Station6_6_4 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_6_4 <= _GEN_308;
        end
      end else begin
        Station6_6_4 <= _GEN_308;
      end
    end else begin
      Station6_6_4 <= _GEN_308;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2358 & _GEN_2273) begin // @[stationary_dpe.scala 152:32]
          Station6_6_5 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_6_5 <= _GEN_309;
        end
      end else begin
        Station6_6_5 <= _GEN_309;
      end
    end else begin
      Station6_6_5 <= _GEN_309;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2358 & _GEN_2275) begin // @[stationary_dpe.scala 152:32]
          Station6_6_6 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_6_6 <= _GEN_310;
        end
      end else begin
        Station6_6_6 <= _GEN_310;
      end
    end else begin
      Station6_6_6 <= _GEN_310;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2358 & _GEN_2277) begin // @[stationary_dpe.scala 152:32]
          Station6_6_7 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_6_7 <= _GEN_311;
        end
      end else begin
        Station6_6_7 <= _GEN_311;
      end
    end else begin
      Station6_6_7 <= _GEN_311;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2374 & _GEN_2279) begin // @[stationary_dpe.scala 152:32]
          Station6_7_0 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_7_0 <= _GEN_312;
        end
      end else begin
        Station6_7_0 <= _GEN_312;
      end
    end else begin
      Station6_7_0 <= _GEN_312;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2374 & _GEN_2265) begin // @[stationary_dpe.scala 152:32]
          Station6_7_1 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_7_1 <= _GEN_313;
        end
      end else begin
        Station6_7_1 <= _GEN_313;
      end
    end else begin
      Station6_7_1 <= _GEN_313;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2374 & _GEN_2267) begin // @[stationary_dpe.scala 152:32]
          Station6_7_2 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_7_2 <= _GEN_314;
        end
      end else begin
        Station6_7_2 <= _GEN_314;
      end
    end else begin
      Station6_7_2 <= _GEN_314;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2374 & _GEN_2269) begin // @[stationary_dpe.scala 152:32]
          Station6_7_3 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_7_3 <= _GEN_315;
        end
      end else begin
        Station6_7_3 <= _GEN_315;
      end
    end else begin
      Station6_7_3 <= _GEN_315;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2374 & _GEN_2271) begin // @[stationary_dpe.scala 152:32]
          Station6_7_4 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_7_4 <= _GEN_316;
        end
      end else begin
        Station6_7_4 <= _GEN_316;
      end
    end else begin
      Station6_7_4 <= _GEN_316;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2374 & _GEN_2273) begin // @[stationary_dpe.scala 152:32]
          Station6_7_5 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_7_5 <= _GEN_317;
        end
      end else begin
        Station6_7_5 <= _GEN_317;
      end
    end else begin
      Station6_7_5 <= _GEN_317;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2374 & _GEN_2275) begin // @[stationary_dpe.scala 152:32]
          Station6_7_6 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_7_6 <= _GEN_318;
        end
      end else begin
        Station6_7_6 <= _GEN_318;
      end
    end else begin
      Station6_7_6 <= _GEN_318;
    end
    if (~valid4) begin // @[stationary_dpe.scala 150:28]
      if (_GEN_1543 != 16'h0) begin // @[stationary_dpe.scala 151:39]
        if (_GEN_2374 & _GEN_2277) begin // @[stationary_dpe.scala 152:32]
          Station6_7_7 <= 16'h0; // @[stationary_dpe.scala 152:32]
        end else begin
          Station6_7_7 <= _GEN_319;
        end
      end else begin
        Station6_7_7 <= _GEN_319;
      end
    end else begin
      Station6_7_7 <= _GEN_319;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2264 & _GEN_2279) begin // @[stationary_dpe.scala 164:32]
          Station7_0_0 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_0_0 <= _GEN_320;
        end
      end else begin
        Station7_0_0 <= _GEN_320;
      end
    end else begin
      Station7_0_0 <= _GEN_320;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2264 & _GEN_2265) begin // @[stationary_dpe.scala 164:32]
          Station7_0_1 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_0_1 <= _GEN_321;
        end
      end else begin
        Station7_0_1 <= _GEN_321;
      end
    end else begin
      Station7_0_1 <= _GEN_321;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2264 & _GEN_2267) begin // @[stationary_dpe.scala 164:32]
          Station7_0_2 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_0_2 <= _GEN_322;
        end
      end else begin
        Station7_0_2 <= _GEN_322;
      end
    end else begin
      Station7_0_2 <= _GEN_322;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2264 & _GEN_2269) begin // @[stationary_dpe.scala 164:32]
          Station7_0_3 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_0_3 <= _GEN_323;
        end
      end else begin
        Station7_0_3 <= _GEN_323;
      end
    end else begin
      Station7_0_3 <= _GEN_323;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2264 & _GEN_2271) begin // @[stationary_dpe.scala 164:32]
          Station7_0_4 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_0_4 <= _GEN_324;
        end
      end else begin
        Station7_0_4 <= _GEN_324;
      end
    end else begin
      Station7_0_4 <= _GEN_324;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2264 & _GEN_2273) begin // @[stationary_dpe.scala 164:32]
          Station7_0_5 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_0_5 <= _GEN_325;
        end
      end else begin
        Station7_0_5 <= _GEN_325;
      end
    end else begin
      Station7_0_5 <= _GEN_325;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2264 & _GEN_2275) begin // @[stationary_dpe.scala 164:32]
          Station7_0_6 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_0_6 <= _GEN_326;
        end
      end else begin
        Station7_0_6 <= _GEN_326;
      end
    end else begin
      Station7_0_6 <= _GEN_326;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2264 & _GEN_2277) begin // @[stationary_dpe.scala 164:32]
          Station7_0_7 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_0_7 <= _GEN_327;
        end
      end else begin
        Station7_0_7 <= _GEN_327;
      end
    end else begin
      Station7_0_7 <= _GEN_327;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2278 & _GEN_2279) begin // @[stationary_dpe.scala 164:32]
          Station7_1_0 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_1_0 <= _GEN_328;
        end
      end else begin
        Station7_1_0 <= _GEN_328;
      end
    end else begin
      Station7_1_0 <= _GEN_328;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2278 & _GEN_2265) begin // @[stationary_dpe.scala 164:32]
          Station7_1_1 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_1_1 <= _GEN_329;
        end
      end else begin
        Station7_1_1 <= _GEN_329;
      end
    end else begin
      Station7_1_1 <= _GEN_329;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2278 & _GEN_2267) begin // @[stationary_dpe.scala 164:32]
          Station7_1_2 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_1_2 <= _GEN_330;
        end
      end else begin
        Station7_1_2 <= _GEN_330;
      end
    end else begin
      Station7_1_2 <= _GEN_330;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2278 & _GEN_2269) begin // @[stationary_dpe.scala 164:32]
          Station7_1_3 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_1_3 <= _GEN_331;
        end
      end else begin
        Station7_1_3 <= _GEN_331;
      end
    end else begin
      Station7_1_3 <= _GEN_331;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2278 & _GEN_2271) begin // @[stationary_dpe.scala 164:32]
          Station7_1_4 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_1_4 <= _GEN_332;
        end
      end else begin
        Station7_1_4 <= _GEN_332;
      end
    end else begin
      Station7_1_4 <= _GEN_332;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2278 & _GEN_2273) begin // @[stationary_dpe.scala 164:32]
          Station7_1_5 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_1_5 <= _GEN_333;
        end
      end else begin
        Station7_1_5 <= _GEN_333;
      end
    end else begin
      Station7_1_5 <= _GEN_333;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2278 & _GEN_2275) begin // @[stationary_dpe.scala 164:32]
          Station7_1_6 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_1_6 <= _GEN_334;
        end
      end else begin
        Station7_1_6 <= _GEN_334;
      end
    end else begin
      Station7_1_6 <= _GEN_334;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2278 & _GEN_2277) begin // @[stationary_dpe.scala 164:32]
          Station7_1_7 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_1_7 <= _GEN_335;
        end
      end else begin
        Station7_1_7 <= _GEN_335;
      end
    end else begin
      Station7_1_7 <= _GEN_335;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2294 & _GEN_2279) begin // @[stationary_dpe.scala 164:32]
          Station7_2_0 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_2_0 <= _GEN_336;
        end
      end else begin
        Station7_2_0 <= _GEN_336;
      end
    end else begin
      Station7_2_0 <= _GEN_336;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2294 & _GEN_2265) begin // @[stationary_dpe.scala 164:32]
          Station7_2_1 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_2_1 <= _GEN_337;
        end
      end else begin
        Station7_2_1 <= _GEN_337;
      end
    end else begin
      Station7_2_1 <= _GEN_337;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2294 & _GEN_2267) begin // @[stationary_dpe.scala 164:32]
          Station7_2_2 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_2_2 <= _GEN_338;
        end
      end else begin
        Station7_2_2 <= _GEN_338;
      end
    end else begin
      Station7_2_2 <= _GEN_338;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2294 & _GEN_2269) begin // @[stationary_dpe.scala 164:32]
          Station7_2_3 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_2_3 <= _GEN_339;
        end
      end else begin
        Station7_2_3 <= _GEN_339;
      end
    end else begin
      Station7_2_3 <= _GEN_339;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2294 & _GEN_2271) begin // @[stationary_dpe.scala 164:32]
          Station7_2_4 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_2_4 <= _GEN_340;
        end
      end else begin
        Station7_2_4 <= _GEN_340;
      end
    end else begin
      Station7_2_4 <= _GEN_340;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2294 & _GEN_2273) begin // @[stationary_dpe.scala 164:32]
          Station7_2_5 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_2_5 <= _GEN_341;
        end
      end else begin
        Station7_2_5 <= _GEN_341;
      end
    end else begin
      Station7_2_5 <= _GEN_341;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2294 & _GEN_2275) begin // @[stationary_dpe.scala 164:32]
          Station7_2_6 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_2_6 <= _GEN_342;
        end
      end else begin
        Station7_2_6 <= _GEN_342;
      end
    end else begin
      Station7_2_6 <= _GEN_342;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2294 & _GEN_2277) begin // @[stationary_dpe.scala 164:32]
          Station7_2_7 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_2_7 <= _GEN_343;
        end
      end else begin
        Station7_2_7 <= _GEN_343;
      end
    end else begin
      Station7_2_7 <= _GEN_343;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2310 & _GEN_2279) begin // @[stationary_dpe.scala 164:32]
          Station7_3_0 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_3_0 <= _GEN_344;
        end
      end else begin
        Station7_3_0 <= _GEN_344;
      end
    end else begin
      Station7_3_0 <= _GEN_344;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2310 & _GEN_2265) begin // @[stationary_dpe.scala 164:32]
          Station7_3_1 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_3_1 <= _GEN_345;
        end
      end else begin
        Station7_3_1 <= _GEN_345;
      end
    end else begin
      Station7_3_1 <= _GEN_345;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2310 & _GEN_2267) begin // @[stationary_dpe.scala 164:32]
          Station7_3_2 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_3_2 <= _GEN_346;
        end
      end else begin
        Station7_3_2 <= _GEN_346;
      end
    end else begin
      Station7_3_2 <= _GEN_346;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2310 & _GEN_2269) begin // @[stationary_dpe.scala 164:32]
          Station7_3_3 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_3_3 <= _GEN_347;
        end
      end else begin
        Station7_3_3 <= _GEN_347;
      end
    end else begin
      Station7_3_3 <= _GEN_347;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2310 & _GEN_2271) begin // @[stationary_dpe.scala 164:32]
          Station7_3_4 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_3_4 <= _GEN_348;
        end
      end else begin
        Station7_3_4 <= _GEN_348;
      end
    end else begin
      Station7_3_4 <= _GEN_348;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2310 & _GEN_2273) begin // @[stationary_dpe.scala 164:32]
          Station7_3_5 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_3_5 <= _GEN_349;
        end
      end else begin
        Station7_3_5 <= _GEN_349;
      end
    end else begin
      Station7_3_5 <= _GEN_349;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2310 & _GEN_2275) begin // @[stationary_dpe.scala 164:32]
          Station7_3_6 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_3_6 <= _GEN_350;
        end
      end else begin
        Station7_3_6 <= _GEN_350;
      end
    end else begin
      Station7_3_6 <= _GEN_350;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2310 & _GEN_2277) begin // @[stationary_dpe.scala 164:32]
          Station7_3_7 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_3_7 <= _GEN_351;
        end
      end else begin
        Station7_3_7 <= _GEN_351;
      end
    end else begin
      Station7_3_7 <= _GEN_351;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2326 & _GEN_2279) begin // @[stationary_dpe.scala 164:32]
          Station7_4_0 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_4_0 <= _GEN_352;
        end
      end else begin
        Station7_4_0 <= _GEN_352;
      end
    end else begin
      Station7_4_0 <= _GEN_352;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2326 & _GEN_2265) begin // @[stationary_dpe.scala 164:32]
          Station7_4_1 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_4_1 <= _GEN_353;
        end
      end else begin
        Station7_4_1 <= _GEN_353;
      end
    end else begin
      Station7_4_1 <= _GEN_353;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2326 & _GEN_2267) begin // @[stationary_dpe.scala 164:32]
          Station7_4_2 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_4_2 <= _GEN_354;
        end
      end else begin
        Station7_4_2 <= _GEN_354;
      end
    end else begin
      Station7_4_2 <= _GEN_354;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2326 & _GEN_2269) begin // @[stationary_dpe.scala 164:32]
          Station7_4_3 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_4_3 <= _GEN_355;
        end
      end else begin
        Station7_4_3 <= _GEN_355;
      end
    end else begin
      Station7_4_3 <= _GEN_355;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2326 & _GEN_2271) begin // @[stationary_dpe.scala 164:32]
          Station7_4_4 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_4_4 <= _GEN_356;
        end
      end else begin
        Station7_4_4 <= _GEN_356;
      end
    end else begin
      Station7_4_4 <= _GEN_356;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2326 & _GEN_2273) begin // @[stationary_dpe.scala 164:32]
          Station7_4_5 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_4_5 <= _GEN_357;
        end
      end else begin
        Station7_4_5 <= _GEN_357;
      end
    end else begin
      Station7_4_5 <= _GEN_357;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2326 & _GEN_2275) begin // @[stationary_dpe.scala 164:32]
          Station7_4_6 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_4_6 <= _GEN_358;
        end
      end else begin
        Station7_4_6 <= _GEN_358;
      end
    end else begin
      Station7_4_6 <= _GEN_358;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2326 & _GEN_2277) begin // @[stationary_dpe.scala 164:32]
          Station7_4_7 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_4_7 <= _GEN_359;
        end
      end else begin
        Station7_4_7 <= _GEN_359;
      end
    end else begin
      Station7_4_7 <= _GEN_359;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2342 & _GEN_2279) begin // @[stationary_dpe.scala 164:32]
          Station7_5_0 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_5_0 <= _GEN_360;
        end
      end else begin
        Station7_5_0 <= _GEN_360;
      end
    end else begin
      Station7_5_0 <= _GEN_360;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2342 & _GEN_2265) begin // @[stationary_dpe.scala 164:32]
          Station7_5_1 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_5_1 <= _GEN_361;
        end
      end else begin
        Station7_5_1 <= _GEN_361;
      end
    end else begin
      Station7_5_1 <= _GEN_361;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2342 & _GEN_2267) begin // @[stationary_dpe.scala 164:32]
          Station7_5_2 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_5_2 <= _GEN_362;
        end
      end else begin
        Station7_5_2 <= _GEN_362;
      end
    end else begin
      Station7_5_2 <= _GEN_362;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2342 & _GEN_2269) begin // @[stationary_dpe.scala 164:32]
          Station7_5_3 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_5_3 <= _GEN_363;
        end
      end else begin
        Station7_5_3 <= _GEN_363;
      end
    end else begin
      Station7_5_3 <= _GEN_363;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2342 & _GEN_2271) begin // @[stationary_dpe.scala 164:32]
          Station7_5_4 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_5_4 <= _GEN_364;
        end
      end else begin
        Station7_5_4 <= _GEN_364;
      end
    end else begin
      Station7_5_4 <= _GEN_364;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2342 & _GEN_2273) begin // @[stationary_dpe.scala 164:32]
          Station7_5_5 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_5_5 <= _GEN_365;
        end
      end else begin
        Station7_5_5 <= _GEN_365;
      end
    end else begin
      Station7_5_5 <= _GEN_365;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2342 & _GEN_2275) begin // @[stationary_dpe.scala 164:32]
          Station7_5_6 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_5_6 <= _GEN_366;
        end
      end else begin
        Station7_5_6 <= _GEN_366;
      end
    end else begin
      Station7_5_6 <= _GEN_366;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2342 & _GEN_2277) begin // @[stationary_dpe.scala 164:32]
          Station7_5_7 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_5_7 <= _GEN_367;
        end
      end else begin
        Station7_5_7 <= _GEN_367;
      end
    end else begin
      Station7_5_7 <= _GEN_367;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2358 & _GEN_2279) begin // @[stationary_dpe.scala 164:32]
          Station7_6_0 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_6_0 <= _GEN_368;
        end
      end else begin
        Station7_6_0 <= _GEN_368;
      end
    end else begin
      Station7_6_0 <= _GEN_368;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2358 & _GEN_2265) begin // @[stationary_dpe.scala 164:32]
          Station7_6_1 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_6_1 <= _GEN_369;
        end
      end else begin
        Station7_6_1 <= _GEN_369;
      end
    end else begin
      Station7_6_1 <= _GEN_369;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2358 & _GEN_2267) begin // @[stationary_dpe.scala 164:32]
          Station7_6_2 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_6_2 <= _GEN_370;
        end
      end else begin
        Station7_6_2 <= _GEN_370;
      end
    end else begin
      Station7_6_2 <= _GEN_370;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2358 & _GEN_2269) begin // @[stationary_dpe.scala 164:32]
          Station7_6_3 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_6_3 <= _GEN_371;
        end
      end else begin
        Station7_6_3 <= _GEN_371;
      end
    end else begin
      Station7_6_3 <= _GEN_371;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2358 & _GEN_2271) begin // @[stationary_dpe.scala 164:32]
          Station7_6_4 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_6_4 <= _GEN_372;
        end
      end else begin
        Station7_6_4 <= _GEN_372;
      end
    end else begin
      Station7_6_4 <= _GEN_372;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2358 & _GEN_2273) begin // @[stationary_dpe.scala 164:32]
          Station7_6_5 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_6_5 <= _GEN_373;
        end
      end else begin
        Station7_6_5 <= _GEN_373;
      end
    end else begin
      Station7_6_5 <= _GEN_373;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2358 & _GEN_2275) begin // @[stationary_dpe.scala 164:32]
          Station7_6_6 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_6_6 <= _GEN_374;
        end
      end else begin
        Station7_6_6 <= _GEN_374;
      end
    end else begin
      Station7_6_6 <= _GEN_374;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2358 & _GEN_2277) begin // @[stationary_dpe.scala 164:32]
          Station7_6_7 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_6_7 <= _GEN_375;
        end
      end else begin
        Station7_6_7 <= _GEN_375;
      end
    end else begin
      Station7_6_7 <= _GEN_375;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2374 & _GEN_2279) begin // @[stationary_dpe.scala 164:32]
          Station7_7_0 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_7_0 <= _GEN_376;
        end
      end else begin
        Station7_7_0 <= _GEN_376;
      end
    end else begin
      Station7_7_0 <= _GEN_376;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2374 & _GEN_2265) begin // @[stationary_dpe.scala 164:32]
          Station7_7_1 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_7_1 <= _GEN_377;
        end
      end else begin
        Station7_7_1 <= _GEN_377;
      end
    end else begin
      Station7_7_1 <= _GEN_377;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2374 & _GEN_2267) begin // @[stationary_dpe.scala 164:32]
          Station7_7_2 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_7_2 <= _GEN_378;
        end
      end else begin
        Station7_7_2 <= _GEN_378;
      end
    end else begin
      Station7_7_2 <= _GEN_378;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2374 & _GEN_2269) begin // @[stationary_dpe.scala 164:32]
          Station7_7_3 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_7_3 <= _GEN_379;
        end
      end else begin
        Station7_7_3 <= _GEN_379;
      end
    end else begin
      Station7_7_3 <= _GEN_379;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2374 & _GEN_2271) begin // @[stationary_dpe.scala 164:32]
          Station7_7_4 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_7_4 <= _GEN_380;
        end
      end else begin
        Station7_7_4 <= _GEN_380;
      end
    end else begin
      Station7_7_4 <= _GEN_380;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2374 & _GEN_2273) begin // @[stationary_dpe.scala 164:32]
          Station7_7_5 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_7_5 <= _GEN_381;
        end
      end else begin
        Station7_7_5 <= _GEN_381;
      end
    end else begin
      Station7_7_5 <= _GEN_381;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2374 & _GEN_2275) begin // @[stationary_dpe.scala 164:32]
          Station7_7_6 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_7_6 <= _GEN_382;
        end
      end else begin
        Station7_7_6 <= _GEN_382;
      end
    end else begin
      Station7_7_6 <= _GEN_382;
    end
    if (~valid5) begin // @[stationary_dpe.scala 162:28]
      if (_GEN_1801 != 16'h0) begin // @[stationary_dpe.scala 163:39]
        if (_GEN_2374 & _GEN_2277) begin // @[stationary_dpe.scala 164:32]
          Station7_7_7 <= 16'h0; // @[stationary_dpe.scala 164:32]
        end else begin
          Station7_7_7 <= _GEN_383;
        end
      end else begin
        Station7_7_7 <= _GEN_383;
      end
    end else begin
      Station7_7_7 <= _GEN_383;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2264 & _GEN_2279) begin // @[stationary_dpe.scala 176:32]
          Station8_0_0 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_0_0 <= _GEN_384;
        end
      end else begin
        Station8_0_0 <= _GEN_384;
      end
    end else begin
      Station8_0_0 <= _GEN_384;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2264 & _GEN_2265) begin // @[stationary_dpe.scala 176:32]
          Station8_0_1 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_0_1 <= _GEN_385;
        end
      end else begin
        Station8_0_1 <= _GEN_385;
      end
    end else begin
      Station8_0_1 <= _GEN_385;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2264 & _GEN_2267) begin // @[stationary_dpe.scala 176:32]
          Station8_0_2 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_0_2 <= _GEN_386;
        end
      end else begin
        Station8_0_2 <= _GEN_386;
      end
    end else begin
      Station8_0_2 <= _GEN_386;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2264 & _GEN_2269) begin // @[stationary_dpe.scala 176:32]
          Station8_0_3 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_0_3 <= _GEN_387;
        end
      end else begin
        Station8_0_3 <= _GEN_387;
      end
    end else begin
      Station8_0_3 <= _GEN_387;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2264 & _GEN_2271) begin // @[stationary_dpe.scala 176:32]
          Station8_0_4 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_0_4 <= _GEN_388;
        end
      end else begin
        Station8_0_4 <= _GEN_388;
      end
    end else begin
      Station8_0_4 <= _GEN_388;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2264 & _GEN_2273) begin // @[stationary_dpe.scala 176:32]
          Station8_0_5 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_0_5 <= _GEN_389;
        end
      end else begin
        Station8_0_5 <= _GEN_389;
      end
    end else begin
      Station8_0_5 <= _GEN_389;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2264 & _GEN_2275) begin // @[stationary_dpe.scala 176:32]
          Station8_0_6 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_0_6 <= _GEN_390;
        end
      end else begin
        Station8_0_6 <= _GEN_390;
      end
    end else begin
      Station8_0_6 <= _GEN_390;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2264 & _GEN_2277) begin // @[stationary_dpe.scala 176:32]
          Station8_0_7 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_0_7 <= _GEN_391;
        end
      end else begin
        Station8_0_7 <= _GEN_391;
      end
    end else begin
      Station8_0_7 <= _GEN_391;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2278 & _GEN_2279) begin // @[stationary_dpe.scala 176:32]
          Station8_1_0 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_1_0 <= _GEN_392;
        end
      end else begin
        Station8_1_0 <= _GEN_392;
      end
    end else begin
      Station8_1_0 <= _GEN_392;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2278 & _GEN_2265) begin // @[stationary_dpe.scala 176:32]
          Station8_1_1 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_1_1 <= _GEN_393;
        end
      end else begin
        Station8_1_1 <= _GEN_393;
      end
    end else begin
      Station8_1_1 <= _GEN_393;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2278 & _GEN_2267) begin // @[stationary_dpe.scala 176:32]
          Station8_1_2 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_1_2 <= _GEN_394;
        end
      end else begin
        Station8_1_2 <= _GEN_394;
      end
    end else begin
      Station8_1_2 <= _GEN_394;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2278 & _GEN_2269) begin // @[stationary_dpe.scala 176:32]
          Station8_1_3 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_1_3 <= _GEN_395;
        end
      end else begin
        Station8_1_3 <= _GEN_395;
      end
    end else begin
      Station8_1_3 <= _GEN_395;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2278 & _GEN_2271) begin // @[stationary_dpe.scala 176:32]
          Station8_1_4 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_1_4 <= _GEN_396;
        end
      end else begin
        Station8_1_4 <= _GEN_396;
      end
    end else begin
      Station8_1_4 <= _GEN_396;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2278 & _GEN_2273) begin // @[stationary_dpe.scala 176:32]
          Station8_1_5 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_1_5 <= _GEN_397;
        end
      end else begin
        Station8_1_5 <= _GEN_397;
      end
    end else begin
      Station8_1_5 <= _GEN_397;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2278 & _GEN_2275) begin // @[stationary_dpe.scala 176:32]
          Station8_1_6 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_1_6 <= _GEN_398;
        end
      end else begin
        Station8_1_6 <= _GEN_398;
      end
    end else begin
      Station8_1_6 <= _GEN_398;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2278 & _GEN_2277) begin // @[stationary_dpe.scala 176:32]
          Station8_1_7 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_1_7 <= _GEN_399;
        end
      end else begin
        Station8_1_7 <= _GEN_399;
      end
    end else begin
      Station8_1_7 <= _GEN_399;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2294 & _GEN_2279) begin // @[stationary_dpe.scala 176:32]
          Station8_2_0 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_2_0 <= _GEN_400;
        end
      end else begin
        Station8_2_0 <= _GEN_400;
      end
    end else begin
      Station8_2_0 <= _GEN_400;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2294 & _GEN_2265) begin // @[stationary_dpe.scala 176:32]
          Station8_2_1 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_2_1 <= _GEN_401;
        end
      end else begin
        Station8_2_1 <= _GEN_401;
      end
    end else begin
      Station8_2_1 <= _GEN_401;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2294 & _GEN_2267) begin // @[stationary_dpe.scala 176:32]
          Station8_2_2 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_2_2 <= _GEN_402;
        end
      end else begin
        Station8_2_2 <= _GEN_402;
      end
    end else begin
      Station8_2_2 <= _GEN_402;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2294 & _GEN_2269) begin // @[stationary_dpe.scala 176:32]
          Station8_2_3 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_2_3 <= _GEN_403;
        end
      end else begin
        Station8_2_3 <= _GEN_403;
      end
    end else begin
      Station8_2_3 <= _GEN_403;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2294 & _GEN_2271) begin // @[stationary_dpe.scala 176:32]
          Station8_2_4 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_2_4 <= _GEN_404;
        end
      end else begin
        Station8_2_4 <= _GEN_404;
      end
    end else begin
      Station8_2_4 <= _GEN_404;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2294 & _GEN_2273) begin // @[stationary_dpe.scala 176:32]
          Station8_2_5 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_2_5 <= _GEN_405;
        end
      end else begin
        Station8_2_5 <= _GEN_405;
      end
    end else begin
      Station8_2_5 <= _GEN_405;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2294 & _GEN_2275) begin // @[stationary_dpe.scala 176:32]
          Station8_2_6 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_2_6 <= _GEN_406;
        end
      end else begin
        Station8_2_6 <= _GEN_406;
      end
    end else begin
      Station8_2_6 <= _GEN_406;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2294 & _GEN_2277) begin // @[stationary_dpe.scala 176:32]
          Station8_2_7 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_2_7 <= _GEN_407;
        end
      end else begin
        Station8_2_7 <= _GEN_407;
      end
    end else begin
      Station8_2_7 <= _GEN_407;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2310 & _GEN_2279) begin // @[stationary_dpe.scala 176:32]
          Station8_3_0 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_3_0 <= _GEN_408;
        end
      end else begin
        Station8_3_0 <= _GEN_408;
      end
    end else begin
      Station8_3_0 <= _GEN_408;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2310 & _GEN_2265) begin // @[stationary_dpe.scala 176:32]
          Station8_3_1 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_3_1 <= _GEN_409;
        end
      end else begin
        Station8_3_1 <= _GEN_409;
      end
    end else begin
      Station8_3_1 <= _GEN_409;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2310 & _GEN_2267) begin // @[stationary_dpe.scala 176:32]
          Station8_3_2 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_3_2 <= _GEN_410;
        end
      end else begin
        Station8_3_2 <= _GEN_410;
      end
    end else begin
      Station8_3_2 <= _GEN_410;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2310 & _GEN_2269) begin // @[stationary_dpe.scala 176:32]
          Station8_3_3 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_3_3 <= _GEN_411;
        end
      end else begin
        Station8_3_3 <= _GEN_411;
      end
    end else begin
      Station8_3_3 <= _GEN_411;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2310 & _GEN_2271) begin // @[stationary_dpe.scala 176:32]
          Station8_3_4 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_3_4 <= _GEN_412;
        end
      end else begin
        Station8_3_4 <= _GEN_412;
      end
    end else begin
      Station8_3_4 <= _GEN_412;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2310 & _GEN_2273) begin // @[stationary_dpe.scala 176:32]
          Station8_3_5 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_3_5 <= _GEN_413;
        end
      end else begin
        Station8_3_5 <= _GEN_413;
      end
    end else begin
      Station8_3_5 <= _GEN_413;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2310 & _GEN_2275) begin // @[stationary_dpe.scala 176:32]
          Station8_3_6 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_3_6 <= _GEN_414;
        end
      end else begin
        Station8_3_6 <= _GEN_414;
      end
    end else begin
      Station8_3_6 <= _GEN_414;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2310 & _GEN_2277) begin // @[stationary_dpe.scala 176:32]
          Station8_3_7 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_3_7 <= _GEN_415;
        end
      end else begin
        Station8_3_7 <= _GEN_415;
      end
    end else begin
      Station8_3_7 <= _GEN_415;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2326 & _GEN_2279) begin // @[stationary_dpe.scala 176:32]
          Station8_4_0 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_4_0 <= _GEN_416;
        end
      end else begin
        Station8_4_0 <= _GEN_416;
      end
    end else begin
      Station8_4_0 <= _GEN_416;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2326 & _GEN_2265) begin // @[stationary_dpe.scala 176:32]
          Station8_4_1 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_4_1 <= _GEN_417;
        end
      end else begin
        Station8_4_1 <= _GEN_417;
      end
    end else begin
      Station8_4_1 <= _GEN_417;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2326 & _GEN_2267) begin // @[stationary_dpe.scala 176:32]
          Station8_4_2 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_4_2 <= _GEN_418;
        end
      end else begin
        Station8_4_2 <= _GEN_418;
      end
    end else begin
      Station8_4_2 <= _GEN_418;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2326 & _GEN_2269) begin // @[stationary_dpe.scala 176:32]
          Station8_4_3 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_4_3 <= _GEN_419;
        end
      end else begin
        Station8_4_3 <= _GEN_419;
      end
    end else begin
      Station8_4_3 <= _GEN_419;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2326 & _GEN_2271) begin // @[stationary_dpe.scala 176:32]
          Station8_4_4 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_4_4 <= _GEN_420;
        end
      end else begin
        Station8_4_4 <= _GEN_420;
      end
    end else begin
      Station8_4_4 <= _GEN_420;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2326 & _GEN_2273) begin // @[stationary_dpe.scala 176:32]
          Station8_4_5 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_4_5 <= _GEN_421;
        end
      end else begin
        Station8_4_5 <= _GEN_421;
      end
    end else begin
      Station8_4_5 <= _GEN_421;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2326 & _GEN_2275) begin // @[stationary_dpe.scala 176:32]
          Station8_4_6 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_4_6 <= _GEN_422;
        end
      end else begin
        Station8_4_6 <= _GEN_422;
      end
    end else begin
      Station8_4_6 <= _GEN_422;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2326 & _GEN_2277) begin // @[stationary_dpe.scala 176:32]
          Station8_4_7 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_4_7 <= _GEN_423;
        end
      end else begin
        Station8_4_7 <= _GEN_423;
      end
    end else begin
      Station8_4_7 <= _GEN_423;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2342 & _GEN_2279) begin // @[stationary_dpe.scala 176:32]
          Station8_5_0 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_5_0 <= _GEN_424;
        end
      end else begin
        Station8_5_0 <= _GEN_424;
      end
    end else begin
      Station8_5_0 <= _GEN_424;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2342 & _GEN_2265) begin // @[stationary_dpe.scala 176:32]
          Station8_5_1 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_5_1 <= _GEN_425;
        end
      end else begin
        Station8_5_1 <= _GEN_425;
      end
    end else begin
      Station8_5_1 <= _GEN_425;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2342 & _GEN_2267) begin // @[stationary_dpe.scala 176:32]
          Station8_5_2 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_5_2 <= _GEN_426;
        end
      end else begin
        Station8_5_2 <= _GEN_426;
      end
    end else begin
      Station8_5_2 <= _GEN_426;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2342 & _GEN_2269) begin // @[stationary_dpe.scala 176:32]
          Station8_5_3 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_5_3 <= _GEN_427;
        end
      end else begin
        Station8_5_3 <= _GEN_427;
      end
    end else begin
      Station8_5_3 <= _GEN_427;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2342 & _GEN_2271) begin // @[stationary_dpe.scala 176:32]
          Station8_5_4 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_5_4 <= _GEN_428;
        end
      end else begin
        Station8_5_4 <= _GEN_428;
      end
    end else begin
      Station8_5_4 <= _GEN_428;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2342 & _GEN_2273) begin // @[stationary_dpe.scala 176:32]
          Station8_5_5 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_5_5 <= _GEN_429;
        end
      end else begin
        Station8_5_5 <= _GEN_429;
      end
    end else begin
      Station8_5_5 <= _GEN_429;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2342 & _GEN_2275) begin // @[stationary_dpe.scala 176:32]
          Station8_5_6 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_5_6 <= _GEN_430;
        end
      end else begin
        Station8_5_6 <= _GEN_430;
      end
    end else begin
      Station8_5_6 <= _GEN_430;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2342 & _GEN_2277) begin // @[stationary_dpe.scala 176:32]
          Station8_5_7 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_5_7 <= _GEN_431;
        end
      end else begin
        Station8_5_7 <= _GEN_431;
      end
    end else begin
      Station8_5_7 <= _GEN_431;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2358 & _GEN_2279) begin // @[stationary_dpe.scala 176:32]
          Station8_6_0 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_6_0 <= _GEN_432;
        end
      end else begin
        Station8_6_0 <= _GEN_432;
      end
    end else begin
      Station8_6_0 <= _GEN_432;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2358 & _GEN_2265) begin // @[stationary_dpe.scala 176:32]
          Station8_6_1 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_6_1 <= _GEN_433;
        end
      end else begin
        Station8_6_1 <= _GEN_433;
      end
    end else begin
      Station8_6_1 <= _GEN_433;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2358 & _GEN_2267) begin // @[stationary_dpe.scala 176:32]
          Station8_6_2 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_6_2 <= _GEN_434;
        end
      end else begin
        Station8_6_2 <= _GEN_434;
      end
    end else begin
      Station8_6_2 <= _GEN_434;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2358 & _GEN_2269) begin // @[stationary_dpe.scala 176:32]
          Station8_6_3 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_6_3 <= _GEN_435;
        end
      end else begin
        Station8_6_3 <= _GEN_435;
      end
    end else begin
      Station8_6_3 <= _GEN_435;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2358 & _GEN_2271) begin // @[stationary_dpe.scala 176:32]
          Station8_6_4 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_6_4 <= _GEN_436;
        end
      end else begin
        Station8_6_4 <= _GEN_436;
      end
    end else begin
      Station8_6_4 <= _GEN_436;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2358 & _GEN_2273) begin // @[stationary_dpe.scala 176:32]
          Station8_6_5 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_6_5 <= _GEN_437;
        end
      end else begin
        Station8_6_5 <= _GEN_437;
      end
    end else begin
      Station8_6_5 <= _GEN_437;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2358 & _GEN_2275) begin // @[stationary_dpe.scala 176:32]
          Station8_6_6 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_6_6 <= _GEN_438;
        end
      end else begin
        Station8_6_6 <= _GEN_438;
      end
    end else begin
      Station8_6_6 <= _GEN_438;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2358 & _GEN_2277) begin // @[stationary_dpe.scala 176:32]
          Station8_6_7 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_6_7 <= _GEN_439;
        end
      end else begin
        Station8_6_7 <= _GEN_439;
      end
    end else begin
      Station8_6_7 <= _GEN_439;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2374 & _GEN_2279) begin // @[stationary_dpe.scala 176:32]
          Station8_7_0 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_7_0 <= _GEN_440;
        end
      end else begin
        Station8_7_0 <= _GEN_440;
      end
    end else begin
      Station8_7_0 <= _GEN_440;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2374 & _GEN_2265) begin // @[stationary_dpe.scala 176:32]
          Station8_7_1 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_7_1 <= _GEN_441;
        end
      end else begin
        Station8_7_1 <= _GEN_441;
      end
    end else begin
      Station8_7_1 <= _GEN_441;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2374 & _GEN_2267) begin // @[stationary_dpe.scala 176:32]
          Station8_7_2 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_7_2 <= _GEN_442;
        end
      end else begin
        Station8_7_2 <= _GEN_442;
      end
    end else begin
      Station8_7_2 <= _GEN_442;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2374 & _GEN_2269) begin // @[stationary_dpe.scala 176:32]
          Station8_7_3 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_7_3 <= _GEN_443;
        end
      end else begin
        Station8_7_3 <= _GEN_443;
      end
    end else begin
      Station8_7_3 <= _GEN_443;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2374 & _GEN_2271) begin // @[stationary_dpe.scala 176:32]
          Station8_7_4 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_7_4 <= _GEN_444;
        end
      end else begin
        Station8_7_4 <= _GEN_444;
      end
    end else begin
      Station8_7_4 <= _GEN_444;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2374 & _GEN_2273) begin // @[stationary_dpe.scala 176:32]
          Station8_7_5 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_7_5 <= _GEN_445;
        end
      end else begin
        Station8_7_5 <= _GEN_445;
      end
    end else begin
      Station8_7_5 <= _GEN_445;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2374 & _GEN_2275) begin // @[stationary_dpe.scala 176:32]
          Station8_7_6 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_7_6 <= _GEN_446;
        end
      end else begin
        Station8_7_6 <= _GEN_446;
      end
    end else begin
      Station8_7_6 <= _GEN_446;
    end
    if (~valid6) begin // @[stationary_dpe.scala 174:28]
      if (_GEN_2059 != 16'h0) begin // @[stationary_dpe.scala 175:39]
        if (_GEN_2374 & _GEN_2277) begin // @[stationary_dpe.scala 176:32]
          Station8_7_7 <= 16'h0; // @[stationary_dpe.scala 176:32]
        end else begin
          Station8_7_7 <= _GEN_447;
        end
      end else begin
        Station8_7_7 <= _GEN_447;
      end
    end else begin
      Station8_7_7 <= _GEN_447;
    end
    if (reset) begin // @[stationary_dpe.scala 79:20]
      i <= 32'h0; // @[stationary_dpe.scala 79:20]
    end else if (i < 32'h7 & j == 32'h7) begin // @[stationary_dpe.scala 222:74]
      i <= _i_T_1; // @[stationary_dpe.scala 223:11]
    end
    if (reset) begin // @[stationary_dpe.scala 80:20]
      j <= 32'h0; // @[stationary_dpe.scala 80:20]
    end else if (j < 32'h7 & i <= 32'h7) begin // @[stationary_dpe.scala 226:71]
      j <= _j_T_1; // @[stationary_dpe.scala 227:11]
    end else if (!(i == 32'h7 & _T_57)) begin // @[stationary_dpe.scala 229:81]
      j <= 32'h0; // @[stationary_dpe.scala 233:11]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  Station2_0_0 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  Station2_0_1 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  Station2_0_2 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  Station2_0_3 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  Station2_0_4 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  Station2_0_5 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  Station2_0_6 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  Station2_0_7 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  Station2_1_0 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  Station2_1_1 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  Station2_1_2 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  Station2_1_3 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  Station2_1_4 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  Station2_1_5 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  Station2_1_6 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  Station2_1_7 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  Station2_2_0 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  Station2_2_1 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  Station2_2_2 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  Station2_2_3 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  Station2_2_4 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  Station2_2_5 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  Station2_2_6 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  Station2_2_7 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  Station2_3_0 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  Station2_3_1 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  Station2_3_2 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  Station2_3_3 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  Station2_3_4 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  Station2_3_5 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  Station2_3_6 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  Station2_3_7 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  Station2_4_0 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  Station2_4_1 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  Station2_4_2 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  Station2_4_3 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  Station2_4_4 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  Station2_4_5 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  Station2_4_6 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  Station2_4_7 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  Station2_5_0 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  Station2_5_1 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  Station2_5_2 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  Station2_5_3 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  Station2_5_4 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  Station2_5_5 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  Station2_5_6 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  Station2_5_7 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  Station2_6_0 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  Station2_6_1 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  Station2_6_2 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  Station2_6_3 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  Station2_6_4 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  Station2_6_5 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  Station2_6_6 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  Station2_6_7 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  Station2_7_0 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  Station2_7_1 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  Station2_7_2 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  Station2_7_3 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  Station2_7_4 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  Station2_7_5 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  Station2_7_6 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  Station2_7_7 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  Station3_0_0 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  Station3_0_1 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  Station3_0_2 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  Station3_0_3 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  Station3_0_4 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  Station3_0_5 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  Station3_0_6 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  Station3_0_7 = _RAND_72[15:0];
  _RAND_73 = {1{`RANDOM}};
  Station3_1_0 = _RAND_73[15:0];
  _RAND_74 = {1{`RANDOM}};
  Station3_1_1 = _RAND_74[15:0];
  _RAND_75 = {1{`RANDOM}};
  Station3_1_2 = _RAND_75[15:0];
  _RAND_76 = {1{`RANDOM}};
  Station3_1_3 = _RAND_76[15:0];
  _RAND_77 = {1{`RANDOM}};
  Station3_1_4 = _RAND_77[15:0];
  _RAND_78 = {1{`RANDOM}};
  Station3_1_5 = _RAND_78[15:0];
  _RAND_79 = {1{`RANDOM}};
  Station3_1_6 = _RAND_79[15:0];
  _RAND_80 = {1{`RANDOM}};
  Station3_1_7 = _RAND_80[15:0];
  _RAND_81 = {1{`RANDOM}};
  Station3_2_0 = _RAND_81[15:0];
  _RAND_82 = {1{`RANDOM}};
  Station3_2_1 = _RAND_82[15:0];
  _RAND_83 = {1{`RANDOM}};
  Station3_2_2 = _RAND_83[15:0];
  _RAND_84 = {1{`RANDOM}};
  Station3_2_3 = _RAND_84[15:0];
  _RAND_85 = {1{`RANDOM}};
  Station3_2_4 = _RAND_85[15:0];
  _RAND_86 = {1{`RANDOM}};
  Station3_2_5 = _RAND_86[15:0];
  _RAND_87 = {1{`RANDOM}};
  Station3_2_6 = _RAND_87[15:0];
  _RAND_88 = {1{`RANDOM}};
  Station3_2_7 = _RAND_88[15:0];
  _RAND_89 = {1{`RANDOM}};
  Station3_3_0 = _RAND_89[15:0];
  _RAND_90 = {1{`RANDOM}};
  Station3_3_1 = _RAND_90[15:0];
  _RAND_91 = {1{`RANDOM}};
  Station3_3_2 = _RAND_91[15:0];
  _RAND_92 = {1{`RANDOM}};
  Station3_3_3 = _RAND_92[15:0];
  _RAND_93 = {1{`RANDOM}};
  Station3_3_4 = _RAND_93[15:0];
  _RAND_94 = {1{`RANDOM}};
  Station3_3_5 = _RAND_94[15:0];
  _RAND_95 = {1{`RANDOM}};
  Station3_3_6 = _RAND_95[15:0];
  _RAND_96 = {1{`RANDOM}};
  Station3_3_7 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  Station3_4_0 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  Station3_4_1 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  Station3_4_2 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  Station3_4_3 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  Station3_4_4 = _RAND_101[15:0];
  _RAND_102 = {1{`RANDOM}};
  Station3_4_5 = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  Station3_4_6 = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  Station3_4_7 = _RAND_104[15:0];
  _RAND_105 = {1{`RANDOM}};
  Station3_5_0 = _RAND_105[15:0];
  _RAND_106 = {1{`RANDOM}};
  Station3_5_1 = _RAND_106[15:0];
  _RAND_107 = {1{`RANDOM}};
  Station3_5_2 = _RAND_107[15:0];
  _RAND_108 = {1{`RANDOM}};
  Station3_5_3 = _RAND_108[15:0];
  _RAND_109 = {1{`RANDOM}};
  Station3_5_4 = _RAND_109[15:0];
  _RAND_110 = {1{`RANDOM}};
  Station3_5_5 = _RAND_110[15:0];
  _RAND_111 = {1{`RANDOM}};
  Station3_5_6 = _RAND_111[15:0];
  _RAND_112 = {1{`RANDOM}};
  Station3_5_7 = _RAND_112[15:0];
  _RAND_113 = {1{`RANDOM}};
  Station3_6_0 = _RAND_113[15:0];
  _RAND_114 = {1{`RANDOM}};
  Station3_6_1 = _RAND_114[15:0];
  _RAND_115 = {1{`RANDOM}};
  Station3_6_2 = _RAND_115[15:0];
  _RAND_116 = {1{`RANDOM}};
  Station3_6_3 = _RAND_116[15:0];
  _RAND_117 = {1{`RANDOM}};
  Station3_6_4 = _RAND_117[15:0];
  _RAND_118 = {1{`RANDOM}};
  Station3_6_5 = _RAND_118[15:0];
  _RAND_119 = {1{`RANDOM}};
  Station3_6_6 = _RAND_119[15:0];
  _RAND_120 = {1{`RANDOM}};
  Station3_6_7 = _RAND_120[15:0];
  _RAND_121 = {1{`RANDOM}};
  Station3_7_0 = _RAND_121[15:0];
  _RAND_122 = {1{`RANDOM}};
  Station3_7_1 = _RAND_122[15:0];
  _RAND_123 = {1{`RANDOM}};
  Station3_7_2 = _RAND_123[15:0];
  _RAND_124 = {1{`RANDOM}};
  Station3_7_3 = _RAND_124[15:0];
  _RAND_125 = {1{`RANDOM}};
  Station3_7_4 = _RAND_125[15:0];
  _RAND_126 = {1{`RANDOM}};
  Station3_7_5 = _RAND_126[15:0];
  _RAND_127 = {1{`RANDOM}};
  Station3_7_6 = _RAND_127[15:0];
  _RAND_128 = {1{`RANDOM}};
  Station3_7_7 = _RAND_128[15:0];
  _RAND_129 = {1{`RANDOM}};
  Station4_0_0 = _RAND_129[15:0];
  _RAND_130 = {1{`RANDOM}};
  Station4_0_1 = _RAND_130[15:0];
  _RAND_131 = {1{`RANDOM}};
  Station4_0_2 = _RAND_131[15:0];
  _RAND_132 = {1{`RANDOM}};
  Station4_0_3 = _RAND_132[15:0];
  _RAND_133 = {1{`RANDOM}};
  Station4_0_4 = _RAND_133[15:0];
  _RAND_134 = {1{`RANDOM}};
  Station4_0_5 = _RAND_134[15:0];
  _RAND_135 = {1{`RANDOM}};
  Station4_0_6 = _RAND_135[15:0];
  _RAND_136 = {1{`RANDOM}};
  Station4_0_7 = _RAND_136[15:0];
  _RAND_137 = {1{`RANDOM}};
  Station4_1_0 = _RAND_137[15:0];
  _RAND_138 = {1{`RANDOM}};
  Station4_1_1 = _RAND_138[15:0];
  _RAND_139 = {1{`RANDOM}};
  Station4_1_2 = _RAND_139[15:0];
  _RAND_140 = {1{`RANDOM}};
  Station4_1_3 = _RAND_140[15:0];
  _RAND_141 = {1{`RANDOM}};
  Station4_1_4 = _RAND_141[15:0];
  _RAND_142 = {1{`RANDOM}};
  Station4_1_5 = _RAND_142[15:0];
  _RAND_143 = {1{`RANDOM}};
  Station4_1_6 = _RAND_143[15:0];
  _RAND_144 = {1{`RANDOM}};
  Station4_1_7 = _RAND_144[15:0];
  _RAND_145 = {1{`RANDOM}};
  Station4_2_0 = _RAND_145[15:0];
  _RAND_146 = {1{`RANDOM}};
  Station4_2_1 = _RAND_146[15:0];
  _RAND_147 = {1{`RANDOM}};
  Station4_2_2 = _RAND_147[15:0];
  _RAND_148 = {1{`RANDOM}};
  Station4_2_3 = _RAND_148[15:0];
  _RAND_149 = {1{`RANDOM}};
  Station4_2_4 = _RAND_149[15:0];
  _RAND_150 = {1{`RANDOM}};
  Station4_2_5 = _RAND_150[15:0];
  _RAND_151 = {1{`RANDOM}};
  Station4_2_6 = _RAND_151[15:0];
  _RAND_152 = {1{`RANDOM}};
  Station4_2_7 = _RAND_152[15:0];
  _RAND_153 = {1{`RANDOM}};
  Station4_3_0 = _RAND_153[15:0];
  _RAND_154 = {1{`RANDOM}};
  Station4_3_1 = _RAND_154[15:0];
  _RAND_155 = {1{`RANDOM}};
  Station4_3_2 = _RAND_155[15:0];
  _RAND_156 = {1{`RANDOM}};
  Station4_3_3 = _RAND_156[15:0];
  _RAND_157 = {1{`RANDOM}};
  Station4_3_4 = _RAND_157[15:0];
  _RAND_158 = {1{`RANDOM}};
  Station4_3_5 = _RAND_158[15:0];
  _RAND_159 = {1{`RANDOM}};
  Station4_3_6 = _RAND_159[15:0];
  _RAND_160 = {1{`RANDOM}};
  Station4_3_7 = _RAND_160[15:0];
  _RAND_161 = {1{`RANDOM}};
  Station4_4_0 = _RAND_161[15:0];
  _RAND_162 = {1{`RANDOM}};
  Station4_4_1 = _RAND_162[15:0];
  _RAND_163 = {1{`RANDOM}};
  Station4_4_2 = _RAND_163[15:0];
  _RAND_164 = {1{`RANDOM}};
  Station4_4_3 = _RAND_164[15:0];
  _RAND_165 = {1{`RANDOM}};
  Station4_4_4 = _RAND_165[15:0];
  _RAND_166 = {1{`RANDOM}};
  Station4_4_5 = _RAND_166[15:0];
  _RAND_167 = {1{`RANDOM}};
  Station4_4_6 = _RAND_167[15:0];
  _RAND_168 = {1{`RANDOM}};
  Station4_4_7 = _RAND_168[15:0];
  _RAND_169 = {1{`RANDOM}};
  Station4_5_0 = _RAND_169[15:0];
  _RAND_170 = {1{`RANDOM}};
  Station4_5_1 = _RAND_170[15:0];
  _RAND_171 = {1{`RANDOM}};
  Station4_5_2 = _RAND_171[15:0];
  _RAND_172 = {1{`RANDOM}};
  Station4_5_3 = _RAND_172[15:0];
  _RAND_173 = {1{`RANDOM}};
  Station4_5_4 = _RAND_173[15:0];
  _RAND_174 = {1{`RANDOM}};
  Station4_5_5 = _RAND_174[15:0];
  _RAND_175 = {1{`RANDOM}};
  Station4_5_6 = _RAND_175[15:0];
  _RAND_176 = {1{`RANDOM}};
  Station4_5_7 = _RAND_176[15:0];
  _RAND_177 = {1{`RANDOM}};
  Station4_6_0 = _RAND_177[15:0];
  _RAND_178 = {1{`RANDOM}};
  Station4_6_1 = _RAND_178[15:0];
  _RAND_179 = {1{`RANDOM}};
  Station4_6_2 = _RAND_179[15:0];
  _RAND_180 = {1{`RANDOM}};
  Station4_6_3 = _RAND_180[15:0];
  _RAND_181 = {1{`RANDOM}};
  Station4_6_4 = _RAND_181[15:0];
  _RAND_182 = {1{`RANDOM}};
  Station4_6_5 = _RAND_182[15:0];
  _RAND_183 = {1{`RANDOM}};
  Station4_6_6 = _RAND_183[15:0];
  _RAND_184 = {1{`RANDOM}};
  Station4_6_7 = _RAND_184[15:0];
  _RAND_185 = {1{`RANDOM}};
  Station4_7_0 = _RAND_185[15:0];
  _RAND_186 = {1{`RANDOM}};
  Station4_7_1 = _RAND_186[15:0];
  _RAND_187 = {1{`RANDOM}};
  Station4_7_2 = _RAND_187[15:0];
  _RAND_188 = {1{`RANDOM}};
  Station4_7_3 = _RAND_188[15:0];
  _RAND_189 = {1{`RANDOM}};
  Station4_7_4 = _RAND_189[15:0];
  _RAND_190 = {1{`RANDOM}};
  Station4_7_5 = _RAND_190[15:0];
  _RAND_191 = {1{`RANDOM}};
  Station4_7_6 = _RAND_191[15:0];
  _RAND_192 = {1{`RANDOM}};
  Station4_7_7 = _RAND_192[15:0];
  _RAND_193 = {1{`RANDOM}};
  Station5_0_0 = _RAND_193[15:0];
  _RAND_194 = {1{`RANDOM}};
  Station5_0_1 = _RAND_194[15:0];
  _RAND_195 = {1{`RANDOM}};
  Station5_0_2 = _RAND_195[15:0];
  _RAND_196 = {1{`RANDOM}};
  Station5_0_3 = _RAND_196[15:0];
  _RAND_197 = {1{`RANDOM}};
  Station5_0_4 = _RAND_197[15:0];
  _RAND_198 = {1{`RANDOM}};
  Station5_0_5 = _RAND_198[15:0];
  _RAND_199 = {1{`RANDOM}};
  Station5_0_6 = _RAND_199[15:0];
  _RAND_200 = {1{`RANDOM}};
  Station5_0_7 = _RAND_200[15:0];
  _RAND_201 = {1{`RANDOM}};
  Station5_1_0 = _RAND_201[15:0];
  _RAND_202 = {1{`RANDOM}};
  Station5_1_1 = _RAND_202[15:0];
  _RAND_203 = {1{`RANDOM}};
  Station5_1_2 = _RAND_203[15:0];
  _RAND_204 = {1{`RANDOM}};
  Station5_1_3 = _RAND_204[15:0];
  _RAND_205 = {1{`RANDOM}};
  Station5_1_4 = _RAND_205[15:0];
  _RAND_206 = {1{`RANDOM}};
  Station5_1_5 = _RAND_206[15:0];
  _RAND_207 = {1{`RANDOM}};
  Station5_1_6 = _RAND_207[15:0];
  _RAND_208 = {1{`RANDOM}};
  Station5_1_7 = _RAND_208[15:0];
  _RAND_209 = {1{`RANDOM}};
  Station5_2_0 = _RAND_209[15:0];
  _RAND_210 = {1{`RANDOM}};
  Station5_2_1 = _RAND_210[15:0];
  _RAND_211 = {1{`RANDOM}};
  Station5_2_2 = _RAND_211[15:0];
  _RAND_212 = {1{`RANDOM}};
  Station5_2_3 = _RAND_212[15:0];
  _RAND_213 = {1{`RANDOM}};
  Station5_2_4 = _RAND_213[15:0];
  _RAND_214 = {1{`RANDOM}};
  Station5_2_5 = _RAND_214[15:0];
  _RAND_215 = {1{`RANDOM}};
  Station5_2_6 = _RAND_215[15:0];
  _RAND_216 = {1{`RANDOM}};
  Station5_2_7 = _RAND_216[15:0];
  _RAND_217 = {1{`RANDOM}};
  Station5_3_0 = _RAND_217[15:0];
  _RAND_218 = {1{`RANDOM}};
  Station5_3_1 = _RAND_218[15:0];
  _RAND_219 = {1{`RANDOM}};
  Station5_3_2 = _RAND_219[15:0];
  _RAND_220 = {1{`RANDOM}};
  Station5_3_3 = _RAND_220[15:0];
  _RAND_221 = {1{`RANDOM}};
  Station5_3_4 = _RAND_221[15:0];
  _RAND_222 = {1{`RANDOM}};
  Station5_3_5 = _RAND_222[15:0];
  _RAND_223 = {1{`RANDOM}};
  Station5_3_6 = _RAND_223[15:0];
  _RAND_224 = {1{`RANDOM}};
  Station5_3_7 = _RAND_224[15:0];
  _RAND_225 = {1{`RANDOM}};
  Station5_4_0 = _RAND_225[15:0];
  _RAND_226 = {1{`RANDOM}};
  Station5_4_1 = _RAND_226[15:0];
  _RAND_227 = {1{`RANDOM}};
  Station5_4_2 = _RAND_227[15:0];
  _RAND_228 = {1{`RANDOM}};
  Station5_4_3 = _RAND_228[15:0];
  _RAND_229 = {1{`RANDOM}};
  Station5_4_4 = _RAND_229[15:0];
  _RAND_230 = {1{`RANDOM}};
  Station5_4_5 = _RAND_230[15:0];
  _RAND_231 = {1{`RANDOM}};
  Station5_4_6 = _RAND_231[15:0];
  _RAND_232 = {1{`RANDOM}};
  Station5_4_7 = _RAND_232[15:0];
  _RAND_233 = {1{`RANDOM}};
  Station5_5_0 = _RAND_233[15:0];
  _RAND_234 = {1{`RANDOM}};
  Station5_5_1 = _RAND_234[15:0];
  _RAND_235 = {1{`RANDOM}};
  Station5_5_2 = _RAND_235[15:0];
  _RAND_236 = {1{`RANDOM}};
  Station5_5_3 = _RAND_236[15:0];
  _RAND_237 = {1{`RANDOM}};
  Station5_5_4 = _RAND_237[15:0];
  _RAND_238 = {1{`RANDOM}};
  Station5_5_5 = _RAND_238[15:0];
  _RAND_239 = {1{`RANDOM}};
  Station5_5_6 = _RAND_239[15:0];
  _RAND_240 = {1{`RANDOM}};
  Station5_5_7 = _RAND_240[15:0];
  _RAND_241 = {1{`RANDOM}};
  Station5_6_0 = _RAND_241[15:0];
  _RAND_242 = {1{`RANDOM}};
  Station5_6_1 = _RAND_242[15:0];
  _RAND_243 = {1{`RANDOM}};
  Station5_6_2 = _RAND_243[15:0];
  _RAND_244 = {1{`RANDOM}};
  Station5_6_3 = _RAND_244[15:0];
  _RAND_245 = {1{`RANDOM}};
  Station5_6_4 = _RAND_245[15:0];
  _RAND_246 = {1{`RANDOM}};
  Station5_6_5 = _RAND_246[15:0];
  _RAND_247 = {1{`RANDOM}};
  Station5_6_6 = _RAND_247[15:0];
  _RAND_248 = {1{`RANDOM}};
  Station5_6_7 = _RAND_248[15:0];
  _RAND_249 = {1{`RANDOM}};
  Station5_7_0 = _RAND_249[15:0];
  _RAND_250 = {1{`RANDOM}};
  Station5_7_1 = _RAND_250[15:0];
  _RAND_251 = {1{`RANDOM}};
  Station5_7_2 = _RAND_251[15:0];
  _RAND_252 = {1{`RANDOM}};
  Station5_7_3 = _RAND_252[15:0];
  _RAND_253 = {1{`RANDOM}};
  Station5_7_4 = _RAND_253[15:0];
  _RAND_254 = {1{`RANDOM}};
  Station5_7_5 = _RAND_254[15:0];
  _RAND_255 = {1{`RANDOM}};
  Station5_7_6 = _RAND_255[15:0];
  _RAND_256 = {1{`RANDOM}};
  Station5_7_7 = _RAND_256[15:0];
  _RAND_257 = {1{`RANDOM}};
  Station6_0_0 = _RAND_257[15:0];
  _RAND_258 = {1{`RANDOM}};
  Station6_0_1 = _RAND_258[15:0];
  _RAND_259 = {1{`RANDOM}};
  Station6_0_2 = _RAND_259[15:0];
  _RAND_260 = {1{`RANDOM}};
  Station6_0_3 = _RAND_260[15:0];
  _RAND_261 = {1{`RANDOM}};
  Station6_0_4 = _RAND_261[15:0];
  _RAND_262 = {1{`RANDOM}};
  Station6_0_5 = _RAND_262[15:0];
  _RAND_263 = {1{`RANDOM}};
  Station6_0_6 = _RAND_263[15:0];
  _RAND_264 = {1{`RANDOM}};
  Station6_0_7 = _RAND_264[15:0];
  _RAND_265 = {1{`RANDOM}};
  Station6_1_0 = _RAND_265[15:0];
  _RAND_266 = {1{`RANDOM}};
  Station6_1_1 = _RAND_266[15:0];
  _RAND_267 = {1{`RANDOM}};
  Station6_1_2 = _RAND_267[15:0];
  _RAND_268 = {1{`RANDOM}};
  Station6_1_3 = _RAND_268[15:0];
  _RAND_269 = {1{`RANDOM}};
  Station6_1_4 = _RAND_269[15:0];
  _RAND_270 = {1{`RANDOM}};
  Station6_1_5 = _RAND_270[15:0];
  _RAND_271 = {1{`RANDOM}};
  Station6_1_6 = _RAND_271[15:0];
  _RAND_272 = {1{`RANDOM}};
  Station6_1_7 = _RAND_272[15:0];
  _RAND_273 = {1{`RANDOM}};
  Station6_2_0 = _RAND_273[15:0];
  _RAND_274 = {1{`RANDOM}};
  Station6_2_1 = _RAND_274[15:0];
  _RAND_275 = {1{`RANDOM}};
  Station6_2_2 = _RAND_275[15:0];
  _RAND_276 = {1{`RANDOM}};
  Station6_2_3 = _RAND_276[15:0];
  _RAND_277 = {1{`RANDOM}};
  Station6_2_4 = _RAND_277[15:0];
  _RAND_278 = {1{`RANDOM}};
  Station6_2_5 = _RAND_278[15:0];
  _RAND_279 = {1{`RANDOM}};
  Station6_2_6 = _RAND_279[15:0];
  _RAND_280 = {1{`RANDOM}};
  Station6_2_7 = _RAND_280[15:0];
  _RAND_281 = {1{`RANDOM}};
  Station6_3_0 = _RAND_281[15:0];
  _RAND_282 = {1{`RANDOM}};
  Station6_3_1 = _RAND_282[15:0];
  _RAND_283 = {1{`RANDOM}};
  Station6_3_2 = _RAND_283[15:0];
  _RAND_284 = {1{`RANDOM}};
  Station6_3_3 = _RAND_284[15:0];
  _RAND_285 = {1{`RANDOM}};
  Station6_3_4 = _RAND_285[15:0];
  _RAND_286 = {1{`RANDOM}};
  Station6_3_5 = _RAND_286[15:0];
  _RAND_287 = {1{`RANDOM}};
  Station6_3_6 = _RAND_287[15:0];
  _RAND_288 = {1{`RANDOM}};
  Station6_3_7 = _RAND_288[15:0];
  _RAND_289 = {1{`RANDOM}};
  Station6_4_0 = _RAND_289[15:0];
  _RAND_290 = {1{`RANDOM}};
  Station6_4_1 = _RAND_290[15:0];
  _RAND_291 = {1{`RANDOM}};
  Station6_4_2 = _RAND_291[15:0];
  _RAND_292 = {1{`RANDOM}};
  Station6_4_3 = _RAND_292[15:0];
  _RAND_293 = {1{`RANDOM}};
  Station6_4_4 = _RAND_293[15:0];
  _RAND_294 = {1{`RANDOM}};
  Station6_4_5 = _RAND_294[15:0];
  _RAND_295 = {1{`RANDOM}};
  Station6_4_6 = _RAND_295[15:0];
  _RAND_296 = {1{`RANDOM}};
  Station6_4_7 = _RAND_296[15:0];
  _RAND_297 = {1{`RANDOM}};
  Station6_5_0 = _RAND_297[15:0];
  _RAND_298 = {1{`RANDOM}};
  Station6_5_1 = _RAND_298[15:0];
  _RAND_299 = {1{`RANDOM}};
  Station6_5_2 = _RAND_299[15:0];
  _RAND_300 = {1{`RANDOM}};
  Station6_5_3 = _RAND_300[15:0];
  _RAND_301 = {1{`RANDOM}};
  Station6_5_4 = _RAND_301[15:0];
  _RAND_302 = {1{`RANDOM}};
  Station6_5_5 = _RAND_302[15:0];
  _RAND_303 = {1{`RANDOM}};
  Station6_5_6 = _RAND_303[15:0];
  _RAND_304 = {1{`RANDOM}};
  Station6_5_7 = _RAND_304[15:0];
  _RAND_305 = {1{`RANDOM}};
  Station6_6_0 = _RAND_305[15:0];
  _RAND_306 = {1{`RANDOM}};
  Station6_6_1 = _RAND_306[15:0];
  _RAND_307 = {1{`RANDOM}};
  Station6_6_2 = _RAND_307[15:0];
  _RAND_308 = {1{`RANDOM}};
  Station6_6_3 = _RAND_308[15:0];
  _RAND_309 = {1{`RANDOM}};
  Station6_6_4 = _RAND_309[15:0];
  _RAND_310 = {1{`RANDOM}};
  Station6_6_5 = _RAND_310[15:0];
  _RAND_311 = {1{`RANDOM}};
  Station6_6_6 = _RAND_311[15:0];
  _RAND_312 = {1{`RANDOM}};
  Station6_6_7 = _RAND_312[15:0];
  _RAND_313 = {1{`RANDOM}};
  Station6_7_0 = _RAND_313[15:0];
  _RAND_314 = {1{`RANDOM}};
  Station6_7_1 = _RAND_314[15:0];
  _RAND_315 = {1{`RANDOM}};
  Station6_7_2 = _RAND_315[15:0];
  _RAND_316 = {1{`RANDOM}};
  Station6_7_3 = _RAND_316[15:0];
  _RAND_317 = {1{`RANDOM}};
  Station6_7_4 = _RAND_317[15:0];
  _RAND_318 = {1{`RANDOM}};
  Station6_7_5 = _RAND_318[15:0];
  _RAND_319 = {1{`RANDOM}};
  Station6_7_6 = _RAND_319[15:0];
  _RAND_320 = {1{`RANDOM}};
  Station6_7_7 = _RAND_320[15:0];
  _RAND_321 = {1{`RANDOM}};
  Station7_0_0 = _RAND_321[15:0];
  _RAND_322 = {1{`RANDOM}};
  Station7_0_1 = _RAND_322[15:0];
  _RAND_323 = {1{`RANDOM}};
  Station7_0_2 = _RAND_323[15:0];
  _RAND_324 = {1{`RANDOM}};
  Station7_0_3 = _RAND_324[15:0];
  _RAND_325 = {1{`RANDOM}};
  Station7_0_4 = _RAND_325[15:0];
  _RAND_326 = {1{`RANDOM}};
  Station7_0_5 = _RAND_326[15:0];
  _RAND_327 = {1{`RANDOM}};
  Station7_0_6 = _RAND_327[15:0];
  _RAND_328 = {1{`RANDOM}};
  Station7_0_7 = _RAND_328[15:0];
  _RAND_329 = {1{`RANDOM}};
  Station7_1_0 = _RAND_329[15:0];
  _RAND_330 = {1{`RANDOM}};
  Station7_1_1 = _RAND_330[15:0];
  _RAND_331 = {1{`RANDOM}};
  Station7_1_2 = _RAND_331[15:0];
  _RAND_332 = {1{`RANDOM}};
  Station7_1_3 = _RAND_332[15:0];
  _RAND_333 = {1{`RANDOM}};
  Station7_1_4 = _RAND_333[15:0];
  _RAND_334 = {1{`RANDOM}};
  Station7_1_5 = _RAND_334[15:0];
  _RAND_335 = {1{`RANDOM}};
  Station7_1_6 = _RAND_335[15:0];
  _RAND_336 = {1{`RANDOM}};
  Station7_1_7 = _RAND_336[15:0];
  _RAND_337 = {1{`RANDOM}};
  Station7_2_0 = _RAND_337[15:0];
  _RAND_338 = {1{`RANDOM}};
  Station7_2_1 = _RAND_338[15:0];
  _RAND_339 = {1{`RANDOM}};
  Station7_2_2 = _RAND_339[15:0];
  _RAND_340 = {1{`RANDOM}};
  Station7_2_3 = _RAND_340[15:0];
  _RAND_341 = {1{`RANDOM}};
  Station7_2_4 = _RAND_341[15:0];
  _RAND_342 = {1{`RANDOM}};
  Station7_2_5 = _RAND_342[15:0];
  _RAND_343 = {1{`RANDOM}};
  Station7_2_6 = _RAND_343[15:0];
  _RAND_344 = {1{`RANDOM}};
  Station7_2_7 = _RAND_344[15:0];
  _RAND_345 = {1{`RANDOM}};
  Station7_3_0 = _RAND_345[15:0];
  _RAND_346 = {1{`RANDOM}};
  Station7_3_1 = _RAND_346[15:0];
  _RAND_347 = {1{`RANDOM}};
  Station7_3_2 = _RAND_347[15:0];
  _RAND_348 = {1{`RANDOM}};
  Station7_3_3 = _RAND_348[15:0];
  _RAND_349 = {1{`RANDOM}};
  Station7_3_4 = _RAND_349[15:0];
  _RAND_350 = {1{`RANDOM}};
  Station7_3_5 = _RAND_350[15:0];
  _RAND_351 = {1{`RANDOM}};
  Station7_3_6 = _RAND_351[15:0];
  _RAND_352 = {1{`RANDOM}};
  Station7_3_7 = _RAND_352[15:0];
  _RAND_353 = {1{`RANDOM}};
  Station7_4_0 = _RAND_353[15:0];
  _RAND_354 = {1{`RANDOM}};
  Station7_4_1 = _RAND_354[15:0];
  _RAND_355 = {1{`RANDOM}};
  Station7_4_2 = _RAND_355[15:0];
  _RAND_356 = {1{`RANDOM}};
  Station7_4_3 = _RAND_356[15:0];
  _RAND_357 = {1{`RANDOM}};
  Station7_4_4 = _RAND_357[15:0];
  _RAND_358 = {1{`RANDOM}};
  Station7_4_5 = _RAND_358[15:0];
  _RAND_359 = {1{`RANDOM}};
  Station7_4_6 = _RAND_359[15:0];
  _RAND_360 = {1{`RANDOM}};
  Station7_4_7 = _RAND_360[15:0];
  _RAND_361 = {1{`RANDOM}};
  Station7_5_0 = _RAND_361[15:0];
  _RAND_362 = {1{`RANDOM}};
  Station7_5_1 = _RAND_362[15:0];
  _RAND_363 = {1{`RANDOM}};
  Station7_5_2 = _RAND_363[15:0];
  _RAND_364 = {1{`RANDOM}};
  Station7_5_3 = _RAND_364[15:0];
  _RAND_365 = {1{`RANDOM}};
  Station7_5_4 = _RAND_365[15:0];
  _RAND_366 = {1{`RANDOM}};
  Station7_5_5 = _RAND_366[15:0];
  _RAND_367 = {1{`RANDOM}};
  Station7_5_6 = _RAND_367[15:0];
  _RAND_368 = {1{`RANDOM}};
  Station7_5_7 = _RAND_368[15:0];
  _RAND_369 = {1{`RANDOM}};
  Station7_6_0 = _RAND_369[15:0];
  _RAND_370 = {1{`RANDOM}};
  Station7_6_1 = _RAND_370[15:0];
  _RAND_371 = {1{`RANDOM}};
  Station7_6_2 = _RAND_371[15:0];
  _RAND_372 = {1{`RANDOM}};
  Station7_6_3 = _RAND_372[15:0];
  _RAND_373 = {1{`RANDOM}};
  Station7_6_4 = _RAND_373[15:0];
  _RAND_374 = {1{`RANDOM}};
  Station7_6_5 = _RAND_374[15:0];
  _RAND_375 = {1{`RANDOM}};
  Station7_6_6 = _RAND_375[15:0];
  _RAND_376 = {1{`RANDOM}};
  Station7_6_7 = _RAND_376[15:0];
  _RAND_377 = {1{`RANDOM}};
  Station7_7_0 = _RAND_377[15:0];
  _RAND_378 = {1{`RANDOM}};
  Station7_7_1 = _RAND_378[15:0];
  _RAND_379 = {1{`RANDOM}};
  Station7_7_2 = _RAND_379[15:0];
  _RAND_380 = {1{`RANDOM}};
  Station7_7_3 = _RAND_380[15:0];
  _RAND_381 = {1{`RANDOM}};
  Station7_7_4 = _RAND_381[15:0];
  _RAND_382 = {1{`RANDOM}};
  Station7_7_5 = _RAND_382[15:0];
  _RAND_383 = {1{`RANDOM}};
  Station7_7_6 = _RAND_383[15:0];
  _RAND_384 = {1{`RANDOM}};
  Station7_7_7 = _RAND_384[15:0];
  _RAND_385 = {1{`RANDOM}};
  Station8_0_0 = _RAND_385[15:0];
  _RAND_386 = {1{`RANDOM}};
  Station8_0_1 = _RAND_386[15:0];
  _RAND_387 = {1{`RANDOM}};
  Station8_0_2 = _RAND_387[15:0];
  _RAND_388 = {1{`RANDOM}};
  Station8_0_3 = _RAND_388[15:0];
  _RAND_389 = {1{`RANDOM}};
  Station8_0_4 = _RAND_389[15:0];
  _RAND_390 = {1{`RANDOM}};
  Station8_0_5 = _RAND_390[15:0];
  _RAND_391 = {1{`RANDOM}};
  Station8_0_6 = _RAND_391[15:0];
  _RAND_392 = {1{`RANDOM}};
  Station8_0_7 = _RAND_392[15:0];
  _RAND_393 = {1{`RANDOM}};
  Station8_1_0 = _RAND_393[15:0];
  _RAND_394 = {1{`RANDOM}};
  Station8_1_1 = _RAND_394[15:0];
  _RAND_395 = {1{`RANDOM}};
  Station8_1_2 = _RAND_395[15:0];
  _RAND_396 = {1{`RANDOM}};
  Station8_1_3 = _RAND_396[15:0];
  _RAND_397 = {1{`RANDOM}};
  Station8_1_4 = _RAND_397[15:0];
  _RAND_398 = {1{`RANDOM}};
  Station8_1_5 = _RAND_398[15:0];
  _RAND_399 = {1{`RANDOM}};
  Station8_1_6 = _RAND_399[15:0];
  _RAND_400 = {1{`RANDOM}};
  Station8_1_7 = _RAND_400[15:0];
  _RAND_401 = {1{`RANDOM}};
  Station8_2_0 = _RAND_401[15:0];
  _RAND_402 = {1{`RANDOM}};
  Station8_2_1 = _RAND_402[15:0];
  _RAND_403 = {1{`RANDOM}};
  Station8_2_2 = _RAND_403[15:0];
  _RAND_404 = {1{`RANDOM}};
  Station8_2_3 = _RAND_404[15:0];
  _RAND_405 = {1{`RANDOM}};
  Station8_2_4 = _RAND_405[15:0];
  _RAND_406 = {1{`RANDOM}};
  Station8_2_5 = _RAND_406[15:0];
  _RAND_407 = {1{`RANDOM}};
  Station8_2_6 = _RAND_407[15:0];
  _RAND_408 = {1{`RANDOM}};
  Station8_2_7 = _RAND_408[15:0];
  _RAND_409 = {1{`RANDOM}};
  Station8_3_0 = _RAND_409[15:0];
  _RAND_410 = {1{`RANDOM}};
  Station8_3_1 = _RAND_410[15:0];
  _RAND_411 = {1{`RANDOM}};
  Station8_3_2 = _RAND_411[15:0];
  _RAND_412 = {1{`RANDOM}};
  Station8_3_3 = _RAND_412[15:0];
  _RAND_413 = {1{`RANDOM}};
  Station8_3_4 = _RAND_413[15:0];
  _RAND_414 = {1{`RANDOM}};
  Station8_3_5 = _RAND_414[15:0];
  _RAND_415 = {1{`RANDOM}};
  Station8_3_6 = _RAND_415[15:0];
  _RAND_416 = {1{`RANDOM}};
  Station8_3_7 = _RAND_416[15:0];
  _RAND_417 = {1{`RANDOM}};
  Station8_4_0 = _RAND_417[15:0];
  _RAND_418 = {1{`RANDOM}};
  Station8_4_1 = _RAND_418[15:0];
  _RAND_419 = {1{`RANDOM}};
  Station8_4_2 = _RAND_419[15:0];
  _RAND_420 = {1{`RANDOM}};
  Station8_4_3 = _RAND_420[15:0];
  _RAND_421 = {1{`RANDOM}};
  Station8_4_4 = _RAND_421[15:0];
  _RAND_422 = {1{`RANDOM}};
  Station8_4_5 = _RAND_422[15:0];
  _RAND_423 = {1{`RANDOM}};
  Station8_4_6 = _RAND_423[15:0];
  _RAND_424 = {1{`RANDOM}};
  Station8_4_7 = _RAND_424[15:0];
  _RAND_425 = {1{`RANDOM}};
  Station8_5_0 = _RAND_425[15:0];
  _RAND_426 = {1{`RANDOM}};
  Station8_5_1 = _RAND_426[15:0];
  _RAND_427 = {1{`RANDOM}};
  Station8_5_2 = _RAND_427[15:0];
  _RAND_428 = {1{`RANDOM}};
  Station8_5_3 = _RAND_428[15:0];
  _RAND_429 = {1{`RANDOM}};
  Station8_5_4 = _RAND_429[15:0];
  _RAND_430 = {1{`RANDOM}};
  Station8_5_5 = _RAND_430[15:0];
  _RAND_431 = {1{`RANDOM}};
  Station8_5_6 = _RAND_431[15:0];
  _RAND_432 = {1{`RANDOM}};
  Station8_5_7 = _RAND_432[15:0];
  _RAND_433 = {1{`RANDOM}};
  Station8_6_0 = _RAND_433[15:0];
  _RAND_434 = {1{`RANDOM}};
  Station8_6_1 = _RAND_434[15:0];
  _RAND_435 = {1{`RANDOM}};
  Station8_6_2 = _RAND_435[15:0];
  _RAND_436 = {1{`RANDOM}};
  Station8_6_3 = _RAND_436[15:0];
  _RAND_437 = {1{`RANDOM}};
  Station8_6_4 = _RAND_437[15:0];
  _RAND_438 = {1{`RANDOM}};
  Station8_6_5 = _RAND_438[15:0];
  _RAND_439 = {1{`RANDOM}};
  Station8_6_6 = _RAND_439[15:0];
  _RAND_440 = {1{`RANDOM}};
  Station8_6_7 = _RAND_440[15:0];
  _RAND_441 = {1{`RANDOM}};
  Station8_7_0 = _RAND_441[15:0];
  _RAND_442 = {1{`RANDOM}};
  Station8_7_1 = _RAND_442[15:0];
  _RAND_443 = {1{`RANDOM}};
  Station8_7_2 = _RAND_443[15:0];
  _RAND_444 = {1{`RANDOM}};
  Station8_7_3 = _RAND_444[15:0];
  _RAND_445 = {1{`RANDOM}};
  Station8_7_4 = _RAND_445[15:0];
  _RAND_446 = {1{`RANDOM}};
  Station8_7_5 = _RAND_446[15:0];
  _RAND_447 = {1{`RANDOM}};
  Station8_7_6 = _RAND_447[15:0];
  _RAND_448 = {1{`RANDOM}};
  Station8_7_7 = _RAND_448[15:0];
  _RAND_449 = {1{`RANDOM}};
  i = _RAND_449[31:0];
  _RAND_450 = {1{`RANDOM}};
  j = _RAND_450[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ivncontrol4(
  input         clock,
  input         reset,
  input  [15:0] io_Stationary_matrix_0_0,
  input  [15:0] io_Stationary_matrix_0_1,
  input  [15:0] io_Stationary_matrix_0_2,
  input  [15:0] io_Stationary_matrix_0_3,
  input  [15:0] io_Stationary_matrix_0_4,
  input  [15:0] io_Stationary_matrix_0_5,
  input  [15:0] io_Stationary_matrix_0_6,
  input  [15:0] io_Stationary_matrix_0_7,
  input  [15:0] io_Stationary_matrix_1_0,
  input  [15:0] io_Stationary_matrix_1_1,
  input  [15:0] io_Stationary_matrix_1_2,
  input  [15:0] io_Stationary_matrix_1_3,
  input  [15:0] io_Stationary_matrix_1_4,
  input  [15:0] io_Stationary_matrix_1_5,
  input  [15:0] io_Stationary_matrix_1_6,
  input  [15:0] io_Stationary_matrix_1_7,
  input  [15:0] io_Stationary_matrix_2_0,
  input  [15:0] io_Stationary_matrix_2_1,
  input  [15:0] io_Stationary_matrix_2_2,
  input  [15:0] io_Stationary_matrix_2_3,
  input  [15:0] io_Stationary_matrix_2_4,
  input  [15:0] io_Stationary_matrix_2_5,
  input  [15:0] io_Stationary_matrix_2_6,
  input  [15:0] io_Stationary_matrix_2_7,
  input  [15:0] io_Stationary_matrix_3_0,
  input  [15:0] io_Stationary_matrix_3_1,
  input  [15:0] io_Stationary_matrix_3_2,
  input  [15:0] io_Stationary_matrix_3_3,
  input  [15:0] io_Stationary_matrix_3_4,
  input  [15:0] io_Stationary_matrix_3_5,
  input  [15:0] io_Stationary_matrix_3_6,
  input  [15:0] io_Stationary_matrix_3_7,
  input  [15:0] io_Stationary_matrix_4_0,
  input  [15:0] io_Stationary_matrix_4_1,
  input  [15:0] io_Stationary_matrix_4_2,
  input  [15:0] io_Stationary_matrix_4_3,
  input  [15:0] io_Stationary_matrix_4_4,
  input  [15:0] io_Stationary_matrix_4_5,
  input  [15:0] io_Stationary_matrix_4_6,
  input  [15:0] io_Stationary_matrix_4_7,
  input  [15:0] io_Stationary_matrix_5_0,
  input  [15:0] io_Stationary_matrix_5_1,
  input  [15:0] io_Stationary_matrix_5_2,
  input  [15:0] io_Stationary_matrix_5_3,
  input  [15:0] io_Stationary_matrix_5_4,
  input  [15:0] io_Stationary_matrix_5_5,
  input  [15:0] io_Stationary_matrix_5_6,
  input  [15:0] io_Stationary_matrix_5_7,
  input  [15:0] io_Stationary_matrix_6_0,
  input  [15:0] io_Stationary_matrix_6_1,
  input  [15:0] io_Stationary_matrix_6_2,
  input  [15:0] io_Stationary_matrix_6_3,
  input  [15:0] io_Stationary_matrix_6_4,
  input  [15:0] io_Stationary_matrix_6_5,
  input  [15:0] io_Stationary_matrix_6_6,
  input  [15:0] io_Stationary_matrix_6_7,
  input  [15:0] io_Stationary_matrix_7_0,
  input  [15:0] io_Stationary_matrix_7_1,
  input  [15:0] io_Stationary_matrix_7_2,
  input  [15:0] io_Stationary_matrix_7_3,
  input  [15:0] io_Stationary_matrix_7_4,
  input  [15:0] io_Stationary_matrix_7_5,
  input  [15:0] io_Stationary_matrix_7_6,
  input  [15:0] io_Stationary_matrix_7_7,
  output [4:0]  io_o_vn_0,
  output [4:0]  io_o_vn_1,
  output [4:0]  io_o_vn_2,
  output [4:0]  io_o_vn_3,
  output [4:0]  io_o_vn2_0,
  output [4:0]  io_o_vn2_1,
  output [4:0]  io_o_vn2_2,
  output [4:0]  io_o_vn2_3,
  output        io_ProcessValid,
  input         io_validpin
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
`endif // RANDOMIZE_REG_INIT
  reg [4:0] i_vn_0; // @[ivncontrol4.scala 17:23]
  reg [4:0] i_vn_1; // @[ivncontrol4.scala 17:23]
  reg [4:0] i_vn_2; // @[ivncontrol4.scala 17:23]
  reg [4:0] i_vn_3; // @[ivncontrol4.scala 17:23]
  reg [4:0] i_vn2_0; // @[ivncontrol4.scala 18:24]
  reg [4:0] i_vn2_1; // @[ivncontrol4.scala 18:24]
  reg [4:0] i_vn2_2; // @[ivncontrol4.scala 18:24]
  reg [4:0] i_vn2_3; // @[ivncontrol4.scala 18:24]
  reg [15:0] solution_0_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_0_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_0_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_0_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_0_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_0_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_0_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_0_7; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_7; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_7; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_7; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_7; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_7; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_7; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_7; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_0; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_1; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_2; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_3; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_4; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_5; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_6; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_7; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_8; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_9; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_10; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_11; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_12; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_13; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_14; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_15; // @[ivncontrol4.scala 27:27]
  reg [31:0] pin; // @[ivncontrol4.scala 37:22]
  reg [31:0] i; // @[ivncontrol4.scala 41:20]
  reg [31:0] j; // @[ivncontrol4.scala 42:20]
  wire  _io_ProcessValid_T = i == 32'h7; // @[ivncontrol4.scala 44:27]
  wire  _io_ProcessValid_T_1 = j == 32'h7; // @[ivncontrol4.scala 44:42]
  wire  _io_ProcessValid_T_2 = i == 32'h7 & j == 32'h7; // @[ivncontrol4.scala 44:36]
  reg [31:0] mat_0_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_0_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_0_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_0_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_0_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_0_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_0_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_0_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] count_0; // @[ivncontrol4.scala 58:20]
  reg [31:0] count_1; // @[ivncontrol4.scala 58:20]
  reg [31:0] count_2; // @[ivncontrol4.scala 58:20]
  reg [31:0] count_3; // @[ivncontrol4.scala 58:20]
  reg [31:0] count_4; // @[ivncontrol4.scala 58:20]
  reg [31:0] count_5; // @[ivncontrol4.scala 58:20]
  reg [31:0] count_6; // @[ivncontrol4.scala 58:20]
  reg [31:0] count_7; // @[ivncontrol4.scala 58:20]
  wire  _GEN_3825 = 3'h0 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_65 = 3'h0 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_0_1 : io_Stationary_matrix_0_0; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_66 = 3'h0 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_0_2 : _GEN_65; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_67 = 3'h0 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_0_3 : _GEN_66; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_68 = 3'h0 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_0_4 : _GEN_67; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_69 = 3'h0 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_0_5 : _GEN_68; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_70 = 3'h0 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_0_6 : _GEN_69; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_71 = 3'h0 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_0_7 : _GEN_70; // @[ivncontrol4.scala 63:{17,17}]
  wire  _GEN_3839 = 3'h1 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_72 = 3'h1 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_1_0 : _GEN_71; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_73 = 3'h1 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_1_1 : _GEN_72; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_74 = 3'h1 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_1_2 : _GEN_73; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_75 = 3'h1 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_1_3 : _GEN_74; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_76 = 3'h1 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_1_4 : _GEN_75; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_77 = 3'h1 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_1_5 : _GEN_76; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_78 = 3'h1 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_1_6 : _GEN_77; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_79 = 3'h1 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_1_7 : _GEN_78; // @[ivncontrol4.scala 63:{17,17}]
  wire  _GEN_3855 = 3'h2 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_80 = 3'h2 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_2_0 : _GEN_79; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_81 = 3'h2 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_2_1 : _GEN_80; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_82 = 3'h2 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_2_2 : _GEN_81; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_83 = 3'h2 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_2_3 : _GEN_82; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_84 = 3'h2 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_2_4 : _GEN_83; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_85 = 3'h2 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_2_5 : _GEN_84; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_86 = 3'h2 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_2_6 : _GEN_85; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_87 = 3'h2 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_2_7 : _GEN_86; // @[ivncontrol4.scala 63:{17,17}]
  wire  _GEN_3871 = 3'h3 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_88 = 3'h3 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_3_0 : _GEN_87; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_89 = 3'h3 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_3_1 : _GEN_88; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_90 = 3'h3 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_3_2 : _GEN_89; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_91 = 3'h3 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_3_3 : _GEN_90; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_92 = 3'h3 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_3_4 : _GEN_91; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_93 = 3'h3 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_3_5 : _GEN_92; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_94 = 3'h3 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_3_6 : _GEN_93; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_95 = 3'h3 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_3_7 : _GEN_94; // @[ivncontrol4.scala 63:{17,17}]
  wire  _GEN_3887 = 3'h4 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_96 = 3'h4 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_4_0 : _GEN_95; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_97 = 3'h4 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_4_1 : _GEN_96; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_98 = 3'h4 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_4_2 : _GEN_97; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_99 = 3'h4 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_4_3 : _GEN_98; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_100 = 3'h4 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_4_4 : _GEN_99; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_101 = 3'h4 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_4_5 : _GEN_100; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_102 = 3'h4 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_4_6 : _GEN_101; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_103 = 3'h4 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_4_7 : _GEN_102; // @[ivncontrol4.scala 63:{17,17}]
  wire  _GEN_3903 = 3'h5 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_104 = 3'h5 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_5_0 : _GEN_103; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_105 = 3'h5 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_5_1 : _GEN_104; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_106 = 3'h5 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_5_2 : _GEN_105; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_107 = 3'h5 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_5_3 : _GEN_106; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_108 = 3'h5 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_5_4 : _GEN_107; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_109 = 3'h5 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_5_5 : _GEN_108; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_110 = 3'h5 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_5_6 : _GEN_109; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_111 = 3'h5 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_5_7 : _GEN_110; // @[ivncontrol4.scala 63:{17,17}]
  wire  _GEN_3919 = 3'h6 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_112 = 3'h6 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_6_0 : _GEN_111; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_113 = 3'h6 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_6_1 : _GEN_112; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_114 = 3'h6 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_6_2 : _GEN_113; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_115 = 3'h6 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_6_3 : _GEN_114; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_116 = 3'h6 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_6_4 : _GEN_115; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_117 = 3'h6 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_6_5 : _GEN_116; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_118 = 3'h6 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_6_6 : _GEN_117; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_119 = 3'h6 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_6_7 : _GEN_118; // @[ivncontrol4.scala 63:{17,17}]
  wire  _GEN_3935 = 3'h7 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_120 = 3'h7 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_7_0 : _GEN_119; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_121 = 3'h7 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_7_1 : _GEN_120; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_122 = 3'h7 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_7_2 : _GEN_121; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_123 = 3'h7 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_7_3 : _GEN_122; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_124 = 3'h7 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_7_4 : _GEN_123; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_125 = 3'h7 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_7_5 : _GEN_124; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_126 = 3'h7 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_7_6 : _GEN_125; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_127 = 3'h7 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_7_7 : _GEN_126; // @[ivncontrol4.scala 63:{17,17}]
  wire [31:0] _mat_T_1_T_2 = {{16'd0}, _GEN_127}; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_129 = _GEN_3825 & 4'h1 == j[3:0] ? solution_0_1 : solution_0_0; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_130 = _GEN_3825 & 4'h2 == j[3:0] ? solution_0_2 : _GEN_129; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_131 = _GEN_3825 & 4'h3 == j[3:0] ? solution_0_3 : _GEN_130; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_132 = _GEN_3825 & 4'h4 == j[3:0] ? solution_0_4 : _GEN_131; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_133 = _GEN_3825 & 4'h5 == j[3:0] ? solution_0_5 : _GEN_132; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_134 = _GEN_3825 & 4'h6 == j[3:0] ? solution_0_6 : _GEN_133; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_135 = _GEN_3825 & 4'h7 == j[3:0] ? solution_0_7 : _GEN_134; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_136 = _GEN_3825 & 4'h8 == j[3:0] ? 16'h0 : _GEN_135; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_137 = _GEN_3839 & 4'h0 == j[3:0] ? solution_1_0 : _GEN_136; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_138 = _GEN_3839 & 4'h1 == j[3:0] ? solution_1_1 : _GEN_137; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_139 = _GEN_3839 & 4'h2 == j[3:0] ? solution_1_2 : _GEN_138; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_140 = _GEN_3839 & 4'h3 == j[3:0] ? solution_1_3 : _GEN_139; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_141 = _GEN_3839 & 4'h4 == j[3:0] ? solution_1_4 : _GEN_140; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_142 = _GEN_3839 & 4'h5 == j[3:0] ? solution_1_5 : _GEN_141; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_143 = _GEN_3839 & 4'h6 == j[3:0] ? solution_1_6 : _GEN_142; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_144 = _GEN_3839 & 4'h7 == j[3:0] ? solution_1_7 : _GEN_143; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_145 = _GEN_3839 & 4'h8 == j[3:0] ? 16'h0 : _GEN_144; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_146 = _GEN_3855 & 4'h0 == j[3:0] ? solution_2_0 : _GEN_145; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_147 = _GEN_3855 & 4'h1 == j[3:0] ? solution_2_1 : _GEN_146; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_148 = _GEN_3855 & 4'h2 == j[3:0] ? solution_2_2 : _GEN_147; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_149 = _GEN_3855 & 4'h3 == j[3:0] ? solution_2_3 : _GEN_148; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_150 = _GEN_3855 & 4'h4 == j[3:0] ? solution_2_4 : _GEN_149; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_151 = _GEN_3855 & 4'h5 == j[3:0] ? solution_2_5 : _GEN_150; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_152 = _GEN_3855 & 4'h6 == j[3:0] ? solution_2_6 : _GEN_151; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_153 = _GEN_3855 & 4'h7 == j[3:0] ? solution_2_7 : _GEN_152; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_154 = _GEN_3855 & 4'h8 == j[3:0] ? 16'h0 : _GEN_153; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_155 = _GEN_3871 & 4'h0 == j[3:0] ? solution_3_0 : _GEN_154; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_156 = _GEN_3871 & 4'h1 == j[3:0] ? solution_3_1 : _GEN_155; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_157 = _GEN_3871 & 4'h2 == j[3:0] ? solution_3_2 : _GEN_156; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_158 = _GEN_3871 & 4'h3 == j[3:0] ? solution_3_3 : _GEN_157; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_159 = _GEN_3871 & 4'h4 == j[3:0] ? solution_3_4 : _GEN_158; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_160 = _GEN_3871 & 4'h5 == j[3:0] ? solution_3_5 : _GEN_159; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_161 = _GEN_3871 & 4'h6 == j[3:0] ? solution_3_6 : _GEN_160; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_162 = _GEN_3871 & 4'h7 == j[3:0] ? solution_3_7 : _GEN_161; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_163 = _GEN_3871 & 4'h8 == j[3:0] ? 16'h0 : _GEN_162; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_164 = _GEN_3887 & 4'h0 == j[3:0] ? solution_4_0 : _GEN_163; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_165 = _GEN_3887 & 4'h1 == j[3:0] ? solution_4_1 : _GEN_164; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_166 = _GEN_3887 & 4'h2 == j[3:0] ? solution_4_2 : _GEN_165; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_167 = _GEN_3887 & 4'h3 == j[3:0] ? solution_4_3 : _GEN_166; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_168 = _GEN_3887 & 4'h4 == j[3:0] ? solution_4_4 : _GEN_167; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_169 = _GEN_3887 & 4'h5 == j[3:0] ? solution_4_5 : _GEN_168; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_170 = _GEN_3887 & 4'h6 == j[3:0] ? solution_4_6 : _GEN_169; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_171 = _GEN_3887 & 4'h7 == j[3:0] ? solution_4_7 : _GEN_170; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_172 = _GEN_3887 & 4'h8 == j[3:0] ? 16'h0 : _GEN_171; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_173 = _GEN_3903 & 4'h0 == j[3:0] ? solution_5_0 : _GEN_172; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_174 = _GEN_3903 & 4'h1 == j[3:0] ? solution_5_1 : _GEN_173; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_175 = _GEN_3903 & 4'h2 == j[3:0] ? solution_5_2 : _GEN_174; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_176 = _GEN_3903 & 4'h3 == j[3:0] ? solution_5_3 : _GEN_175; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_177 = _GEN_3903 & 4'h4 == j[3:0] ? solution_5_4 : _GEN_176; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_178 = _GEN_3903 & 4'h5 == j[3:0] ? solution_5_5 : _GEN_177; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_179 = _GEN_3903 & 4'h6 == j[3:0] ? solution_5_6 : _GEN_178; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_180 = _GEN_3903 & 4'h7 == j[3:0] ? solution_5_7 : _GEN_179; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_181 = _GEN_3903 & 4'h8 == j[3:0] ? 16'h0 : _GEN_180; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_182 = _GEN_3919 & 4'h0 == j[3:0] ? solution_6_0 : _GEN_181; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_183 = _GEN_3919 & 4'h1 == j[3:0] ? solution_6_1 : _GEN_182; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_184 = _GEN_3919 & 4'h2 == j[3:0] ? solution_6_2 : _GEN_183; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_185 = _GEN_3919 & 4'h3 == j[3:0] ? solution_6_3 : _GEN_184; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_186 = _GEN_3919 & 4'h4 == j[3:0] ? solution_6_4 : _GEN_185; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_187 = _GEN_3919 & 4'h5 == j[3:0] ? solution_6_5 : _GEN_186; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_188 = _GEN_3919 & 4'h6 == j[3:0] ? solution_6_6 : _GEN_187; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_189 = _GEN_3919 & 4'h7 == j[3:0] ? solution_6_7 : _GEN_188; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_190 = _GEN_3919 & 4'h8 == j[3:0] ? 16'h0 : _GEN_189; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_191 = _GEN_3935 & 4'h0 == j[3:0] ? solution_7_0 : _GEN_190; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_192 = _GEN_3935 & 4'h1 == j[3:0] ? solution_7_1 : _GEN_191; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_193 = _GEN_3935 & 4'h2 == j[3:0] ? solution_7_2 : _GEN_192; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_194 = _GEN_3935 & 4'h3 == j[3:0] ? solution_7_3 : _GEN_193; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_195 = _GEN_3935 & 4'h4 == j[3:0] ? solution_7_4 : _GEN_194; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_196 = _GEN_3935 & 4'h5 == j[3:0] ? solution_7_5 : _GEN_195; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_197 = _GEN_3935 & 4'h6 == j[3:0] ? solution_7_6 : _GEN_196; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_198 = _GEN_3935 & 4'h7 == j[3:0] ? solution_7_7 : _GEN_197; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_199 = _GEN_3935 & 4'h8 == j[3:0] ? 16'h0 : _GEN_198; // @[ivncontrol4.scala 65:{31,31}]
  wire [31:0] _GEN_201 = 3'h1 == i[2:0] ? count_1 : count_0; // @[ivncontrol4.scala 66:{33,33}]
  wire [31:0] _GEN_202 = 3'h2 == i[2:0] ? count_2 : _GEN_201; // @[ivncontrol4.scala 66:{33,33}]
  wire [31:0] _GEN_203 = 3'h3 == i[2:0] ? count_3 : _GEN_202; // @[ivncontrol4.scala 66:{33,33}]
  wire [31:0] _GEN_204 = 3'h4 == i[2:0] ? count_4 : _GEN_203; // @[ivncontrol4.scala 66:{33,33}]
  wire [31:0] _GEN_205 = 3'h5 == i[2:0] ? count_5 : _GEN_204; // @[ivncontrol4.scala 66:{33,33}]
  wire [31:0] _GEN_206 = 3'h6 == i[2:0] ? count_6 : _GEN_205; // @[ivncontrol4.scala 66:{33,33}]
  wire [31:0] _GEN_207 = 3'h7 == i[2:0] ? count_7 : _GEN_206; // @[ivncontrol4.scala 66:{33,33}]
  wire [31:0] _count_T_2 = _GEN_207 + 32'h1; // @[ivncontrol4.scala 66:33]
  wire [31:0] _GEN_208 = 3'h0 == i[2:0] ? _count_T_2 : count_0; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_209 = 3'h1 == i[2:0] ? _count_T_2 : count_1; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_210 = 3'h2 == i[2:0] ? _count_T_2 : count_2; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_211 = 3'h3 == i[2:0] ? _count_T_2 : count_3; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_212 = 3'h4 == i[2:0] ? _count_T_2 : count_4; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_213 = 3'h5 == i[2:0] ? _count_T_2 : count_5; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_214 = 3'h6 == i[2:0] ? _count_T_2 : count_6; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_215 = 3'h7 == i[2:0] ? _count_T_2 : count_7; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_216 = _GEN_199 != 16'h0 ? _GEN_208 : count_0; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_217 = _GEN_199 != 16'h0 ? _GEN_209 : count_1; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_218 = _GEN_199 != 16'h0 ? _GEN_210 : count_2; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_219 = _GEN_199 != 16'h0 ? _GEN_211 : count_3; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_220 = _GEN_199 != 16'h0 ? _GEN_212 : count_4; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_221 = _GEN_199 != 16'h0 ? _GEN_213 : count_5; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_222 = _GEN_199 != 16'h0 ? _GEN_214 : count_6; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_223 = _GEN_199 != 16'h0 ? _GEN_215 : count_7; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_224 = io_validpin ? _GEN_216 : count_0; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _GEN_225 = io_validpin ? _GEN_217 : count_1; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _GEN_226 = io_validpin ? _GEN_218 : count_2; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _GEN_227 = io_validpin ? _GEN_219 : count_3; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _GEN_228 = io_validpin ? _GEN_220 : count_4; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _GEN_229 = io_validpin ? _GEN_221 : count_5; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _GEN_230 = io_validpin ? _GEN_222 : count_6; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _GEN_231 = io_validpin ? _GEN_223 : count_7; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _i_T_1 = i + 32'h1; // @[ivncontrol4.scala 113:16]
  wire [31:0] _GEN_247 = i < 32'h7 & _io_ProcessValid_T_1 ? _i_T_1 : i; // @[ivncontrol4.scala 112:74 113:11 41:20]
  wire [31:0] _j_T_1 = j + 32'h1; // @[ivncontrol4.scala 118:16]
  wire [3:0] _GEN_264 = _io_ProcessValid_T & j == 32'h8 ? 4'h8 : 4'h0; // @[ivncontrol4.scala 120:77 121:11 129:11]
  wire [31:0] _GEN_265 = _io_ProcessValid_T & j == 32'h8 ? 32'h7 : _GEN_247; // @[ivncontrol4.scala 120:77 122:11]
  wire  _GEN_312 = _io_ProcessValid_T_2; // @[ivncontrol4.scala 153:41]
  wire [31:0] _GEN_313 = rowcount_0 != 32'h0 ? 32'h0 : pin; // @[ivncontrol4.scala 162:30 163:13 37:22]
  wire  _T_27 = rowcount_0 == 32'h0; // @[ivncontrol4.scala 165:23]
  wire [31:0] _GEN_314 = rowcount_0 == 32'h0 & rowcount_1 != 32'h0 ? 32'h1 : _GEN_313; // @[ivncontrol4.scala 165:54 166:13]
  wire  _T_32 = _T_27 & rowcount_1 == 32'h0; // @[ivncontrol4.scala 168:31]
  wire [31:0] _GEN_315 = _T_27 & rowcount_1 == 32'h0 & rowcount_2 != 32'h0 ? 32'h2 : _GEN_314; // @[ivncontrol4.scala 168:77 169:13]
  wire  _T_39 = _T_32 & rowcount_2 == 32'h0; // @[ivncontrol4.scala 171:54]
  wire [31:0] _GEN_316 = _T_32 & rowcount_2 == 32'h0 & rowcount_3 != 32'h0 ? 32'h3 : _GEN_315; // @[ivncontrol4.scala 171:100 172:13]
  wire  _T_48 = _T_39 & rowcount_3 == 32'h0; // @[ivncontrol4.scala 174:77]
  wire [31:0] _GEN_317 = _T_39 & rowcount_3 == 32'h0 & rowcount_4 != 32'h0 ? 32'h4 : _GEN_316; // @[ivncontrol4.scala 174:123 175:13]
  wire  _T_59 = _T_48 & rowcount_4 == 32'h0; // @[ivncontrol4.scala 177:100]
  wire  _T_72 = _T_59 & rowcount_5 == 32'h0; // @[ivncontrol4.scala 180:123]
  wire  valid = _io_ProcessValid_T_2; // @[ivncontrol4.scala 153:41]
  wire [32:0] _T_91 = {{1'd0}, pin}; // @[ivncontrol4.scala 191:27]
  wire [31:0] _GEN_322 = 4'h1 == _T_91[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_323 = 4'h2 == _T_91[3:0] ? rowcount_2 : _GEN_322; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_324 = 4'h3 == _T_91[3:0] ? rowcount_3 : _GEN_323; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_325 = 4'h4 == _T_91[3:0] ? rowcount_4 : _GEN_324; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_326 = 4'h5 == _T_91[3:0] ? rowcount_5 : _GEN_325; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_327 = 4'h6 == _T_91[3:0] ? rowcount_6 : _GEN_326; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_328 = 4'h7 == _T_91[3:0] ? rowcount_7 : _GEN_327; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_329 = 4'h8 == _T_91[3:0] ? rowcount_8 : _GEN_328; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_330 = 4'h9 == _T_91[3:0] ? rowcount_9 : _GEN_329; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_331 = 4'ha == _T_91[3:0] ? rowcount_10 : _GEN_330; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_332 = 4'hb == _T_91[3:0] ? rowcount_11 : _GEN_331; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_333 = 4'hc == _T_91[3:0] ? rowcount_12 : _GEN_332; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_334 = 4'hd == _T_91[3:0] ? rowcount_13 : _GEN_333; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_335 = 4'he == _T_91[3:0] ? rowcount_14 : _GEN_334; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_336 = 4'hf == _T_91[3:0] ? rowcount_15 : _GEN_335; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_449 = _GEN_336 == 32'h1 ? _T_91[31:0] : 32'ha; // @[ivncontrol4.scala 142:17 241:50 242:21]
  wire [31:0] _GEN_450 = _GEN_336 == 32'h2 ? _T_91[31:0] : _GEN_449; // @[ivncontrol4.scala 237:51 238:21]
  wire [31:0] _GEN_451 = _GEN_336 == 32'h2 ? _T_91[31:0] : 32'h1c; // @[ivncontrol4.scala 142:17 237:51 239:21]
  wire [31:0] _GEN_452 = _GEN_336 == 32'h3 ? _T_91[31:0] : _GEN_450; // @[ivncontrol4.scala 232:50 233:21]
  wire [31:0] _GEN_453 = _GEN_336 == 32'h3 ? _T_91[31:0] : _GEN_451; // @[ivncontrol4.scala 232:50 234:21]
  wire [31:0] _GEN_454 = _GEN_336 == 32'h3 ? _T_91[31:0] : 32'h14; // @[ivncontrol4.scala 142:17 232:50 235:21]
  wire [31:0] _GEN_455 = _GEN_336 == 32'h4 ? _T_91[31:0] : _GEN_452; // @[ivncontrol4.scala 224:50 225:21]
  wire [31:0] _GEN_456 = _GEN_336 == 32'h4 ? _T_91[31:0] : _GEN_453; // @[ivncontrol4.scala 224:50 226:21]
  wire [31:0] _GEN_457 = _GEN_336 == 32'h4 ? _T_91[31:0] : _GEN_454; // @[ivncontrol4.scala 224:50 227:21]
  wire [31:0] _GEN_458 = _GEN_336 == 32'h4 ? _T_91[31:0] : 32'h0; // @[ivncontrol4.scala 142:17 224:50 228:21]
  wire [31:0] _GEN_459 = _GEN_336 == 32'h5 ? _T_91[31:0] : _GEN_455; // @[ivncontrol4.scala 217:50 218:21]
  wire [31:0] _GEN_460 = _GEN_336 == 32'h5 ? _T_91[31:0] : _GEN_456; // @[ivncontrol4.scala 217:50 219:21]
  wire [31:0] _GEN_461 = _GEN_336 == 32'h5 ? _T_91[31:0] : _GEN_457; // @[ivncontrol4.scala 217:50 220:21]
  wire [31:0] _GEN_462 = _GEN_336 == 32'h5 ? _T_91[31:0] : _GEN_458; // @[ivncontrol4.scala 217:50 221:21]
  wire [31:0] _GEN_463 = _GEN_336 == 32'h5 ? _T_91[31:0] : 32'h1d; // @[ivncontrol4.scala 143:18 217:50 222:22]
  wire [31:0] _GEN_464 = _GEN_336 == 32'h6 ? _T_91[31:0] : _GEN_459; // @[ivncontrol4.scala 209:52 210:21]
  wire [31:0] _GEN_465 = _GEN_336 == 32'h6 ? _T_91[31:0] : _GEN_460; // @[ivncontrol4.scala 209:52 211:21]
  wire [31:0] _GEN_466 = _GEN_336 == 32'h6 ? _T_91[31:0] : _GEN_461; // @[ivncontrol4.scala 209:52 212:21]
  wire [31:0] _GEN_467 = _GEN_336 == 32'h6 ? _T_91[31:0] : _GEN_462; // @[ivncontrol4.scala 209:52 213:21]
  wire [31:0] _GEN_468 = _GEN_336 == 32'h6 ? _T_91[31:0] : _GEN_463; // @[ivncontrol4.scala 209:52 214:22]
  wire [31:0] _GEN_469 = _GEN_336 == 32'h6 ? _T_91[31:0] : 32'he; // @[ivncontrol4.scala 143:18 209:52 215:22]
  wire [31:0] _GEN_470 = _GEN_336 == 32'h7 ? _T_91[31:0] : _GEN_464; // @[ivncontrol4.scala 201:52 202:21]
  wire [31:0] _GEN_471 = _GEN_336 == 32'h7 ? _T_91[31:0] : _GEN_465; // @[ivncontrol4.scala 201:52 203:21]
  wire [31:0] _GEN_472 = _GEN_336 == 32'h7 ? _T_91[31:0] : _GEN_466; // @[ivncontrol4.scala 201:52 204:21]
  wire [31:0] _GEN_473 = _GEN_336 == 32'h7 ? _T_91[31:0] : _GEN_467; // @[ivncontrol4.scala 201:52 205:21]
  wire [31:0] _GEN_474 = _GEN_336 == 32'h7 ? _T_91[31:0] : _GEN_468; // @[ivncontrol4.scala 201:52 206:22]
  wire [31:0] _GEN_475 = _GEN_336 == 32'h7 ? _T_91[31:0] : _GEN_469; // @[ivncontrol4.scala 201:52 207:22]
  wire [31:0] _GEN_476 = _GEN_336 == 32'h7 ? _T_91[31:0] : 32'h8; // @[ivncontrol4.scala 143:18 201:52 208:22]
  wire [31:0] _GEN_477 = _GEN_336 >= 32'h8 ? _T_91[31:0] : _GEN_470; // @[ivncontrol4.scala 191:42 192:21]
  wire [31:0] _GEN_478 = _GEN_336 >= 32'h8 ? _T_91[31:0] : _GEN_471; // @[ivncontrol4.scala 191:42 193:21]
  wire [31:0] _GEN_479 = _GEN_336 >= 32'h8 ? _T_91[31:0] : _GEN_472; // @[ivncontrol4.scala 191:42 194:21]
  wire [31:0] _GEN_480 = _GEN_336 >= 32'h8 ? _T_91[31:0] : _GEN_473; // @[ivncontrol4.scala 191:42 195:21]
  wire [31:0] _GEN_481 = _GEN_336 >= 32'h8 ? _T_91[31:0] : _GEN_474; // @[ivncontrol4.scala 191:42 196:22]
  wire [31:0] _GEN_482 = _GEN_336 >= 32'h8 ? _T_91[31:0] : _GEN_475; // @[ivncontrol4.scala 191:42 197:22]
  wire [31:0] _GEN_483 = _GEN_336 >= 32'h8 ? _T_91[31:0] : _GEN_476; // @[ivncontrol4.scala 191:42 198:22]
  wire [31:0] _GEN_484 = _GEN_336 >= 32'h8 ? _T_91[31:0] : 32'h5; // @[ivncontrol4.scala 143:18 191:42 199:22]
  wire [31:0] _T_127 = 32'h8 - _GEN_336; // @[ivncontrol4.scala 245:18]
  wire [31:0] _i_vn_1_T_15 = 32'h1 + pin; // @[ivncontrol4.scala 246:29]
  wire [31:0] _GEN_597 = _T_127 == 32'h1 ? _i_vn_1_T_15 : _GEN_484; // @[ivncontrol4.scala 286:54 289:22]
  wire [31:0] _GEN_598 = _T_127 == 32'h2 ? _i_vn_1_T_15 : _GEN_483; // @[ivncontrol4.scala 281:54 284:22]
  wire [31:0] _GEN_599 = _T_127 == 32'h2 ? _i_vn_1_T_15 : _GEN_597; // @[ivncontrol4.scala 281:54 285:22]
  wire [31:0] _GEN_600 = _T_127 == 32'h3 ? _i_vn_1_T_15 : _GEN_482; // @[ivncontrol4.scala 274:54 276:22]
  wire [31:0] _GEN_601 = _T_127 == 32'h3 ? _i_vn_1_T_15 : _GEN_598; // @[ivncontrol4.scala 274:54 277:22]
  wire [31:0] _GEN_602 = _T_127 == 32'h3 ? _i_vn_1_T_15 : _GEN_599; // @[ivncontrol4.scala 274:54 278:22]
  wire [31:0] _GEN_603 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_481; // @[ivncontrol4.scala 268:54 270:22]
  wire [31:0] _GEN_604 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_600; // @[ivncontrol4.scala 268:54 271:22]
  wire [31:0] _GEN_605 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_601; // @[ivncontrol4.scala 268:54 272:22]
  wire [31:0] _GEN_606 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_602; // @[ivncontrol4.scala 268:54 273:22]
  wire [31:0] _GEN_607 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_480; // @[ivncontrol4.scala 261:54 263:21]
  wire [31:0] _GEN_608 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_603; // @[ivncontrol4.scala 261:54 264:22]
  wire [31:0] _GEN_609 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_604; // @[ivncontrol4.scala 261:54 265:22]
  wire [31:0] _GEN_610 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_605; // @[ivncontrol4.scala 261:54 266:22]
  wire [31:0] _GEN_611 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_606; // @[ivncontrol4.scala 261:54 267:22]
  wire [31:0] _GEN_612 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_479; // @[ivncontrol4.scala 254:54 255:22]
  wire [31:0] _GEN_613 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_607; // @[ivncontrol4.scala 254:54 256:21]
  wire [31:0] _GEN_614 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_608; // @[ivncontrol4.scala 254:54 257:22]
  wire [31:0] _GEN_615 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_609; // @[ivncontrol4.scala 254:54 258:22]
  wire [31:0] _GEN_616 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_610; // @[ivncontrol4.scala 254:54 259:22]
  wire [31:0] _GEN_617 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_611; // @[ivncontrol4.scala 254:54 260:22]
  wire [31:0] _GEN_618 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_478; // @[ivncontrol4.scala 245:49 246:22]
  wire [31:0] _GEN_619 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_612; // @[ivncontrol4.scala 245:49 247:21]
  wire [31:0] _GEN_620 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_613; // @[ivncontrol4.scala 245:49 248:21]
  wire [31:0] _GEN_621 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_614; // @[ivncontrol4.scala 245:49 249:22]
  wire [31:0] _GEN_622 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_615; // @[ivncontrol4.scala 245:49 250:22]
  wire [31:0] _GEN_623 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_616; // @[ivncontrol4.scala 245:49 251:22]
  wire [31:0] _GEN_624 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_617; // @[ivncontrol4.scala 245:49 252:22]
  wire [31:0] _GEN_642 = 4'h1 == _i_vn_1_T_15[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_643 = 4'h2 == _i_vn_1_T_15[3:0] ? rowcount_2 : _GEN_642; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_644 = 4'h3 == _i_vn_1_T_15[3:0] ? rowcount_3 : _GEN_643; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_645 = 4'h4 == _i_vn_1_T_15[3:0] ? rowcount_4 : _GEN_644; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_646 = 4'h5 == _i_vn_1_T_15[3:0] ? rowcount_5 : _GEN_645; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_647 = 4'h6 == _i_vn_1_T_15[3:0] ? rowcount_6 : _GEN_646; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_648 = 4'h7 == _i_vn_1_T_15[3:0] ? rowcount_7 : _GEN_647; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_649 = 4'h8 == _i_vn_1_T_15[3:0] ? rowcount_8 : _GEN_648; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_650 = 4'h9 == _i_vn_1_T_15[3:0] ? rowcount_9 : _GEN_649; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_651 = 4'ha == _i_vn_1_T_15[3:0] ? rowcount_10 : _GEN_650; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_652 = 4'hb == _i_vn_1_T_15[3:0] ? rowcount_11 : _GEN_651; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_653 = 4'hc == _i_vn_1_T_15[3:0] ? rowcount_12 : _GEN_652; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_654 = 4'hd == _i_vn_1_T_15[3:0] ? rowcount_13 : _GEN_653; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_655 = 4'he == _i_vn_1_T_15[3:0] ? rowcount_14 : _GEN_654; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_656 = 4'hf == _i_vn_1_T_15[3:0] ? rowcount_15 : _GEN_655; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _T_172 = _GEN_336 + _GEN_656; // @[ivncontrol4.scala 292:41]
  wire [31:0] _T_174 = 32'h8 - _T_172; // @[ivncontrol4.scala 292:18]
  wire [31:0] _i_vn_1_T_17 = 32'h2 + pin; // @[ivncontrol4.scala 293:29]
  wire [31:0] _GEN_849 = _T_174 == 32'h1 ? _i_vn_1_T_17 : _GEN_624; // @[ivncontrol4.scala 335:78 338:22]
  wire [31:0] _GEN_850 = _T_174 == 32'h2 ? _i_vn_1_T_17 : _GEN_623; // @[ivncontrol4.scala 329:76 332:22]
  wire [31:0] _GEN_851 = _T_174 == 32'h2 ? _i_vn_1_T_17 : _GEN_849; // @[ivncontrol4.scala 329:76 333:22]
  wire [31:0] _GEN_852 = _T_174 == 32'h3 ? _i_vn_1_T_17 : _GEN_622; // @[ivncontrol4.scala 322:78 324:23]
  wire [31:0] _GEN_853 = _T_174 == 32'h3 ? _i_vn_1_T_17 : _GEN_850; // @[ivncontrol4.scala 322:78 325:22]
  wire [31:0] _GEN_854 = _T_174 == 32'h3 ? _i_vn_1_T_17 : _GEN_851; // @[ivncontrol4.scala 322:78 326:22]
  wire [31:0] _GEN_855 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_621; // @[ivncontrol4.scala 316:78 318:22]
  wire [31:0] _GEN_856 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_852; // @[ivncontrol4.scala 316:78 319:22]
  wire [31:0] _GEN_857 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_853; // @[ivncontrol4.scala 316:78 320:22]
  wire [31:0] _GEN_858 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_854; // @[ivncontrol4.scala 316:78 321:22]
  wire [31:0] _GEN_859 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_620; // @[ivncontrol4.scala 309:76 311:23]
  wire [31:0] _GEN_860 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_855; // @[ivncontrol4.scala 309:76 312:22]
  wire [31:0] _GEN_861 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_856; // @[ivncontrol4.scala 309:76 313:22]
  wire [31:0] _GEN_862 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_857; // @[ivncontrol4.scala 309:76 314:22]
  wire [31:0] _GEN_863 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_858; // @[ivncontrol4.scala 309:76 315:22]
  wire [31:0] _GEN_864 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_619; // @[ivncontrol4.scala 301:77 303:22]
  wire [31:0] _GEN_865 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_859; // @[ivncontrol4.scala 301:77 304:21]
  wire [31:0] _GEN_866 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_860; // @[ivncontrol4.scala 301:77 305:22]
  wire [31:0] _GEN_867 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_861; // @[ivncontrol4.scala 301:77 306:22]
  wire [31:0] _GEN_868 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_862; // @[ivncontrol4.scala 301:77 307:22]
  wire [31:0] _GEN_869 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_863; // @[ivncontrol4.scala 301:77 308:22]
  wire [31:0] _GEN_870 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_618; // @[ivncontrol4.scala 292:73 293:22]
  wire [31:0] _GEN_871 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_864; // @[ivncontrol4.scala 292:73 294:21]
  wire [31:0] _GEN_872 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_865; // @[ivncontrol4.scala 292:73 295:21]
  wire [31:0] _GEN_873 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_866; // @[ivncontrol4.scala 292:73 296:22]
  wire [31:0] _GEN_874 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_867; // @[ivncontrol4.scala 292:73 297:22]
  wire [31:0] _GEN_875 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_868; // @[ivncontrol4.scala 292:73 298:22]
  wire [31:0] _GEN_876 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_869; // @[ivncontrol4.scala 292:73 299:22]
  wire [31:0] _GEN_910 = 4'h1 == _i_vn_1_T_17[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_911 = 4'h2 == _i_vn_1_T_17[3:0] ? rowcount_2 : _GEN_910; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_912 = 4'h3 == _i_vn_1_T_17[3:0] ? rowcount_3 : _GEN_911; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_913 = 4'h4 == _i_vn_1_T_17[3:0] ? rowcount_4 : _GEN_912; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_914 = 4'h5 == _i_vn_1_T_17[3:0] ? rowcount_5 : _GEN_913; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_915 = 4'h6 == _i_vn_1_T_17[3:0] ? rowcount_6 : _GEN_914; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_916 = 4'h7 == _i_vn_1_T_17[3:0] ? rowcount_7 : _GEN_915; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_917 = 4'h8 == _i_vn_1_T_17[3:0] ? rowcount_8 : _GEN_916; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_918 = 4'h9 == _i_vn_1_T_17[3:0] ? rowcount_9 : _GEN_917; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_919 = 4'ha == _i_vn_1_T_17[3:0] ? rowcount_10 : _GEN_918; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_920 = 4'hb == _i_vn_1_T_17[3:0] ? rowcount_11 : _GEN_919; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_921 = 4'hc == _i_vn_1_T_17[3:0] ? rowcount_12 : _GEN_920; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_922 = 4'hd == _i_vn_1_T_17[3:0] ? rowcount_13 : _GEN_921; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_923 = 4'he == _i_vn_1_T_17[3:0] ? rowcount_14 : _GEN_922; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_924 = 4'hf == _i_vn_1_T_17[3:0] ? rowcount_15 : _GEN_923; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _T_254 = _T_172 + _GEN_924; // @[ivncontrol4.scala 343:62]
  wire [31:0] _T_256 = 32'h8 - _T_254; // @[ivncontrol4.scala 343:17]
  wire [31:0] _i_vn_1_T_19 = 32'h3 + pin; // @[ivncontrol4.scala 344:29]
  wire [31:0] _GEN_1213 = _T_256 == 32'h1 ? _i_vn_1_T_19 : _GEN_876; // @[ivncontrol4.scala 386:100 389:22]
  wire [31:0] _GEN_1214 = _T_256 == 32'h2 ? _i_vn_1_T_19 : _GEN_875; // @[ivncontrol4.scala 380:98 383:22]
  wire [31:0] _GEN_1215 = _T_256 == 32'h2 ? _i_vn_1_T_19 : _GEN_1213; // @[ivncontrol4.scala 380:98 384:22]
  wire [31:0] _GEN_1216 = _T_256 == 32'h3 ? _i_vn_1_T_19 : _GEN_874; // @[ivncontrol4.scala 373:100 375:23]
  wire [31:0] _GEN_1217 = _T_256 == 32'h3 ? _i_vn_1_T_19 : _GEN_1214; // @[ivncontrol4.scala 373:100 376:22]
  wire [31:0] _GEN_1218 = _T_256 == 32'h3 ? _i_vn_1_T_19 : _GEN_1215; // @[ivncontrol4.scala 373:100 377:22]
  wire [31:0] _GEN_1219 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_873; // @[ivncontrol4.scala 367:100 369:22]
  wire [31:0] _GEN_1220 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_1216; // @[ivncontrol4.scala 367:100 370:22]
  wire [31:0] _GEN_1221 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_1217; // @[ivncontrol4.scala 367:100 371:22]
  wire [31:0] _GEN_1222 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_1218; // @[ivncontrol4.scala 367:100 372:22]
  wire [31:0] _GEN_1223 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_872; // @[ivncontrol4.scala 360:98 362:23]
  wire [31:0] _GEN_1224 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1219; // @[ivncontrol4.scala 360:98 363:22]
  wire [31:0] _GEN_1225 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1220; // @[ivncontrol4.scala 360:98 364:22]
  wire [31:0] _GEN_1226 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1221; // @[ivncontrol4.scala 360:98 365:22]
  wire [31:0] _GEN_1227 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1222; // @[ivncontrol4.scala 360:98 366:22]
  wire [31:0] _GEN_1228 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_871; // @[ivncontrol4.scala 352:99 354:22]
  wire [31:0] _GEN_1229 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1223; // @[ivncontrol4.scala 352:99 355:21]
  wire [31:0] _GEN_1230 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1224; // @[ivncontrol4.scala 352:99 356:22]
  wire [31:0] _GEN_1231 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1225; // @[ivncontrol4.scala 352:99 357:22]
  wire [31:0] _GEN_1232 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1226; // @[ivncontrol4.scala 352:99 358:22]
  wire [31:0] _GEN_1233 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1227; // @[ivncontrol4.scala 352:99 359:22]
  wire [31:0] _GEN_1234 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_870; // @[ivncontrol4.scala 343:94 344:22]
  wire [31:0] _GEN_1235 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1228; // @[ivncontrol4.scala 343:94 345:21]
  wire [31:0] _GEN_1236 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1229; // @[ivncontrol4.scala 343:94 346:21]
  wire [31:0] _GEN_1237 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1230; // @[ivncontrol4.scala 343:94 347:22]
  wire [31:0] _GEN_1238 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1231; // @[ivncontrol4.scala 343:94 348:22]
  wire [31:0] _GEN_1239 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1232; // @[ivncontrol4.scala 343:94 349:22]
  wire [31:0] _GEN_1240 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1233; // @[ivncontrol4.scala 343:94 350:22]
  wire [31:0] _GEN_1290 = 4'h1 == _i_vn_1_T_19[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1291 = 4'h2 == _i_vn_1_T_19[3:0] ? rowcount_2 : _GEN_1290; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1292 = 4'h3 == _i_vn_1_T_19[3:0] ? rowcount_3 : _GEN_1291; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1293 = 4'h4 == _i_vn_1_T_19[3:0] ? rowcount_4 : _GEN_1292; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1294 = 4'h5 == _i_vn_1_T_19[3:0] ? rowcount_5 : _GEN_1293; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1295 = 4'h6 == _i_vn_1_T_19[3:0] ? rowcount_6 : _GEN_1294; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1296 = 4'h7 == _i_vn_1_T_19[3:0] ? rowcount_7 : _GEN_1295; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1297 = 4'h8 == _i_vn_1_T_19[3:0] ? rowcount_8 : _GEN_1296; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1298 = 4'h9 == _i_vn_1_T_19[3:0] ? rowcount_9 : _GEN_1297; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1299 = 4'ha == _i_vn_1_T_19[3:0] ? rowcount_10 : _GEN_1298; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1300 = 4'hb == _i_vn_1_T_19[3:0] ? rowcount_11 : _GEN_1299; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1301 = 4'hc == _i_vn_1_T_19[3:0] ? rowcount_12 : _GEN_1300; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1302 = 4'hd == _i_vn_1_T_19[3:0] ? rowcount_13 : _GEN_1301; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1303 = 4'he == _i_vn_1_T_19[3:0] ? rowcount_14 : _GEN_1302; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1304 = 4'hf == _i_vn_1_T_19[3:0] ? rowcount_15 : _GEN_1303; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _T_371 = _T_254 + _GEN_1304; // @[ivncontrol4.scala 393:86]
  wire [31:0] _T_373 = 32'h8 - _T_371; // @[ivncontrol4.scala 393:19]
  wire [31:0] _i_vn_1_T_21 = 32'h4 + pin; // @[ivncontrol4.scala 394:29]
  wire [31:0] _GEN_1689 = _T_373 == 32'h1 ? _i_vn_1_T_21 : _GEN_1240; // @[ivncontrol4.scala 436:122 439:22]
  wire [31:0] _GEN_1690 = _T_373 == 32'h2 ? _i_vn_1_T_21 : _GEN_1239; // @[ivncontrol4.scala 430:121 433:22]
  wire [31:0] _GEN_1691 = _T_373 == 32'h2 ? _i_vn_1_T_21 : _GEN_1689; // @[ivncontrol4.scala 430:121 434:22]
  wire [31:0] _GEN_1692 = _T_373 == 32'h3 ? _i_vn_1_T_21 : _GEN_1238; // @[ivncontrol4.scala 423:123 425:23]
  wire [31:0] _GEN_1693 = _T_373 == 32'h3 ? _i_vn_1_T_21 : _GEN_1690; // @[ivncontrol4.scala 423:123 426:22]
  wire [31:0] _GEN_1694 = _T_373 == 32'h3 ? _i_vn_1_T_21 : _GEN_1691; // @[ivncontrol4.scala 423:123 427:22]
  wire [31:0] _GEN_1695 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1237; // @[ivncontrol4.scala 417:122 419:22]
  wire [31:0] _GEN_1696 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1692; // @[ivncontrol4.scala 417:122 420:22]
  wire [31:0] _GEN_1697 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1693; // @[ivncontrol4.scala 417:122 421:22]
  wire [31:0] _GEN_1698 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1694; // @[ivncontrol4.scala 417:122 422:22]
  wire [31:0] _GEN_1699 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1236; // @[ivncontrol4.scala 410:121 412:23]
  wire [31:0] _GEN_1700 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1695; // @[ivncontrol4.scala 410:121 413:22]
  wire [31:0] _GEN_1701 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1696; // @[ivncontrol4.scala 410:121 414:22]
  wire [31:0] _GEN_1702 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1697; // @[ivncontrol4.scala 410:121 415:22]
  wire [31:0] _GEN_1703 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1698; // @[ivncontrol4.scala 410:121 416:22]
  wire [31:0] _GEN_1704 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1235; // @[ivncontrol4.scala 402:121 404:22]
  wire [31:0] _GEN_1705 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1699; // @[ivncontrol4.scala 402:121 405:21]
  wire [31:0] _GEN_1706 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1700; // @[ivncontrol4.scala 402:121 406:22]
  wire [31:0] _GEN_1707 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1701; // @[ivncontrol4.scala 402:121 407:22]
  wire [31:0] _GEN_1708 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1702; // @[ivncontrol4.scala 402:121 408:22]
  wire [31:0] _GEN_1709 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1703; // @[ivncontrol4.scala 402:121 409:22]
  wire [31:0] _GEN_1710 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1234; // @[ivncontrol4.scala 393:118 394:22]
  wire [31:0] _GEN_1711 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1704; // @[ivncontrol4.scala 393:118 395:21]
  wire [31:0] _GEN_1712 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1705; // @[ivncontrol4.scala 393:118 396:21]
  wire [31:0] _GEN_1713 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1706; // @[ivncontrol4.scala 393:118 397:22]
  wire [31:0] _GEN_1714 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1707; // @[ivncontrol4.scala 393:118 398:22]
  wire [31:0] _GEN_1715 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1708; // @[ivncontrol4.scala 393:118 399:22]
  wire [31:0] _GEN_1716 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1709; // @[ivncontrol4.scala 393:118 400:22]
  wire [31:0] _GEN_1782 = 4'h1 == _i_vn_1_T_21[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1783 = 4'h2 == _i_vn_1_T_21[3:0] ? rowcount_2 : _GEN_1782; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1784 = 4'h3 == _i_vn_1_T_21[3:0] ? rowcount_3 : _GEN_1783; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1785 = 4'h4 == _i_vn_1_T_21[3:0] ? rowcount_4 : _GEN_1784; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1786 = 4'h5 == _i_vn_1_T_21[3:0] ? rowcount_5 : _GEN_1785; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1787 = 4'h6 == _i_vn_1_T_21[3:0] ? rowcount_6 : _GEN_1786; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1788 = 4'h7 == _i_vn_1_T_21[3:0] ? rowcount_7 : _GEN_1787; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1789 = 4'h8 == _i_vn_1_T_21[3:0] ? rowcount_8 : _GEN_1788; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1790 = 4'h9 == _i_vn_1_T_21[3:0] ? rowcount_9 : _GEN_1789; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1791 = 4'ha == _i_vn_1_T_21[3:0] ? rowcount_10 : _GEN_1790; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1792 = 4'hb == _i_vn_1_T_21[3:0] ? rowcount_11 : _GEN_1791; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1793 = 4'hc == _i_vn_1_T_21[3:0] ? rowcount_12 : _GEN_1792; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1794 = 4'hd == _i_vn_1_T_21[3:0] ? rowcount_13 : _GEN_1793; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1795 = 4'he == _i_vn_1_T_21[3:0] ? rowcount_14 : _GEN_1794; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1796 = 4'hf == _i_vn_1_T_21[3:0] ? rowcount_15 : _GEN_1795; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _T_523 = _T_371 + _GEN_1796; // @[ivncontrol4.scala 443:108]
  wire [31:0] _T_525 = 32'h8 - _T_523; // @[ivncontrol4.scala 443:19]
  wire [31:0] _i_vn_1_T_23 = 32'h5 + pin; // @[ivncontrol4.scala 444:29]
  wire [31:0] _GEN_2277 = _T_525 == 32'h1 ? _i_vn_1_T_23 : _GEN_1716; // @[ivncontrol4.scala 486:144 489:22]
  wire [31:0] _GEN_2278 = _T_525 == 32'h2 ? _i_vn_1_T_23 : _GEN_1715; // @[ivncontrol4.scala 480:143 483:22]
  wire [31:0] _GEN_2279 = _T_525 == 32'h2 ? _i_vn_1_T_23 : _GEN_2277; // @[ivncontrol4.scala 480:143 484:22]
  wire [31:0] _GEN_2280 = _T_525 == 32'h3 ? _i_vn_1_T_23 : _GEN_1714; // @[ivncontrol4.scala 473:145 475:23]
  wire [31:0] _GEN_2281 = _T_525 == 32'h3 ? _i_vn_1_T_23 : _GEN_2278; // @[ivncontrol4.scala 473:145 476:22]
  wire [31:0] _GEN_2282 = _T_525 == 32'h3 ? _i_vn_1_T_23 : _GEN_2279; // @[ivncontrol4.scala 473:145 477:22]
  wire [31:0] _GEN_2283 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_1713; // @[ivncontrol4.scala 467:143 469:22]
  wire [31:0] _GEN_2284 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_2280; // @[ivncontrol4.scala 467:143 470:22]
  wire [31:0] _GEN_2285 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_2281; // @[ivncontrol4.scala 467:143 471:22]
  wire [31:0] _GEN_2286 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_2282; // @[ivncontrol4.scala 467:143 472:22]
  wire [31:0] _GEN_2287 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_1712; // @[ivncontrol4.scala 460:143 462:23]
  wire [31:0] _GEN_2288 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2283; // @[ivncontrol4.scala 460:143 463:22]
  wire [31:0] _GEN_2289 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2284; // @[ivncontrol4.scala 460:143 464:22]
  wire [31:0] _GEN_2290 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2285; // @[ivncontrol4.scala 460:143 465:22]
  wire [31:0] _GEN_2291 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2286; // @[ivncontrol4.scala 460:143 466:22]
  wire [31:0] _GEN_2292 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_1711; // @[ivncontrol4.scala 452:143 454:22]
  wire [31:0] _GEN_2293 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2287; // @[ivncontrol4.scala 452:143 455:21]
  wire [31:0] _GEN_2294 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2288; // @[ivncontrol4.scala 452:143 456:22]
  wire [31:0] _GEN_2295 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2289; // @[ivncontrol4.scala 452:143 457:22]
  wire [31:0] _GEN_2296 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2290; // @[ivncontrol4.scala 452:143 458:22]
  wire [31:0] _GEN_2297 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2291; // @[ivncontrol4.scala 452:143 459:22]
  wire [31:0] _GEN_2298 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_1710; // @[ivncontrol4.scala 443:140 444:22]
  wire [31:0] _GEN_2299 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2292; // @[ivncontrol4.scala 443:140 445:21]
  wire [31:0] _GEN_2300 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2293; // @[ivncontrol4.scala 443:140 446:21]
  wire [31:0] _GEN_2301 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2294; // @[ivncontrol4.scala 443:140 447:22]
  wire [31:0] _GEN_2302 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2295; // @[ivncontrol4.scala 443:140 448:22]
  wire [31:0] _GEN_2303 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2296; // @[ivncontrol4.scala 443:140 449:22]
  wire [31:0] _GEN_2304 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2297; // @[ivncontrol4.scala 443:140 450:22]
  wire [31:0] _GEN_2386 = 4'h1 == _i_vn_1_T_23[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2387 = 4'h2 == _i_vn_1_T_23[3:0] ? rowcount_2 : _GEN_2386; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2388 = 4'h3 == _i_vn_1_T_23[3:0] ? rowcount_3 : _GEN_2387; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2389 = 4'h4 == _i_vn_1_T_23[3:0] ? rowcount_4 : _GEN_2388; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2390 = 4'h5 == _i_vn_1_T_23[3:0] ? rowcount_5 : _GEN_2389; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2391 = 4'h6 == _i_vn_1_T_23[3:0] ? rowcount_6 : _GEN_2390; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2392 = 4'h7 == _i_vn_1_T_23[3:0] ? rowcount_7 : _GEN_2391; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2393 = 4'h8 == _i_vn_1_T_23[3:0] ? rowcount_8 : _GEN_2392; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2394 = 4'h9 == _i_vn_1_T_23[3:0] ? rowcount_9 : _GEN_2393; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2395 = 4'ha == _i_vn_1_T_23[3:0] ? rowcount_10 : _GEN_2394; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2396 = 4'hb == _i_vn_1_T_23[3:0] ? rowcount_11 : _GEN_2395; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2397 = 4'hc == _i_vn_1_T_23[3:0] ? rowcount_12 : _GEN_2396; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2398 = 4'hd == _i_vn_1_T_23[3:0] ? rowcount_13 : _GEN_2397; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2399 = 4'he == _i_vn_1_T_23[3:0] ? rowcount_14 : _GEN_2398; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2400 = 4'hf == _i_vn_1_T_23[3:0] ? rowcount_15 : _GEN_2399; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _T_710 = _T_523 + _GEN_2400; // @[ivncontrol4.scala 494:130]
  wire [31:0] _T_712 = 32'h8 - _T_710; // @[ivncontrol4.scala 494:19]
  wire [31:0] _i_vn_1_T_25 = 32'h6 + pin; // @[ivncontrol4.scala 495:29]
  wire [31:0] _GEN_2977 = _T_712 == 32'h1 ? _i_vn_1_T_25 : _GEN_2304; // @[ivncontrol4.scala 537:166 540:22]
  wire [31:0] _GEN_2978 = _T_712 == 32'h2 ? _i_vn_1_T_25 : _GEN_2303; // @[ivncontrol4.scala 531:166 534:22]
  wire [31:0] _GEN_2979 = _T_712 == 32'h2 ? _i_vn_1_T_25 : _GEN_2977; // @[ivncontrol4.scala 531:166 535:22]
  wire [31:0] _GEN_2980 = _T_712 == 32'h3 ? _i_vn_1_T_25 : _GEN_2302; // @[ivncontrol4.scala 524:168 526:23]
  wire [31:0] _GEN_2981 = _T_712 == 32'h3 ? _i_vn_1_T_25 : _GEN_2978; // @[ivncontrol4.scala 524:168 527:22]
  wire [31:0] _GEN_2982 = _T_712 == 32'h3 ? _i_vn_1_T_25 : _GEN_2979; // @[ivncontrol4.scala 524:168 528:22]
  wire [31:0] _GEN_2983 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2301; // @[ivncontrol4.scala 518:166 520:22]
  wire [31:0] _GEN_2984 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2980; // @[ivncontrol4.scala 518:166 521:22]
  wire [31:0] _GEN_2985 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2981; // @[ivncontrol4.scala 518:166 522:22]
  wire [31:0] _GEN_2986 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2982; // @[ivncontrol4.scala 518:166 523:22]
  wire [31:0] _GEN_2987 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2300; // @[ivncontrol4.scala 511:166 513:23]
  wire [31:0] _GEN_2988 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2983; // @[ivncontrol4.scala 511:166 514:22]
  wire [31:0] _GEN_2989 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2984; // @[ivncontrol4.scala 511:166 515:22]
  wire [31:0] _GEN_2990 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2985; // @[ivncontrol4.scala 511:166 516:22]
  wire [31:0] _GEN_2991 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2986; // @[ivncontrol4.scala 511:166 517:22]
  wire [31:0] _GEN_2992 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2299; // @[ivncontrol4.scala 503:166 505:22]
  wire [31:0] _GEN_2993 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2987; // @[ivncontrol4.scala 503:166 506:21]
  wire [31:0] _GEN_2994 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2988; // @[ivncontrol4.scala 503:166 507:22]
  wire [31:0] _GEN_2995 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2989; // @[ivncontrol4.scala 503:166 508:22]
  wire [31:0] _GEN_2996 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2990; // @[ivncontrol4.scala 503:166 509:22]
  wire [31:0] _GEN_2997 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2991; // @[ivncontrol4.scala 503:166 510:22]
  wire [31:0] _GEN_2998 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2298; // @[ivncontrol4.scala 494:162 495:22]
  wire [31:0] _GEN_2999 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2992; // @[ivncontrol4.scala 494:162 496:21]
  wire [31:0] _GEN_3000 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2993; // @[ivncontrol4.scala 494:162 497:21]
  wire [31:0] _GEN_3001 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2994; // @[ivncontrol4.scala 494:162 498:22]
  wire [31:0] _GEN_3002 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2995; // @[ivncontrol4.scala 494:162 499:22]
  wire [31:0] _GEN_3003 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2996; // @[ivncontrol4.scala 494:162 500:22]
  wire [31:0] _GEN_3004 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2997; // @[ivncontrol4.scala 494:162 501:22]
  wire [31:0] _GEN_3102 = 4'h1 == _i_vn_1_T_25[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3103 = 4'h2 == _i_vn_1_T_25[3:0] ? rowcount_2 : _GEN_3102; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3104 = 4'h3 == _i_vn_1_T_25[3:0] ? rowcount_3 : _GEN_3103; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3105 = 4'h4 == _i_vn_1_T_25[3:0] ? rowcount_4 : _GEN_3104; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3106 = 4'h5 == _i_vn_1_T_25[3:0] ? rowcount_5 : _GEN_3105; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3107 = 4'h6 == _i_vn_1_T_25[3:0] ? rowcount_6 : _GEN_3106; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3108 = 4'h7 == _i_vn_1_T_25[3:0] ? rowcount_7 : _GEN_3107; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3109 = 4'h8 == _i_vn_1_T_25[3:0] ? rowcount_8 : _GEN_3108; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3110 = 4'h9 == _i_vn_1_T_25[3:0] ? rowcount_9 : _GEN_3109; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3111 = 4'ha == _i_vn_1_T_25[3:0] ? rowcount_10 : _GEN_3110; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3112 = 4'hb == _i_vn_1_T_25[3:0] ? rowcount_11 : _GEN_3111; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3113 = 4'hc == _i_vn_1_T_25[3:0] ? rowcount_12 : _GEN_3112; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3114 = 4'hd == _i_vn_1_T_25[3:0] ? rowcount_13 : _GEN_3113; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3115 = 4'he == _i_vn_1_T_25[3:0] ? rowcount_14 : _GEN_3114; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3116 = 4'hf == _i_vn_1_T_25[3:0] ? rowcount_15 : _GEN_3115; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _T_932 = _T_710 + _GEN_3116; // @[ivncontrol4.scala 545:152]
  wire [31:0] _T_934 = 32'h8 - _T_932; // @[ivncontrol4.scala 545:19]
  wire [31:0] _i_vn_1_T_27 = 32'h7 + pin; // @[ivncontrol4.scala 546:29]
  wire [31:0] _GEN_3789 = _T_934 == 32'h1 ? _i_vn_1_T_27 : _GEN_3004; // @[ivncontrol4.scala 588:188 591:22]
  wire [31:0] _GEN_3790 = _T_934 == 32'h2 ? _i_vn_1_T_27 : _GEN_3003; // @[ivncontrol4.scala 582:188 585:22]
  wire [31:0] _GEN_3791 = _T_934 == 32'h2 ? _i_vn_1_T_27 : _GEN_3789; // @[ivncontrol4.scala 582:188 586:22]
  wire [31:0] _GEN_3792 = _T_934 == 32'h3 ? _i_vn_1_T_27 : _GEN_3002; // @[ivncontrol4.scala 575:190 577:23]
  wire [31:0] _GEN_3793 = _T_934 == 32'h3 ? _i_vn_1_T_27 : _GEN_3790; // @[ivncontrol4.scala 575:190 578:22]
  wire [31:0] _GEN_3794 = _T_934 == 32'h3 ? _i_vn_1_T_27 : _GEN_3791; // @[ivncontrol4.scala 575:190 579:22]
  wire [31:0] _GEN_3795 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_3001; // @[ivncontrol4.scala 569:188 571:22]
  wire [31:0] _GEN_3796 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_3792; // @[ivncontrol4.scala 569:188 572:22]
  wire [31:0] _GEN_3797 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_3793; // @[ivncontrol4.scala 569:188 573:22]
  wire [31:0] _GEN_3798 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_3794; // @[ivncontrol4.scala 569:188 574:22]
  wire [31:0] _GEN_3799 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3000; // @[ivncontrol4.scala 562:188 564:23]
  wire [31:0] _GEN_3800 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3795; // @[ivncontrol4.scala 562:188 565:22]
  wire [31:0] _GEN_3801 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3796; // @[ivncontrol4.scala 562:188 566:22]
  wire [31:0] _GEN_3802 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3797; // @[ivncontrol4.scala 562:188 567:22]
  wire [31:0] _GEN_3803 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3798; // @[ivncontrol4.scala 562:188 568:22]
  wire [31:0] _GEN_3804 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_2999; // @[ivncontrol4.scala 554:188 556:22]
  wire [31:0] _GEN_3805 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3799; // @[ivncontrol4.scala 554:188 557:21]
  wire [31:0] _GEN_3806 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3800; // @[ivncontrol4.scala 554:188 558:22]
  wire [31:0] _GEN_3807 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3801; // @[ivncontrol4.scala 554:188 559:22]
  wire [31:0] _GEN_3808 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3802; // @[ivncontrol4.scala 554:188 560:22]
  wire [31:0] _GEN_3809 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3803; // @[ivncontrol4.scala 554:188 561:22]
  wire [31:0] _GEN_3810 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_2998; // @[ivncontrol4.scala 545:184 546:22]
  wire [31:0] _GEN_3811 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3804; // @[ivncontrol4.scala 545:184 547:21]
  wire [31:0] _GEN_3812 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3805; // @[ivncontrol4.scala 545:184 548:21]
  wire [31:0] _GEN_3813 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3806; // @[ivncontrol4.scala 545:184 549:22]
  wire [31:0] _GEN_3814 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3807; // @[ivncontrol4.scala 545:184 550:22]
  wire [31:0] _GEN_3815 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3808; // @[ivncontrol4.scala 545:184 551:22]
  wire [31:0] _GEN_3816 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3809; // @[ivncontrol4.scala 545:184 552:22]
  wire [31:0] _GEN_3817 = _GEN_312 ? _GEN_477 : 32'ha; // @[ivncontrol4.scala 142:17 189:28]
  wire [31:0] _GEN_3818 = _GEN_312 ? _GEN_3810 : 32'h1c; // @[ivncontrol4.scala 142:17 189:28]
  wire [31:0] _GEN_3819 = _GEN_312 ? _GEN_3811 : 32'h14; // @[ivncontrol4.scala 142:17 189:28]
  wire [31:0] _GEN_3820 = _GEN_312 ? _GEN_3812 : 32'h0; // @[ivncontrol4.scala 142:17 189:28]
  wire [31:0] _GEN_3821 = _GEN_312 ? _GEN_3813 : 32'h1d; // @[ivncontrol4.scala 143:18 189:28]
  wire [31:0] _GEN_3822 = _GEN_312 ? _GEN_3814 : 32'he; // @[ivncontrol4.scala 143:18 189:28]
  wire [31:0] _GEN_3823 = _GEN_312 ? _GEN_3815 : 32'h8; // @[ivncontrol4.scala 143:18 189:28]
  wire [31:0] _GEN_3824 = _GEN_312 ? _GEN_3816 : 32'h5; // @[ivncontrol4.scala 143:18 189:28]
  wire  valid1 = 1'h0;
  wire [31:0] _GEN_4221 = reset ? 32'h0 : _GEN_3817; // @[ivncontrol4.scala 17:{23,23}]
  wire [31:0] _GEN_4222 = reset ? 32'h0 : _GEN_3818; // @[ivncontrol4.scala 17:{23,23}]
  wire [31:0] _GEN_4223 = reset ? 32'h0 : _GEN_3819; // @[ivncontrol4.scala 17:{23,23}]
  wire [31:0] _GEN_4224 = reset ? 32'h0 : _GEN_3820; // @[ivncontrol4.scala 17:{23,23}]
  wire [31:0] _GEN_4225 = reset ? 32'h0 : _GEN_3821; // @[ivncontrol4.scala 18:{24,24}]
  wire [31:0] _GEN_4226 = reset ? 32'h0 : _GEN_3822; // @[ivncontrol4.scala 18:{24,24}]
  wire [31:0] _GEN_4227 = reset ? 32'h0 : _GEN_3823; // @[ivncontrol4.scala 18:{24,24}]
  wire [31:0] _GEN_4228 = reset ? 32'h0 : _GEN_3824; // @[ivncontrol4.scala 18:{24,24}]
  assign io_o_vn_0 = i_vn_0; // @[ivncontrol4.scala 138:13]
  assign io_o_vn_1 = i_vn_1; // @[ivncontrol4.scala 138:13]
  assign io_o_vn_2 = i_vn_2; // @[ivncontrol4.scala 138:13]
  assign io_o_vn_3 = i_vn_3; // @[ivncontrol4.scala 138:13]
  assign io_o_vn2_0 = i_vn2_0; // @[ivncontrol4.scala 139:14]
  assign io_o_vn2_1 = i_vn2_1; // @[ivncontrol4.scala 139:14]
  assign io_o_vn2_2 = i_vn2_2; // @[ivncontrol4.scala 139:14]
  assign io_o_vn2_3 = i_vn2_3; // @[ivncontrol4.scala 139:14]
  assign io_ProcessValid = io_validpin & (i == 32'h7 & j == 32'h7); // @[ivncontrol4.scala 135:21 44:21 46:29]
  always @(posedge clock) begin
    i_vn_0 <= _GEN_4221[4:0]; // @[ivncontrol4.scala 17:{23,23}]
    i_vn_1 <= _GEN_4222[4:0]; // @[ivncontrol4.scala 17:{23,23}]
    i_vn_2 <= _GEN_4223[4:0]; // @[ivncontrol4.scala 17:{23,23}]
    i_vn_3 <= _GEN_4224[4:0]; // @[ivncontrol4.scala 17:{23,23}]
    i_vn2_0 <= _GEN_4225[4:0]; // @[ivncontrol4.scala 18:{24,24}]
    i_vn2_1 <= _GEN_4226[4:0]; // @[ivncontrol4.scala 18:{24,24}]
    i_vn2_2 <= _GEN_4227[4:0]; // @[ivncontrol4.scala 18:{24,24}]
    i_vn2_3 <= _GEN_4228[4:0]; // @[ivncontrol4.scala 18:{24,24}]
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_0 <= io_Stationary_matrix_0_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_1 <= io_Stationary_matrix_0_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_2 <= io_Stationary_matrix_0_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_3 <= io_Stationary_matrix_0_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_4 <= io_Stationary_matrix_0_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_5 <= io_Stationary_matrix_0_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_6 <= io_Stationary_matrix_0_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_7 <= io_Stationary_matrix_0_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_0 <= io_Stationary_matrix_1_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_1 <= io_Stationary_matrix_1_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_2 <= io_Stationary_matrix_1_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_3 <= io_Stationary_matrix_1_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_4 <= io_Stationary_matrix_1_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_5 <= io_Stationary_matrix_1_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_6 <= io_Stationary_matrix_1_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_7 <= io_Stationary_matrix_1_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_0 <= io_Stationary_matrix_2_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_1 <= io_Stationary_matrix_2_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_2 <= io_Stationary_matrix_2_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_3 <= io_Stationary_matrix_2_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_4 <= io_Stationary_matrix_2_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_5 <= io_Stationary_matrix_2_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_6 <= io_Stationary_matrix_2_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_7 <= io_Stationary_matrix_2_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_0 <= io_Stationary_matrix_3_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_1 <= io_Stationary_matrix_3_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_2 <= io_Stationary_matrix_3_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_3 <= io_Stationary_matrix_3_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_4 <= io_Stationary_matrix_3_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_5 <= io_Stationary_matrix_3_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_6 <= io_Stationary_matrix_3_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_7 <= io_Stationary_matrix_3_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_0 <= io_Stationary_matrix_4_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_1 <= io_Stationary_matrix_4_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_2 <= io_Stationary_matrix_4_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_3 <= io_Stationary_matrix_4_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_4 <= io_Stationary_matrix_4_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_5 <= io_Stationary_matrix_4_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_6 <= io_Stationary_matrix_4_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_7 <= io_Stationary_matrix_4_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_0 <= io_Stationary_matrix_5_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_1 <= io_Stationary_matrix_5_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_2 <= io_Stationary_matrix_5_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_3 <= io_Stationary_matrix_5_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_4 <= io_Stationary_matrix_5_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_5 <= io_Stationary_matrix_5_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_6 <= io_Stationary_matrix_5_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_7 <= io_Stationary_matrix_5_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_0 <= io_Stationary_matrix_6_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_1 <= io_Stationary_matrix_6_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_2 <= io_Stationary_matrix_6_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_3 <= io_Stationary_matrix_6_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_4 <= io_Stationary_matrix_6_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_5 <= io_Stationary_matrix_6_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_6 <= io_Stationary_matrix_6_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_7 <= io_Stationary_matrix_6_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_0 <= io_Stationary_matrix_7_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_1 <= io_Stationary_matrix_7_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_2 <= io_Stationary_matrix_7_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_3 <= io_Stationary_matrix_7_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_4 <= io_Stationary_matrix_7_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_5 <= io_Stationary_matrix_7_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_6 <= io_Stationary_matrix_7_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_7 <= io_Stationary_matrix_7_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_0 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_0 <= count_0; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_1 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_1 <= count_1; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_2 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_2 <= count_2; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_3 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_3 <= count_3; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_4 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_4 <= count_4; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_5 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_5 <= count_5; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_6 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_6 <= count_6; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_7 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_7 <= count_7; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_8 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_8 <= 32'h0; // @[ivncontrol4.scala 87:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_9 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_9 <= 32'h0; // @[ivncontrol4.scala 87:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_10 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_10 <= 32'h0; // @[ivncontrol4.scala 87:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_11 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_11 <= 32'h0; // @[ivncontrol4.scala 87:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_12 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_12 <= 32'h0; // @[ivncontrol4.scala 87:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_13 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_13 <= 32'h0; // @[ivncontrol4.scala 87:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_14 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_14 <= 32'h0; // @[ivncontrol4.scala 87:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_15 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end
    if (reset) begin // @[ivncontrol4.scala 37:22]
      pin <= 32'h0; // @[ivncontrol4.scala 37:22]
    end else if (_T_72 & rowcount_6 == 32'h0 & rowcount_7 != 32'h0) begin // @[ivncontrol4.scala 183:192]
      pin <= 32'h7; // @[ivncontrol4.scala 184:13]
    end else if (_T_59 & rowcount_5 == 32'h0 & rowcount_6 != 32'h0) begin // @[ivncontrol4.scala 180:169]
      pin <= 32'h6; // @[ivncontrol4.scala 181:13]
    end else if (_T_48 & rowcount_4 == 32'h0 & rowcount_5 != 32'h0) begin // @[ivncontrol4.scala 177:146]
      pin <= 32'h5; // @[ivncontrol4.scala 178:13]
    end else begin
      pin <= _GEN_317;
    end
    if (reset) begin // @[ivncontrol4.scala 41:20]
      i <= 32'h0; // @[ivncontrol4.scala 41:20]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
        i <= _GEN_247;
      end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
        i <= _GEN_247;
      end else begin
        i <= _GEN_265;
      end
    end
    if (reset) begin // @[ivncontrol4.scala 42:20]
      j <= 32'h0; // @[ivncontrol4.scala 42:20]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
        j <= 32'h8; // @[ivncontrol4.scala 116:11]
      end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
        j <= _j_T_1; // @[ivncontrol4.scala 118:11]
      end else begin
        j <= {{28'd0}, _GEN_264};
      end
    end
    if (3'h0 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h0 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h0 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h0 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h0 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h0 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h0 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h0 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_0 <= _GEN_224;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_0 <= _GEN_224;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h0 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_0 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_0 <= _GEN_224;
      end
    end else begin
      count_0 <= _GEN_224;
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_1 <= _GEN_225;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_1 <= _GEN_225;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h1 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_1 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_1 <= _GEN_225;
      end
    end else begin
      count_1 <= _GEN_225;
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_2 <= _GEN_226;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_2 <= _GEN_226;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h2 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_2 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_2 <= _GEN_226;
      end
    end else begin
      count_2 <= _GEN_226;
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_3 <= _GEN_227;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_3 <= _GEN_227;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h3 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_3 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_3 <= _GEN_227;
      end
    end else begin
      count_3 <= _GEN_227;
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_4 <= _GEN_228;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_4 <= _GEN_228;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h4 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_4 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_4 <= _GEN_228;
      end
    end else begin
      count_4 <= _GEN_228;
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_5 <= _GEN_229;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_5 <= _GEN_229;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h5 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_5 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_5 <= _GEN_229;
      end
    end else begin
      count_5 <= _GEN_229;
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_6 <= _GEN_230;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_6 <= _GEN_230;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h6 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_6 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_6 <= _GEN_230;
      end
    end else begin
      count_6 <= _GEN_230;
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_7 <= _GEN_231;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_7 <= _GEN_231;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h7 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_7 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_7 <= _GEN_231;
      end
    end else begin
      count_7 <= _GEN_231;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  i_vn_0 = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  i_vn_1 = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  i_vn_2 = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  i_vn_3 = _RAND_3[4:0];
  _RAND_4 = {1{`RANDOM}};
  i_vn2_0 = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  i_vn2_1 = _RAND_5[4:0];
  _RAND_6 = {1{`RANDOM}};
  i_vn2_2 = _RAND_6[4:0];
  _RAND_7 = {1{`RANDOM}};
  i_vn2_3 = _RAND_7[4:0];
  _RAND_8 = {1{`RANDOM}};
  solution_0_0 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  solution_0_1 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  solution_0_2 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  solution_0_3 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  solution_0_4 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  solution_0_5 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  solution_0_6 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  solution_0_7 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  solution_1_0 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  solution_1_1 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  solution_1_2 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  solution_1_3 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  solution_1_4 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  solution_1_5 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  solution_1_6 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  solution_1_7 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  solution_2_0 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  solution_2_1 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  solution_2_2 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  solution_2_3 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  solution_2_4 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  solution_2_5 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  solution_2_6 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  solution_2_7 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  solution_3_0 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  solution_3_1 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  solution_3_2 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  solution_3_3 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  solution_3_4 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  solution_3_5 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  solution_3_6 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  solution_3_7 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  solution_4_0 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  solution_4_1 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  solution_4_2 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  solution_4_3 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  solution_4_4 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  solution_4_5 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  solution_4_6 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  solution_4_7 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  solution_5_0 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  solution_5_1 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  solution_5_2 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  solution_5_3 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  solution_5_4 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  solution_5_5 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  solution_5_6 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  solution_5_7 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  solution_6_0 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  solution_6_1 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  solution_6_2 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  solution_6_3 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  solution_6_4 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  solution_6_5 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  solution_6_6 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  solution_6_7 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  solution_7_0 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  solution_7_1 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  solution_7_2 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  solution_7_3 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  solution_7_4 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  solution_7_5 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  solution_7_6 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  solution_7_7 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  rowcount_0 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  rowcount_1 = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  rowcount_2 = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  rowcount_3 = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  rowcount_4 = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  rowcount_5 = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  rowcount_6 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  rowcount_7 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  rowcount_8 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  rowcount_9 = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  rowcount_10 = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  rowcount_11 = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  rowcount_12 = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  rowcount_13 = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  rowcount_14 = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  rowcount_15 = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  pin = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  i = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  j = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  mat_0_0 = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  mat_0_1 = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  mat_0_2 = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  mat_0_3 = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  mat_0_4 = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  mat_0_5 = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  mat_0_6 = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  mat_0_7 = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  mat_1_0 = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  mat_1_1 = _RAND_100[31:0];
  _RAND_101 = {1{`RANDOM}};
  mat_1_2 = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  mat_1_3 = _RAND_102[31:0];
  _RAND_103 = {1{`RANDOM}};
  mat_1_4 = _RAND_103[31:0];
  _RAND_104 = {1{`RANDOM}};
  mat_1_5 = _RAND_104[31:0];
  _RAND_105 = {1{`RANDOM}};
  mat_1_6 = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  mat_1_7 = _RAND_106[31:0];
  _RAND_107 = {1{`RANDOM}};
  mat_2_0 = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  mat_2_1 = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  mat_2_2 = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  mat_2_3 = _RAND_110[31:0];
  _RAND_111 = {1{`RANDOM}};
  mat_2_4 = _RAND_111[31:0];
  _RAND_112 = {1{`RANDOM}};
  mat_2_5 = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  mat_2_6 = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  mat_2_7 = _RAND_114[31:0];
  _RAND_115 = {1{`RANDOM}};
  mat_3_0 = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  mat_3_1 = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  mat_3_2 = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  mat_3_3 = _RAND_118[31:0];
  _RAND_119 = {1{`RANDOM}};
  mat_3_4 = _RAND_119[31:0];
  _RAND_120 = {1{`RANDOM}};
  mat_3_5 = _RAND_120[31:0];
  _RAND_121 = {1{`RANDOM}};
  mat_3_6 = _RAND_121[31:0];
  _RAND_122 = {1{`RANDOM}};
  mat_3_7 = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  mat_4_0 = _RAND_123[31:0];
  _RAND_124 = {1{`RANDOM}};
  mat_4_1 = _RAND_124[31:0];
  _RAND_125 = {1{`RANDOM}};
  mat_4_2 = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  mat_4_3 = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  mat_4_4 = _RAND_127[31:0];
  _RAND_128 = {1{`RANDOM}};
  mat_4_5 = _RAND_128[31:0];
  _RAND_129 = {1{`RANDOM}};
  mat_4_6 = _RAND_129[31:0];
  _RAND_130 = {1{`RANDOM}};
  mat_4_7 = _RAND_130[31:0];
  _RAND_131 = {1{`RANDOM}};
  mat_5_0 = _RAND_131[31:0];
  _RAND_132 = {1{`RANDOM}};
  mat_5_1 = _RAND_132[31:0];
  _RAND_133 = {1{`RANDOM}};
  mat_5_2 = _RAND_133[31:0];
  _RAND_134 = {1{`RANDOM}};
  mat_5_3 = _RAND_134[31:0];
  _RAND_135 = {1{`RANDOM}};
  mat_5_4 = _RAND_135[31:0];
  _RAND_136 = {1{`RANDOM}};
  mat_5_5 = _RAND_136[31:0];
  _RAND_137 = {1{`RANDOM}};
  mat_5_6 = _RAND_137[31:0];
  _RAND_138 = {1{`RANDOM}};
  mat_5_7 = _RAND_138[31:0];
  _RAND_139 = {1{`RANDOM}};
  mat_6_0 = _RAND_139[31:0];
  _RAND_140 = {1{`RANDOM}};
  mat_6_1 = _RAND_140[31:0];
  _RAND_141 = {1{`RANDOM}};
  mat_6_2 = _RAND_141[31:0];
  _RAND_142 = {1{`RANDOM}};
  mat_6_3 = _RAND_142[31:0];
  _RAND_143 = {1{`RANDOM}};
  mat_6_4 = _RAND_143[31:0];
  _RAND_144 = {1{`RANDOM}};
  mat_6_5 = _RAND_144[31:0];
  _RAND_145 = {1{`RANDOM}};
  mat_6_6 = _RAND_145[31:0];
  _RAND_146 = {1{`RANDOM}};
  mat_6_7 = _RAND_146[31:0];
  _RAND_147 = {1{`RANDOM}};
  mat_7_0 = _RAND_147[31:0];
  _RAND_148 = {1{`RANDOM}};
  mat_7_1 = _RAND_148[31:0];
  _RAND_149 = {1{`RANDOM}};
  mat_7_2 = _RAND_149[31:0];
  _RAND_150 = {1{`RANDOM}};
  mat_7_3 = _RAND_150[31:0];
  _RAND_151 = {1{`RANDOM}};
  mat_7_4 = _RAND_151[31:0];
  _RAND_152 = {1{`RANDOM}};
  mat_7_5 = _RAND_152[31:0];
  _RAND_153 = {1{`RANDOM}};
  mat_7_6 = _RAND_153[31:0];
  _RAND_154 = {1{`RANDOM}};
  mat_7_7 = _RAND_154[31:0];
  _RAND_155 = {1{`RANDOM}};
  count_0 = _RAND_155[31:0];
  _RAND_156 = {1{`RANDOM}};
  count_1 = _RAND_156[31:0];
  _RAND_157 = {1{`RANDOM}};
  count_2 = _RAND_157[31:0];
  _RAND_158 = {1{`RANDOM}};
  count_3 = _RAND_158[31:0];
  _RAND_159 = {1{`RANDOM}};
  count_4 = _RAND_159[31:0];
  _RAND_160 = {1{`RANDOM}};
  count_5 = _RAND_160[31:0];
  _RAND_161 = {1{`RANDOM}};
  count_6 = _RAND_161[31:0];
  _RAND_162 = {1{`RANDOM}};
  count_7 = _RAND_162[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ivncontrol4_1(
  input         clock,
  input         reset,
  input  [15:0] io_Stationary_matrix_0_0,
  input  [15:0] io_Stationary_matrix_0_1,
  input  [15:0] io_Stationary_matrix_0_2,
  input  [15:0] io_Stationary_matrix_0_3,
  input  [15:0] io_Stationary_matrix_0_4,
  input  [15:0] io_Stationary_matrix_0_5,
  input  [15:0] io_Stationary_matrix_0_6,
  input  [15:0] io_Stationary_matrix_0_7,
  input  [15:0] io_Stationary_matrix_1_0,
  input  [15:0] io_Stationary_matrix_1_1,
  input  [15:0] io_Stationary_matrix_1_2,
  input  [15:0] io_Stationary_matrix_1_3,
  input  [15:0] io_Stationary_matrix_1_4,
  input  [15:0] io_Stationary_matrix_1_5,
  input  [15:0] io_Stationary_matrix_1_6,
  input  [15:0] io_Stationary_matrix_1_7,
  input  [15:0] io_Stationary_matrix_2_0,
  input  [15:0] io_Stationary_matrix_2_1,
  input  [15:0] io_Stationary_matrix_2_2,
  input  [15:0] io_Stationary_matrix_2_3,
  input  [15:0] io_Stationary_matrix_2_4,
  input  [15:0] io_Stationary_matrix_2_5,
  input  [15:0] io_Stationary_matrix_2_6,
  input  [15:0] io_Stationary_matrix_2_7,
  input  [15:0] io_Stationary_matrix_3_0,
  input  [15:0] io_Stationary_matrix_3_1,
  input  [15:0] io_Stationary_matrix_3_2,
  input  [15:0] io_Stationary_matrix_3_3,
  input  [15:0] io_Stationary_matrix_3_4,
  input  [15:0] io_Stationary_matrix_3_5,
  input  [15:0] io_Stationary_matrix_3_6,
  input  [15:0] io_Stationary_matrix_3_7,
  input  [15:0] io_Stationary_matrix_4_0,
  input  [15:0] io_Stationary_matrix_4_1,
  input  [15:0] io_Stationary_matrix_4_2,
  input  [15:0] io_Stationary_matrix_4_3,
  input  [15:0] io_Stationary_matrix_4_4,
  input  [15:0] io_Stationary_matrix_4_5,
  input  [15:0] io_Stationary_matrix_4_6,
  input  [15:0] io_Stationary_matrix_4_7,
  input  [15:0] io_Stationary_matrix_5_0,
  input  [15:0] io_Stationary_matrix_5_1,
  input  [15:0] io_Stationary_matrix_5_2,
  input  [15:0] io_Stationary_matrix_5_3,
  input  [15:0] io_Stationary_matrix_5_4,
  input  [15:0] io_Stationary_matrix_5_5,
  input  [15:0] io_Stationary_matrix_5_6,
  input  [15:0] io_Stationary_matrix_5_7,
  input  [15:0] io_Stationary_matrix_6_0,
  input  [15:0] io_Stationary_matrix_6_1,
  input  [15:0] io_Stationary_matrix_6_2,
  input  [15:0] io_Stationary_matrix_6_3,
  input  [15:0] io_Stationary_matrix_6_4,
  input  [15:0] io_Stationary_matrix_6_5,
  input  [15:0] io_Stationary_matrix_6_6,
  input  [15:0] io_Stationary_matrix_6_7,
  input  [15:0] io_Stationary_matrix_7_0,
  input  [15:0] io_Stationary_matrix_7_1,
  input  [15:0] io_Stationary_matrix_7_2,
  input  [15:0] io_Stationary_matrix_7_3,
  input  [15:0] io_Stationary_matrix_7_4,
  input  [15:0] io_Stationary_matrix_7_5,
  input  [15:0] io_Stationary_matrix_7_6,
  input  [15:0] io_Stationary_matrix_7_7,
  output [4:0]  io_o_vn_0,
  output [4:0]  io_o_vn_1,
  output [4:0]  io_o_vn_2,
  output [4:0]  io_o_vn_3,
  output [4:0]  io_o_vn2_0,
  output [4:0]  io_o_vn2_1,
  output [4:0]  io_o_vn2_2,
  output [4:0]  io_o_vn2_3,
  input         io_validpin
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
`endif // RANDOMIZE_REG_INIT
  reg [4:0] i_vn_0; // @[ivncontrol4.scala 17:23]
  reg [4:0] i_vn_1; // @[ivncontrol4.scala 17:23]
  reg [4:0] i_vn_2; // @[ivncontrol4.scala 17:23]
  reg [4:0] i_vn_3; // @[ivncontrol4.scala 17:23]
  reg [4:0] i_vn2_0; // @[ivncontrol4.scala 18:24]
  reg [4:0] i_vn2_1; // @[ivncontrol4.scala 18:24]
  reg [4:0] i_vn2_2; // @[ivncontrol4.scala 18:24]
  reg [4:0] i_vn2_3; // @[ivncontrol4.scala 18:24]
  reg [15:0] solution_0_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_0_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_0_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_0_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_0_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_0_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_0_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_0_7; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_7; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_7; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_7; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_7; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_7; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_7; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_7; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_0; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_1; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_2; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_3; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_4; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_5; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_6; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_7; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_8; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_9; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_10; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_11; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_12; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_13; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_14; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_15; // @[ivncontrol4.scala 27:27]
  reg [31:0] pin; // @[ivncontrol4.scala 37:22]
  reg [31:0] i; // @[ivncontrol4.scala 41:20]
  reg [31:0] j; // @[ivncontrol4.scala 42:20]
  wire  _io_ProcessValid_T = i == 32'h7; // @[ivncontrol4.scala 44:27]
  wire  _io_ProcessValid_T_1 = j == 32'h7; // @[ivncontrol4.scala 44:42]
  wire  _io_ProcessValid_T_2 = i == 32'h7 & j == 32'h7; // @[ivncontrol4.scala 44:36]
  reg [31:0] mat_0_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_0_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_0_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_0_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_0_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_0_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_0_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_0_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] count_0; // @[ivncontrol4.scala 58:20]
  reg [31:0] count_1; // @[ivncontrol4.scala 58:20]
  reg [31:0] count_2; // @[ivncontrol4.scala 58:20]
  reg [31:0] count_3; // @[ivncontrol4.scala 58:20]
  reg [31:0] count_4; // @[ivncontrol4.scala 58:20]
  reg [31:0] count_5; // @[ivncontrol4.scala 58:20]
  reg [31:0] count_6; // @[ivncontrol4.scala 58:20]
  reg [31:0] count_7; // @[ivncontrol4.scala 58:20]
  wire  _GEN_3825 = 3'h0 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_65 = 3'h0 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_0_1 : io_Stationary_matrix_0_0; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_66 = 3'h0 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_0_2 : _GEN_65; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_67 = 3'h0 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_0_3 : _GEN_66; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_68 = 3'h0 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_0_4 : _GEN_67; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_69 = 3'h0 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_0_5 : _GEN_68; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_70 = 3'h0 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_0_6 : _GEN_69; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_71 = 3'h0 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_0_7 : _GEN_70; // @[ivncontrol4.scala 63:{17,17}]
  wire  _GEN_3839 = 3'h1 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_72 = 3'h1 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_1_0 : _GEN_71; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_73 = 3'h1 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_1_1 : _GEN_72; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_74 = 3'h1 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_1_2 : _GEN_73; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_75 = 3'h1 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_1_3 : _GEN_74; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_76 = 3'h1 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_1_4 : _GEN_75; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_77 = 3'h1 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_1_5 : _GEN_76; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_78 = 3'h1 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_1_6 : _GEN_77; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_79 = 3'h1 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_1_7 : _GEN_78; // @[ivncontrol4.scala 63:{17,17}]
  wire  _GEN_3855 = 3'h2 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_80 = 3'h2 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_2_0 : _GEN_79; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_81 = 3'h2 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_2_1 : _GEN_80; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_82 = 3'h2 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_2_2 : _GEN_81; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_83 = 3'h2 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_2_3 : _GEN_82; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_84 = 3'h2 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_2_4 : _GEN_83; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_85 = 3'h2 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_2_5 : _GEN_84; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_86 = 3'h2 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_2_6 : _GEN_85; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_87 = 3'h2 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_2_7 : _GEN_86; // @[ivncontrol4.scala 63:{17,17}]
  wire  _GEN_3871 = 3'h3 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_88 = 3'h3 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_3_0 : _GEN_87; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_89 = 3'h3 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_3_1 : _GEN_88; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_90 = 3'h3 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_3_2 : _GEN_89; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_91 = 3'h3 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_3_3 : _GEN_90; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_92 = 3'h3 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_3_4 : _GEN_91; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_93 = 3'h3 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_3_5 : _GEN_92; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_94 = 3'h3 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_3_6 : _GEN_93; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_95 = 3'h3 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_3_7 : _GEN_94; // @[ivncontrol4.scala 63:{17,17}]
  wire  _GEN_3887 = 3'h4 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_96 = 3'h4 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_4_0 : _GEN_95; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_97 = 3'h4 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_4_1 : _GEN_96; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_98 = 3'h4 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_4_2 : _GEN_97; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_99 = 3'h4 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_4_3 : _GEN_98; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_100 = 3'h4 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_4_4 : _GEN_99; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_101 = 3'h4 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_4_5 : _GEN_100; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_102 = 3'h4 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_4_6 : _GEN_101; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_103 = 3'h4 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_4_7 : _GEN_102; // @[ivncontrol4.scala 63:{17,17}]
  wire  _GEN_3903 = 3'h5 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_104 = 3'h5 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_5_0 : _GEN_103; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_105 = 3'h5 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_5_1 : _GEN_104; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_106 = 3'h5 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_5_2 : _GEN_105; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_107 = 3'h5 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_5_3 : _GEN_106; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_108 = 3'h5 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_5_4 : _GEN_107; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_109 = 3'h5 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_5_5 : _GEN_108; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_110 = 3'h5 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_5_6 : _GEN_109; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_111 = 3'h5 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_5_7 : _GEN_110; // @[ivncontrol4.scala 63:{17,17}]
  wire  _GEN_3919 = 3'h6 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_112 = 3'h6 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_6_0 : _GEN_111; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_113 = 3'h6 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_6_1 : _GEN_112; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_114 = 3'h6 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_6_2 : _GEN_113; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_115 = 3'h6 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_6_3 : _GEN_114; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_116 = 3'h6 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_6_4 : _GEN_115; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_117 = 3'h6 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_6_5 : _GEN_116; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_118 = 3'h6 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_6_6 : _GEN_117; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_119 = 3'h6 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_6_7 : _GEN_118; // @[ivncontrol4.scala 63:{17,17}]
  wire  _GEN_3935 = 3'h7 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_120 = 3'h7 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_7_0 : _GEN_119; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_121 = 3'h7 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_7_1 : _GEN_120; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_122 = 3'h7 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_7_2 : _GEN_121; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_123 = 3'h7 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_7_3 : _GEN_122; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_124 = 3'h7 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_7_4 : _GEN_123; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_125 = 3'h7 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_7_5 : _GEN_124; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_126 = 3'h7 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_7_6 : _GEN_125; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_127 = 3'h7 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_7_7 : _GEN_126; // @[ivncontrol4.scala 63:{17,17}]
  wire [31:0] _mat_T_1_T_2 = {{16'd0}, _GEN_127}; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_129 = _GEN_3825 & 4'h1 == j[3:0] ? solution_0_1 : solution_0_0; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_130 = _GEN_3825 & 4'h2 == j[3:0] ? solution_0_2 : _GEN_129; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_131 = _GEN_3825 & 4'h3 == j[3:0] ? solution_0_3 : _GEN_130; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_132 = _GEN_3825 & 4'h4 == j[3:0] ? solution_0_4 : _GEN_131; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_133 = _GEN_3825 & 4'h5 == j[3:0] ? solution_0_5 : _GEN_132; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_134 = _GEN_3825 & 4'h6 == j[3:0] ? solution_0_6 : _GEN_133; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_135 = _GEN_3825 & 4'h7 == j[3:0] ? solution_0_7 : _GEN_134; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_136 = _GEN_3825 & 4'h8 == j[3:0] ? 16'h0 : _GEN_135; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_137 = _GEN_3839 & 4'h0 == j[3:0] ? solution_1_0 : _GEN_136; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_138 = _GEN_3839 & 4'h1 == j[3:0] ? solution_1_1 : _GEN_137; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_139 = _GEN_3839 & 4'h2 == j[3:0] ? solution_1_2 : _GEN_138; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_140 = _GEN_3839 & 4'h3 == j[3:0] ? solution_1_3 : _GEN_139; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_141 = _GEN_3839 & 4'h4 == j[3:0] ? solution_1_4 : _GEN_140; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_142 = _GEN_3839 & 4'h5 == j[3:0] ? solution_1_5 : _GEN_141; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_143 = _GEN_3839 & 4'h6 == j[3:0] ? solution_1_6 : _GEN_142; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_144 = _GEN_3839 & 4'h7 == j[3:0] ? solution_1_7 : _GEN_143; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_145 = _GEN_3839 & 4'h8 == j[3:0] ? 16'h0 : _GEN_144; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_146 = _GEN_3855 & 4'h0 == j[3:0] ? solution_2_0 : _GEN_145; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_147 = _GEN_3855 & 4'h1 == j[3:0] ? solution_2_1 : _GEN_146; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_148 = _GEN_3855 & 4'h2 == j[3:0] ? solution_2_2 : _GEN_147; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_149 = _GEN_3855 & 4'h3 == j[3:0] ? solution_2_3 : _GEN_148; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_150 = _GEN_3855 & 4'h4 == j[3:0] ? solution_2_4 : _GEN_149; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_151 = _GEN_3855 & 4'h5 == j[3:0] ? solution_2_5 : _GEN_150; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_152 = _GEN_3855 & 4'h6 == j[3:0] ? solution_2_6 : _GEN_151; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_153 = _GEN_3855 & 4'h7 == j[3:0] ? solution_2_7 : _GEN_152; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_154 = _GEN_3855 & 4'h8 == j[3:0] ? 16'h0 : _GEN_153; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_155 = _GEN_3871 & 4'h0 == j[3:0] ? solution_3_0 : _GEN_154; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_156 = _GEN_3871 & 4'h1 == j[3:0] ? solution_3_1 : _GEN_155; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_157 = _GEN_3871 & 4'h2 == j[3:0] ? solution_3_2 : _GEN_156; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_158 = _GEN_3871 & 4'h3 == j[3:0] ? solution_3_3 : _GEN_157; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_159 = _GEN_3871 & 4'h4 == j[3:0] ? solution_3_4 : _GEN_158; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_160 = _GEN_3871 & 4'h5 == j[3:0] ? solution_3_5 : _GEN_159; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_161 = _GEN_3871 & 4'h6 == j[3:0] ? solution_3_6 : _GEN_160; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_162 = _GEN_3871 & 4'h7 == j[3:0] ? solution_3_7 : _GEN_161; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_163 = _GEN_3871 & 4'h8 == j[3:0] ? 16'h0 : _GEN_162; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_164 = _GEN_3887 & 4'h0 == j[3:0] ? solution_4_0 : _GEN_163; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_165 = _GEN_3887 & 4'h1 == j[3:0] ? solution_4_1 : _GEN_164; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_166 = _GEN_3887 & 4'h2 == j[3:0] ? solution_4_2 : _GEN_165; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_167 = _GEN_3887 & 4'h3 == j[3:0] ? solution_4_3 : _GEN_166; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_168 = _GEN_3887 & 4'h4 == j[3:0] ? solution_4_4 : _GEN_167; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_169 = _GEN_3887 & 4'h5 == j[3:0] ? solution_4_5 : _GEN_168; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_170 = _GEN_3887 & 4'h6 == j[3:0] ? solution_4_6 : _GEN_169; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_171 = _GEN_3887 & 4'h7 == j[3:0] ? solution_4_7 : _GEN_170; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_172 = _GEN_3887 & 4'h8 == j[3:0] ? 16'h0 : _GEN_171; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_173 = _GEN_3903 & 4'h0 == j[3:0] ? solution_5_0 : _GEN_172; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_174 = _GEN_3903 & 4'h1 == j[3:0] ? solution_5_1 : _GEN_173; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_175 = _GEN_3903 & 4'h2 == j[3:0] ? solution_5_2 : _GEN_174; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_176 = _GEN_3903 & 4'h3 == j[3:0] ? solution_5_3 : _GEN_175; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_177 = _GEN_3903 & 4'h4 == j[3:0] ? solution_5_4 : _GEN_176; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_178 = _GEN_3903 & 4'h5 == j[3:0] ? solution_5_5 : _GEN_177; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_179 = _GEN_3903 & 4'h6 == j[3:0] ? solution_5_6 : _GEN_178; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_180 = _GEN_3903 & 4'h7 == j[3:0] ? solution_5_7 : _GEN_179; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_181 = _GEN_3903 & 4'h8 == j[3:0] ? 16'h0 : _GEN_180; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_182 = _GEN_3919 & 4'h0 == j[3:0] ? solution_6_0 : _GEN_181; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_183 = _GEN_3919 & 4'h1 == j[3:0] ? solution_6_1 : _GEN_182; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_184 = _GEN_3919 & 4'h2 == j[3:0] ? solution_6_2 : _GEN_183; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_185 = _GEN_3919 & 4'h3 == j[3:0] ? solution_6_3 : _GEN_184; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_186 = _GEN_3919 & 4'h4 == j[3:0] ? solution_6_4 : _GEN_185; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_187 = _GEN_3919 & 4'h5 == j[3:0] ? solution_6_5 : _GEN_186; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_188 = _GEN_3919 & 4'h6 == j[3:0] ? solution_6_6 : _GEN_187; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_189 = _GEN_3919 & 4'h7 == j[3:0] ? solution_6_7 : _GEN_188; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_190 = _GEN_3919 & 4'h8 == j[3:0] ? 16'h0 : _GEN_189; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_191 = _GEN_3935 & 4'h0 == j[3:0] ? solution_7_0 : _GEN_190; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_192 = _GEN_3935 & 4'h1 == j[3:0] ? solution_7_1 : _GEN_191; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_193 = _GEN_3935 & 4'h2 == j[3:0] ? solution_7_2 : _GEN_192; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_194 = _GEN_3935 & 4'h3 == j[3:0] ? solution_7_3 : _GEN_193; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_195 = _GEN_3935 & 4'h4 == j[3:0] ? solution_7_4 : _GEN_194; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_196 = _GEN_3935 & 4'h5 == j[3:0] ? solution_7_5 : _GEN_195; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_197 = _GEN_3935 & 4'h6 == j[3:0] ? solution_7_6 : _GEN_196; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_198 = _GEN_3935 & 4'h7 == j[3:0] ? solution_7_7 : _GEN_197; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_199 = _GEN_3935 & 4'h8 == j[3:0] ? 16'h0 : _GEN_198; // @[ivncontrol4.scala 65:{31,31}]
  wire [31:0] _GEN_201 = 3'h1 == i[2:0] ? count_1 : count_0; // @[ivncontrol4.scala 66:{33,33}]
  wire [31:0] _GEN_202 = 3'h2 == i[2:0] ? count_2 : _GEN_201; // @[ivncontrol4.scala 66:{33,33}]
  wire [31:0] _GEN_203 = 3'h3 == i[2:0] ? count_3 : _GEN_202; // @[ivncontrol4.scala 66:{33,33}]
  wire [31:0] _GEN_204 = 3'h4 == i[2:0] ? count_4 : _GEN_203; // @[ivncontrol4.scala 66:{33,33}]
  wire [31:0] _GEN_205 = 3'h5 == i[2:0] ? count_5 : _GEN_204; // @[ivncontrol4.scala 66:{33,33}]
  wire [31:0] _GEN_206 = 3'h6 == i[2:0] ? count_6 : _GEN_205; // @[ivncontrol4.scala 66:{33,33}]
  wire [31:0] _GEN_207 = 3'h7 == i[2:0] ? count_7 : _GEN_206; // @[ivncontrol4.scala 66:{33,33}]
  wire [31:0] _count_T_2 = _GEN_207 + 32'h1; // @[ivncontrol4.scala 66:33]
  wire [31:0] _GEN_208 = 3'h0 == i[2:0] ? _count_T_2 : count_0; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_209 = 3'h1 == i[2:0] ? _count_T_2 : count_1; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_210 = 3'h2 == i[2:0] ? _count_T_2 : count_2; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_211 = 3'h3 == i[2:0] ? _count_T_2 : count_3; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_212 = 3'h4 == i[2:0] ? _count_T_2 : count_4; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_213 = 3'h5 == i[2:0] ? _count_T_2 : count_5; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_214 = 3'h6 == i[2:0] ? _count_T_2 : count_6; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_215 = 3'h7 == i[2:0] ? _count_T_2 : count_7; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_216 = _GEN_199 != 16'h0 ? _GEN_208 : count_0; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_217 = _GEN_199 != 16'h0 ? _GEN_209 : count_1; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_218 = _GEN_199 != 16'h0 ? _GEN_210 : count_2; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_219 = _GEN_199 != 16'h0 ? _GEN_211 : count_3; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_220 = _GEN_199 != 16'h0 ? _GEN_212 : count_4; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_221 = _GEN_199 != 16'h0 ? _GEN_213 : count_5; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_222 = _GEN_199 != 16'h0 ? _GEN_214 : count_6; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_223 = _GEN_199 != 16'h0 ? _GEN_215 : count_7; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_224 = io_validpin ? _GEN_216 : count_0; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _GEN_225 = io_validpin ? _GEN_217 : count_1; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _GEN_226 = io_validpin ? _GEN_218 : count_2; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _GEN_227 = io_validpin ? _GEN_219 : count_3; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _GEN_228 = io_validpin ? _GEN_220 : count_4; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _GEN_229 = io_validpin ? _GEN_221 : count_5; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _GEN_230 = io_validpin ? _GEN_222 : count_6; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _GEN_231 = io_validpin ? _GEN_223 : count_7; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _i_T_1 = i + 32'h1; // @[ivncontrol4.scala 113:16]
  wire [31:0] _GEN_247 = i < 32'h7 & _io_ProcessValid_T_1 ? _i_T_1 : i; // @[ivncontrol4.scala 112:74 113:11 41:20]
  wire [31:0] _j_T_1 = j + 32'h1; // @[ivncontrol4.scala 118:16]
  wire [3:0] _GEN_264 = _io_ProcessValid_T & j == 32'h8 ? 4'h8 : 4'h0; // @[ivncontrol4.scala 120:77 121:11 129:11]
  wire [31:0] _GEN_265 = _io_ProcessValid_T & j == 32'h8 ? 32'h7 : _GEN_247; // @[ivncontrol4.scala 120:77 122:11]
  wire  _GEN_312 = _io_ProcessValid_T_2; // @[ivncontrol4.scala 153:41]
  wire [31:0] _GEN_313 = rowcount_0 != 32'h0 ? 32'h0 : pin; // @[ivncontrol4.scala 162:30 163:13 37:22]
  wire  _T_27 = rowcount_0 == 32'h0; // @[ivncontrol4.scala 165:23]
  wire [31:0] _GEN_314 = rowcount_0 == 32'h0 & rowcount_1 != 32'h0 ? 32'h1 : _GEN_313; // @[ivncontrol4.scala 165:54 166:13]
  wire  _T_32 = _T_27 & rowcount_1 == 32'h0; // @[ivncontrol4.scala 168:31]
  wire [31:0] _GEN_315 = _T_27 & rowcount_1 == 32'h0 & rowcount_2 != 32'h0 ? 32'h2 : _GEN_314; // @[ivncontrol4.scala 168:77 169:13]
  wire  _T_39 = _T_32 & rowcount_2 == 32'h0; // @[ivncontrol4.scala 171:54]
  wire [31:0] _GEN_316 = _T_32 & rowcount_2 == 32'h0 & rowcount_3 != 32'h0 ? 32'h3 : _GEN_315; // @[ivncontrol4.scala 171:100 172:13]
  wire  _T_48 = _T_39 & rowcount_3 == 32'h0; // @[ivncontrol4.scala 174:77]
  wire [31:0] _GEN_317 = _T_39 & rowcount_3 == 32'h0 & rowcount_4 != 32'h0 ? 32'h4 : _GEN_316; // @[ivncontrol4.scala 174:123 175:13]
  wire  _T_59 = _T_48 & rowcount_4 == 32'h0; // @[ivncontrol4.scala 177:100]
  wire  _T_72 = _T_59 & rowcount_5 == 32'h0; // @[ivncontrol4.scala 180:123]
  wire  valid = _io_ProcessValid_T_2; // @[ivncontrol4.scala 153:41]
  wire [32:0] _T_91 = {{1'd0}, pin}; // @[ivncontrol4.scala 191:27]
  wire [31:0] _GEN_322 = 4'h1 == _T_91[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_323 = 4'h2 == _T_91[3:0] ? rowcount_2 : _GEN_322; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_324 = 4'h3 == _T_91[3:0] ? rowcount_3 : _GEN_323; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_325 = 4'h4 == _T_91[3:0] ? rowcount_4 : _GEN_324; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_326 = 4'h5 == _T_91[3:0] ? rowcount_5 : _GEN_325; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_327 = 4'h6 == _T_91[3:0] ? rowcount_6 : _GEN_326; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_328 = 4'h7 == _T_91[3:0] ? rowcount_7 : _GEN_327; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_329 = 4'h8 == _T_91[3:0] ? rowcount_8 : _GEN_328; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_330 = 4'h9 == _T_91[3:0] ? rowcount_9 : _GEN_329; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_331 = 4'ha == _T_91[3:0] ? rowcount_10 : _GEN_330; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_332 = 4'hb == _T_91[3:0] ? rowcount_11 : _GEN_331; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_333 = 4'hc == _T_91[3:0] ? rowcount_12 : _GEN_332; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_334 = 4'hd == _T_91[3:0] ? rowcount_13 : _GEN_333; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_335 = 4'he == _T_91[3:0] ? rowcount_14 : _GEN_334; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_336 = 4'hf == _T_91[3:0] ? rowcount_15 : _GEN_335; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_449 = _GEN_336 == 32'h1 ? _T_91[31:0] : 32'h10; // @[ivncontrol4.scala 142:17 241:50 242:21]
  wire [31:0] _GEN_450 = _GEN_336 == 32'h2 ? _T_91[31:0] : _GEN_449; // @[ivncontrol4.scala 237:51 238:21]
  wire [31:0] _GEN_451 = _GEN_336 == 32'h2 ? _T_91[31:0] : 32'h8; // @[ivncontrol4.scala 142:17 237:51 239:21]
  wire [31:0] _GEN_452 = _GEN_336 == 32'h3 ? _T_91[31:0] : _GEN_450; // @[ivncontrol4.scala 232:50 233:21]
  wire [31:0] _GEN_453 = _GEN_336 == 32'h3 ? _T_91[31:0] : _GEN_451; // @[ivncontrol4.scala 232:50 234:21]
  wire [31:0] _GEN_454 = _GEN_336 == 32'h3 ? _T_91[31:0] : 32'ha; // @[ivncontrol4.scala 142:17 232:50 235:21]
  wire [31:0] _GEN_455 = _GEN_336 == 32'h4 ? _T_91[31:0] : _GEN_452; // @[ivncontrol4.scala 224:50 225:21]
  wire [31:0] _GEN_456 = _GEN_336 == 32'h4 ? _T_91[31:0] : _GEN_453; // @[ivncontrol4.scala 224:50 226:21]
  wire [31:0] _GEN_457 = _GEN_336 == 32'h4 ? _T_91[31:0] : _GEN_454; // @[ivncontrol4.scala 224:50 227:21]
  wire [31:0] _GEN_458 = _GEN_336 == 32'h4 ? _T_91[31:0] : 32'h5; // @[ivncontrol4.scala 142:17 224:50 228:21]
  wire [31:0] _GEN_459 = _GEN_336 == 32'h5 ? _T_91[31:0] : _GEN_455; // @[ivncontrol4.scala 217:50 218:21]
  wire [31:0] _GEN_460 = _GEN_336 == 32'h5 ? _T_91[31:0] : _GEN_456; // @[ivncontrol4.scala 217:50 219:21]
  wire [31:0] _GEN_461 = _GEN_336 == 32'h5 ? _T_91[31:0] : _GEN_457; // @[ivncontrol4.scala 217:50 220:21]
  wire [31:0] _GEN_462 = _GEN_336 == 32'h5 ? _T_91[31:0] : _GEN_458; // @[ivncontrol4.scala 217:50 221:21]
  wire [31:0] _GEN_463 = _GEN_336 == 32'h5 ? _T_91[31:0] : 32'h17; // @[ivncontrol4.scala 143:18 217:50 222:22]
  wire [31:0] _GEN_464 = _GEN_336 == 32'h6 ? _T_91[31:0] : _GEN_459; // @[ivncontrol4.scala 209:52 210:21]
  wire [31:0] _GEN_465 = _GEN_336 == 32'h6 ? _T_91[31:0] : _GEN_460; // @[ivncontrol4.scala 209:52 211:21]
  wire [31:0] _GEN_466 = _GEN_336 == 32'h6 ? _T_91[31:0] : _GEN_461; // @[ivncontrol4.scala 209:52 212:21]
  wire [31:0] _GEN_467 = _GEN_336 == 32'h6 ? _T_91[31:0] : _GEN_462; // @[ivncontrol4.scala 209:52 213:21]
  wire [31:0] _GEN_468 = _GEN_336 == 32'h6 ? _T_91[31:0] : _GEN_463; // @[ivncontrol4.scala 209:52 214:22]
  wire [31:0] _GEN_469 = _GEN_336 == 32'h6 ? _T_91[31:0] : 32'h14; // @[ivncontrol4.scala 143:18 209:52 215:22]
  wire [31:0] _GEN_470 = _GEN_336 == 32'h7 ? _T_91[31:0] : _GEN_464; // @[ivncontrol4.scala 201:52 202:21]
  wire [31:0] _GEN_471 = _GEN_336 == 32'h7 ? _T_91[31:0] : _GEN_465; // @[ivncontrol4.scala 201:52 203:21]
  wire [31:0] _GEN_472 = _GEN_336 == 32'h7 ? _T_91[31:0] : _GEN_466; // @[ivncontrol4.scala 201:52 204:21]
  wire [31:0] _GEN_473 = _GEN_336 == 32'h7 ? _T_91[31:0] : _GEN_467; // @[ivncontrol4.scala 201:52 205:21]
  wire [31:0] _GEN_474 = _GEN_336 == 32'h7 ? _T_91[31:0] : _GEN_468; // @[ivncontrol4.scala 201:52 206:22]
  wire [31:0] _GEN_475 = _GEN_336 == 32'h7 ? _T_91[31:0] : _GEN_469; // @[ivncontrol4.scala 201:52 207:22]
  wire [31:0] _GEN_476 = _GEN_336 == 32'h7 ? _T_91[31:0] : 32'h1; // @[ivncontrol4.scala 143:18 201:52 208:22]
  wire [31:0] _GEN_477 = _GEN_336 >= 32'h8 ? _T_91[31:0] : _GEN_470; // @[ivncontrol4.scala 191:42 192:21]
  wire [31:0] _GEN_478 = _GEN_336 >= 32'h8 ? _T_91[31:0] : _GEN_471; // @[ivncontrol4.scala 191:42 193:21]
  wire [31:0] _GEN_479 = _GEN_336 >= 32'h8 ? _T_91[31:0] : _GEN_472; // @[ivncontrol4.scala 191:42 194:21]
  wire [31:0] _GEN_480 = _GEN_336 >= 32'h8 ? _T_91[31:0] : _GEN_473; // @[ivncontrol4.scala 191:42 195:21]
  wire [31:0] _GEN_481 = _GEN_336 >= 32'h8 ? _T_91[31:0] : _GEN_474; // @[ivncontrol4.scala 191:42 196:22]
  wire [31:0] _GEN_482 = _GEN_336 >= 32'h8 ? _T_91[31:0] : _GEN_475; // @[ivncontrol4.scala 191:42 197:22]
  wire [31:0] _GEN_483 = _GEN_336 >= 32'h8 ? _T_91[31:0] : _GEN_476; // @[ivncontrol4.scala 191:42 198:22]
  wire [31:0] _GEN_484 = _GEN_336 >= 32'h8 ? _T_91[31:0] : 32'hc; // @[ivncontrol4.scala 143:18 191:42 199:22]
  wire [31:0] _T_127 = 32'h8 - _GEN_336; // @[ivncontrol4.scala 245:18]
  wire [31:0] _i_vn_1_T_15 = 32'h1 + pin; // @[ivncontrol4.scala 246:29]
  wire [31:0] _GEN_597 = _T_127 == 32'h1 ? _i_vn_1_T_15 : _GEN_484; // @[ivncontrol4.scala 286:54 289:22]
  wire [31:0] _GEN_598 = _T_127 == 32'h2 ? _i_vn_1_T_15 : _GEN_483; // @[ivncontrol4.scala 281:54 284:22]
  wire [31:0] _GEN_599 = _T_127 == 32'h2 ? _i_vn_1_T_15 : _GEN_597; // @[ivncontrol4.scala 281:54 285:22]
  wire [31:0] _GEN_600 = _T_127 == 32'h3 ? _i_vn_1_T_15 : _GEN_482; // @[ivncontrol4.scala 274:54 276:22]
  wire [31:0] _GEN_601 = _T_127 == 32'h3 ? _i_vn_1_T_15 : _GEN_598; // @[ivncontrol4.scala 274:54 277:22]
  wire [31:0] _GEN_602 = _T_127 == 32'h3 ? _i_vn_1_T_15 : _GEN_599; // @[ivncontrol4.scala 274:54 278:22]
  wire [31:0] _GEN_603 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_481; // @[ivncontrol4.scala 268:54 270:22]
  wire [31:0] _GEN_604 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_600; // @[ivncontrol4.scala 268:54 271:22]
  wire [31:0] _GEN_605 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_601; // @[ivncontrol4.scala 268:54 272:22]
  wire [31:0] _GEN_606 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_602; // @[ivncontrol4.scala 268:54 273:22]
  wire [31:0] _GEN_607 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_480; // @[ivncontrol4.scala 261:54 263:21]
  wire [31:0] _GEN_608 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_603; // @[ivncontrol4.scala 261:54 264:22]
  wire [31:0] _GEN_609 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_604; // @[ivncontrol4.scala 261:54 265:22]
  wire [31:0] _GEN_610 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_605; // @[ivncontrol4.scala 261:54 266:22]
  wire [31:0] _GEN_611 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_606; // @[ivncontrol4.scala 261:54 267:22]
  wire [31:0] _GEN_612 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_479; // @[ivncontrol4.scala 254:54 255:22]
  wire [31:0] _GEN_613 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_607; // @[ivncontrol4.scala 254:54 256:21]
  wire [31:0] _GEN_614 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_608; // @[ivncontrol4.scala 254:54 257:22]
  wire [31:0] _GEN_615 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_609; // @[ivncontrol4.scala 254:54 258:22]
  wire [31:0] _GEN_616 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_610; // @[ivncontrol4.scala 254:54 259:22]
  wire [31:0] _GEN_617 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_611; // @[ivncontrol4.scala 254:54 260:22]
  wire [31:0] _GEN_618 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_478; // @[ivncontrol4.scala 245:49 246:22]
  wire [31:0] _GEN_619 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_612; // @[ivncontrol4.scala 245:49 247:21]
  wire [31:0] _GEN_620 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_613; // @[ivncontrol4.scala 245:49 248:21]
  wire [31:0] _GEN_621 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_614; // @[ivncontrol4.scala 245:49 249:22]
  wire [31:0] _GEN_622 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_615; // @[ivncontrol4.scala 245:49 250:22]
  wire [31:0] _GEN_623 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_616; // @[ivncontrol4.scala 245:49 251:22]
  wire [31:0] _GEN_624 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_617; // @[ivncontrol4.scala 245:49 252:22]
  wire [31:0] _GEN_642 = 4'h1 == _i_vn_1_T_15[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_643 = 4'h2 == _i_vn_1_T_15[3:0] ? rowcount_2 : _GEN_642; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_644 = 4'h3 == _i_vn_1_T_15[3:0] ? rowcount_3 : _GEN_643; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_645 = 4'h4 == _i_vn_1_T_15[3:0] ? rowcount_4 : _GEN_644; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_646 = 4'h5 == _i_vn_1_T_15[3:0] ? rowcount_5 : _GEN_645; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_647 = 4'h6 == _i_vn_1_T_15[3:0] ? rowcount_6 : _GEN_646; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_648 = 4'h7 == _i_vn_1_T_15[3:0] ? rowcount_7 : _GEN_647; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_649 = 4'h8 == _i_vn_1_T_15[3:0] ? rowcount_8 : _GEN_648; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_650 = 4'h9 == _i_vn_1_T_15[3:0] ? rowcount_9 : _GEN_649; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_651 = 4'ha == _i_vn_1_T_15[3:0] ? rowcount_10 : _GEN_650; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_652 = 4'hb == _i_vn_1_T_15[3:0] ? rowcount_11 : _GEN_651; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_653 = 4'hc == _i_vn_1_T_15[3:0] ? rowcount_12 : _GEN_652; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_654 = 4'hd == _i_vn_1_T_15[3:0] ? rowcount_13 : _GEN_653; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_655 = 4'he == _i_vn_1_T_15[3:0] ? rowcount_14 : _GEN_654; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_656 = 4'hf == _i_vn_1_T_15[3:0] ? rowcount_15 : _GEN_655; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _T_172 = _GEN_336 + _GEN_656; // @[ivncontrol4.scala 292:41]
  wire [31:0] _T_174 = 32'h8 - _T_172; // @[ivncontrol4.scala 292:18]
  wire [31:0] _i_vn_1_T_17 = 32'h2 + pin; // @[ivncontrol4.scala 293:29]
  wire [31:0] _GEN_849 = _T_174 == 32'h1 ? _i_vn_1_T_17 : _GEN_624; // @[ivncontrol4.scala 335:78 338:22]
  wire [31:0] _GEN_850 = _T_174 == 32'h2 ? _i_vn_1_T_17 : _GEN_623; // @[ivncontrol4.scala 329:76 332:22]
  wire [31:0] _GEN_851 = _T_174 == 32'h2 ? _i_vn_1_T_17 : _GEN_849; // @[ivncontrol4.scala 329:76 333:22]
  wire [31:0] _GEN_852 = _T_174 == 32'h3 ? _i_vn_1_T_17 : _GEN_622; // @[ivncontrol4.scala 322:78 324:23]
  wire [31:0] _GEN_853 = _T_174 == 32'h3 ? _i_vn_1_T_17 : _GEN_850; // @[ivncontrol4.scala 322:78 325:22]
  wire [31:0] _GEN_854 = _T_174 == 32'h3 ? _i_vn_1_T_17 : _GEN_851; // @[ivncontrol4.scala 322:78 326:22]
  wire [31:0] _GEN_855 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_621; // @[ivncontrol4.scala 316:78 318:22]
  wire [31:0] _GEN_856 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_852; // @[ivncontrol4.scala 316:78 319:22]
  wire [31:0] _GEN_857 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_853; // @[ivncontrol4.scala 316:78 320:22]
  wire [31:0] _GEN_858 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_854; // @[ivncontrol4.scala 316:78 321:22]
  wire [31:0] _GEN_859 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_620; // @[ivncontrol4.scala 309:76 311:23]
  wire [31:0] _GEN_860 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_855; // @[ivncontrol4.scala 309:76 312:22]
  wire [31:0] _GEN_861 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_856; // @[ivncontrol4.scala 309:76 313:22]
  wire [31:0] _GEN_862 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_857; // @[ivncontrol4.scala 309:76 314:22]
  wire [31:0] _GEN_863 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_858; // @[ivncontrol4.scala 309:76 315:22]
  wire [31:0] _GEN_864 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_619; // @[ivncontrol4.scala 301:77 303:22]
  wire [31:0] _GEN_865 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_859; // @[ivncontrol4.scala 301:77 304:21]
  wire [31:0] _GEN_866 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_860; // @[ivncontrol4.scala 301:77 305:22]
  wire [31:0] _GEN_867 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_861; // @[ivncontrol4.scala 301:77 306:22]
  wire [31:0] _GEN_868 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_862; // @[ivncontrol4.scala 301:77 307:22]
  wire [31:0] _GEN_869 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_863; // @[ivncontrol4.scala 301:77 308:22]
  wire [31:0] _GEN_870 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_618; // @[ivncontrol4.scala 292:73 293:22]
  wire [31:0] _GEN_871 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_864; // @[ivncontrol4.scala 292:73 294:21]
  wire [31:0] _GEN_872 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_865; // @[ivncontrol4.scala 292:73 295:21]
  wire [31:0] _GEN_873 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_866; // @[ivncontrol4.scala 292:73 296:22]
  wire [31:0] _GEN_874 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_867; // @[ivncontrol4.scala 292:73 297:22]
  wire [31:0] _GEN_875 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_868; // @[ivncontrol4.scala 292:73 298:22]
  wire [31:0] _GEN_876 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_869; // @[ivncontrol4.scala 292:73 299:22]
  wire [31:0] _GEN_910 = 4'h1 == _i_vn_1_T_17[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_911 = 4'h2 == _i_vn_1_T_17[3:0] ? rowcount_2 : _GEN_910; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_912 = 4'h3 == _i_vn_1_T_17[3:0] ? rowcount_3 : _GEN_911; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_913 = 4'h4 == _i_vn_1_T_17[3:0] ? rowcount_4 : _GEN_912; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_914 = 4'h5 == _i_vn_1_T_17[3:0] ? rowcount_5 : _GEN_913; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_915 = 4'h6 == _i_vn_1_T_17[3:0] ? rowcount_6 : _GEN_914; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_916 = 4'h7 == _i_vn_1_T_17[3:0] ? rowcount_7 : _GEN_915; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_917 = 4'h8 == _i_vn_1_T_17[3:0] ? rowcount_8 : _GEN_916; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_918 = 4'h9 == _i_vn_1_T_17[3:0] ? rowcount_9 : _GEN_917; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_919 = 4'ha == _i_vn_1_T_17[3:0] ? rowcount_10 : _GEN_918; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_920 = 4'hb == _i_vn_1_T_17[3:0] ? rowcount_11 : _GEN_919; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_921 = 4'hc == _i_vn_1_T_17[3:0] ? rowcount_12 : _GEN_920; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_922 = 4'hd == _i_vn_1_T_17[3:0] ? rowcount_13 : _GEN_921; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_923 = 4'he == _i_vn_1_T_17[3:0] ? rowcount_14 : _GEN_922; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_924 = 4'hf == _i_vn_1_T_17[3:0] ? rowcount_15 : _GEN_923; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _T_254 = _T_172 + _GEN_924; // @[ivncontrol4.scala 343:62]
  wire [31:0] _T_256 = 32'h8 - _T_254; // @[ivncontrol4.scala 343:17]
  wire [31:0] _i_vn_1_T_19 = 32'h3 + pin; // @[ivncontrol4.scala 344:29]
  wire [31:0] _GEN_1213 = _T_256 == 32'h1 ? _i_vn_1_T_19 : _GEN_876; // @[ivncontrol4.scala 386:100 389:22]
  wire [31:0] _GEN_1214 = _T_256 == 32'h2 ? _i_vn_1_T_19 : _GEN_875; // @[ivncontrol4.scala 380:98 383:22]
  wire [31:0] _GEN_1215 = _T_256 == 32'h2 ? _i_vn_1_T_19 : _GEN_1213; // @[ivncontrol4.scala 380:98 384:22]
  wire [31:0] _GEN_1216 = _T_256 == 32'h3 ? _i_vn_1_T_19 : _GEN_874; // @[ivncontrol4.scala 373:100 375:23]
  wire [31:0] _GEN_1217 = _T_256 == 32'h3 ? _i_vn_1_T_19 : _GEN_1214; // @[ivncontrol4.scala 373:100 376:22]
  wire [31:0] _GEN_1218 = _T_256 == 32'h3 ? _i_vn_1_T_19 : _GEN_1215; // @[ivncontrol4.scala 373:100 377:22]
  wire [31:0] _GEN_1219 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_873; // @[ivncontrol4.scala 367:100 369:22]
  wire [31:0] _GEN_1220 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_1216; // @[ivncontrol4.scala 367:100 370:22]
  wire [31:0] _GEN_1221 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_1217; // @[ivncontrol4.scala 367:100 371:22]
  wire [31:0] _GEN_1222 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_1218; // @[ivncontrol4.scala 367:100 372:22]
  wire [31:0] _GEN_1223 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_872; // @[ivncontrol4.scala 360:98 362:23]
  wire [31:0] _GEN_1224 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1219; // @[ivncontrol4.scala 360:98 363:22]
  wire [31:0] _GEN_1225 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1220; // @[ivncontrol4.scala 360:98 364:22]
  wire [31:0] _GEN_1226 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1221; // @[ivncontrol4.scala 360:98 365:22]
  wire [31:0] _GEN_1227 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1222; // @[ivncontrol4.scala 360:98 366:22]
  wire [31:0] _GEN_1228 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_871; // @[ivncontrol4.scala 352:99 354:22]
  wire [31:0] _GEN_1229 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1223; // @[ivncontrol4.scala 352:99 355:21]
  wire [31:0] _GEN_1230 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1224; // @[ivncontrol4.scala 352:99 356:22]
  wire [31:0] _GEN_1231 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1225; // @[ivncontrol4.scala 352:99 357:22]
  wire [31:0] _GEN_1232 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1226; // @[ivncontrol4.scala 352:99 358:22]
  wire [31:0] _GEN_1233 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1227; // @[ivncontrol4.scala 352:99 359:22]
  wire [31:0] _GEN_1234 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_870; // @[ivncontrol4.scala 343:94 344:22]
  wire [31:0] _GEN_1235 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1228; // @[ivncontrol4.scala 343:94 345:21]
  wire [31:0] _GEN_1236 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1229; // @[ivncontrol4.scala 343:94 346:21]
  wire [31:0] _GEN_1237 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1230; // @[ivncontrol4.scala 343:94 347:22]
  wire [31:0] _GEN_1238 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1231; // @[ivncontrol4.scala 343:94 348:22]
  wire [31:0] _GEN_1239 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1232; // @[ivncontrol4.scala 343:94 349:22]
  wire [31:0] _GEN_1240 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1233; // @[ivncontrol4.scala 343:94 350:22]
  wire [31:0] _GEN_1290 = 4'h1 == _i_vn_1_T_19[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1291 = 4'h2 == _i_vn_1_T_19[3:0] ? rowcount_2 : _GEN_1290; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1292 = 4'h3 == _i_vn_1_T_19[3:0] ? rowcount_3 : _GEN_1291; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1293 = 4'h4 == _i_vn_1_T_19[3:0] ? rowcount_4 : _GEN_1292; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1294 = 4'h5 == _i_vn_1_T_19[3:0] ? rowcount_5 : _GEN_1293; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1295 = 4'h6 == _i_vn_1_T_19[3:0] ? rowcount_6 : _GEN_1294; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1296 = 4'h7 == _i_vn_1_T_19[3:0] ? rowcount_7 : _GEN_1295; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1297 = 4'h8 == _i_vn_1_T_19[3:0] ? rowcount_8 : _GEN_1296; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1298 = 4'h9 == _i_vn_1_T_19[3:0] ? rowcount_9 : _GEN_1297; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1299 = 4'ha == _i_vn_1_T_19[3:0] ? rowcount_10 : _GEN_1298; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1300 = 4'hb == _i_vn_1_T_19[3:0] ? rowcount_11 : _GEN_1299; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1301 = 4'hc == _i_vn_1_T_19[3:0] ? rowcount_12 : _GEN_1300; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1302 = 4'hd == _i_vn_1_T_19[3:0] ? rowcount_13 : _GEN_1301; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1303 = 4'he == _i_vn_1_T_19[3:0] ? rowcount_14 : _GEN_1302; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1304 = 4'hf == _i_vn_1_T_19[3:0] ? rowcount_15 : _GEN_1303; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _T_371 = _T_254 + _GEN_1304; // @[ivncontrol4.scala 393:86]
  wire [31:0] _T_373 = 32'h8 - _T_371; // @[ivncontrol4.scala 393:19]
  wire [31:0] _i_vn_1_T_21 = 32'h4 + pin; // @[ivncontrol4.scala 394:29]
  wire [31:0] _GEN_1689 = _T_373 == 32'h1 ? _i_vn_1_T_21 : _GEN_1240; // @[ivncontrol4.scala 436:122 439:22]
  wire [31:0] _GEN_1690 = _T_373 == 32'h2 ? _i_vn_1_T_21 : _GEN_1239; // @[ivncontrol4.scala 430:121 433:22]
  wire [31:0] _GEN_1691 = _T_373 == 32'h2 ? _i_vn_1_T_21 : _GEN_1689; // @[ivncontrol4.scala 430:121 434:22]
  wire [31:0] _GEN_1692 = _T_373 == 32'h3 ? _i_vn_1_T_21 : _GEN_1238; // @[ivncontrol4.scala 423:123 425:23]
  wire [31:0] _GEN_1693 = _T_373 == 32'h3 ? _i_vn_1_T_21 : _GEN_1690; // @[ivncontrol4.scala 423:123 426:22]
  wire [31:0] _GEN_1694 = _T_373 == 32'h3 ? _i_vn_1_T_21 : _GEN_1691; // @[ivncontrol4.scala 423:123 427:22]
  wire [31:0] _GEN_1695 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1237; // @[ivncontrol4.scala 417:122 419:22]
  wire [31:0] _GEN_1696 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1692; // @[ivncontrol4.scala 417:122 420:22]
  wire [31:0] _GEN_1697 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1693; // @[ivncontrol4.scala 417:122 421:22]
  wire [31:0] _GEN_1698 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1694; // @[ivncontrol4.scala 417:122 422:22]
  wire [31:0] _GEN_1699 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1236; // @[ivncontrol4.scala 410:121 412:23]
  wire [31:0] _GEN_1700 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1695; // @[ivncontrol4.scala 410:121 413:22]
  wire [31:0] _GEN_1701 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1696; // @[ivncontrol4.scala 410:121 414:22]
  wire [31:0] _GEN_1702 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1697; // @[ivncontrol4.scala 410:121 415:22]
  wire [31:0] _GEN_1703 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1698; // @[ivncontrol4.scala 410:121 416:22]
  wire [31:0] _GEN_1704 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1235; // @[ivncontrol4.scala 402:121 404:22]
  wire [31:0] _GEN_1705 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1699; // @[ivncontrol4.scala 402:121 405:21]
  wire [31:0] _GEN_1706 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1700; // @[ivncontrol4.scala 402:121 406:22]
  wire [31:0] _GEN_1707 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1701; // @[ivncontrol4.scala 402:121 407:22]
  wire [31:0] _GEN_1708 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1702; // @[ivncontrol4.scala 402:121 408:22]
  wire [31:0] _GEN_1709 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1703; // @[ivncontrol4.scala 402:121 409:22]
  wire [31:0] _GEN_1710 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1234; // @[ivncontrol4.scala 393:118 394:22]
  wire [31:0] _GEN_1711 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1704; // @[ivncontrol4.scala 393:118 395:21]
  wire [31:0] _GEN_1712 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1705; // @[ivncontrol4.scala 393:118 396:21]
  wire [31:0] _GEN_1713 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1706; // @[ivncontrol4.scala 393:118 397:22]
  wire [31:0] _GEN_1714 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1707; // @[ivncontrol4.scala 393:118 398:22]
  wire [31:0] _GEN_1715 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1708; // @[ivncontrol4.scala 393:118 399:22]
  wire [31:0] _GEN_1716 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1709; // @[ivncontrol4.scala 393:118 400:22]
  wire [31:0] _GEN_1782 = 4'h1 == _i_vn_1_T_21[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1783 = 4'h2 == _i_vn_1_T_21[3:0] ? rowcount_2 : _GEN_1782; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1784 = 4'h3 == _i_vn_1_T_21[3:0] ? rowcount_3 : _GEN_1783; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1785 = 4'h4 == _i_vn_1_T_21[3:0] ? rowcount_4 : _GEN_1784; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1786 = 4'h5 == _i_vn_1_T_21[3:0] ? rowcount_5 : _GEN_1785; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1787 = 4'h6 == _i_vn_1_T_21[3:0] ? rowcount_6 : _GEN_1786; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1788 = 4'h7 == _i_vn_1_T_21[3:0] ? rowcount_7 : _GEN_1787; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1789 = 4'h8 == _i_vn_1_T_21[3:0] ? rowcount_8 : _GEN_1788; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1790 = 4'h9 == _i_vn_1_T_21[3:0] ? rowcount_9 : _GEN_1789; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1791 = 4'ha == _i_vn_1_T_21[3:0] ? rowcount_10 : _GEN_1790; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1792 = 4'hb == _i_vn_1_T_21[3:0] ? rowcount_11 : _GEN_1791; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1793 = 4'hc == _i_vn_1_T_21[3:0] ? rowcount_12 : _GEN_1792; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1794 = 4'hd == _i_vn_1_T_21[3:0] ? rowcount_13 : _GEN_1793; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1795 = 4'he == _i_vn_1_T_21[3:0] ? rowcount_14 : _GEN_1794; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1796 = 4'hf == _i_vn_1_T_21[3:0] ? rowcount_15 : _GEN_1795; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _T_523 = _T_371 + _GEN_1796; // @[ivncontrol4.scala 443:108]
  wire [31:0] _T_525 = 32'h8 - _T_523; // @[ivncontrol4.scala 443:19]
  wire [31:0] _i_vn_1_T_23 = 32'h5 + pin; // @[ivncontrol4.scala 444:29]
  wire [31:0] _GEN_2277 = _T_525 == 32'h1 ? _i_vn_1_T_23 : _GEN_1716; // @[ivncontrol4.scala 486:144 489:22]
  wire [31:0] _GEN_2278 = _T_525 == 32'h2 ? _i_vn_1_T_23 : _GEN_1715; // @[ivncontrol4.scala 480:143 483:22]
  wire [31:0] _GEN_2279 = _T_525 == 32'h2 ? _i_vn_1_T_23 : _GEN_2277; // @[ivncontrol4.scala 480:143 484:22]
  wire [31:0] _GEN_2280 = _T_525 == 32'h3 ? _i_vn_1_T_23 : _GEN_1714; // @[ivncontrol4.scala 473:145 475:23]
  wire [31:0] _GEN_2281 = _T_525 == 32'h3 ? _i_vn_1_T_23 : _GEN_2278; // @[ivncontrol4.scala 473:145 476:22]
  wire [31:0] _GEN_2282 = _T_525 == 32'h3 ? _i_vn_1_T_23 : _GEN_2279; // @[ivncontrol4.scala 473:145 477:22]
  wire [31:0] _GEN_2283 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_1713; // @[ivncontrol4.scala 467:143 469:22]
  wire [31:0] _GEN_2284 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_2280; // @[ivncontrol4.scala 467:143 470:22]
  wire [31:0] _GEN_2285 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_2281; // @[ivncontrol4.scala 467:143 471:22]
  wire [31:0] _GEN_2286 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_2282; // @[ivncontrol4.scala 467:143 472:22]
  wire [31:0] _GEN_2287 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_1712; // @[ivncontrol4.scala 460:143 462:23]
  wire [31:0] _GEN_2288 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2283; // @[ivncontrol4.scala 460:143 463:22]
  wire [31:0] _GEN_2289 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2284; // @[ivncontrol4.scala 460:143 464:22]
  wire [31:0] _GEN_2290 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2285; // @[ivncontrol4.scala 460:143 465:22]
  wire [31:0] _GEN_2291 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2286; // @[ivncontrol4.scala 460:143 466:22]
  wire [31:0] _GEN_2292 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_1711; // @[ivncontrol4.scala 452:143 454:22]
  wire [31:0] _GEN_2293 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2287; // @[ivncontrol4.scala 452:143 455:21]
  wire [31:0] _GEN_2294 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2288; // @[ivncontrol4.scala 452:143 456:22]
  wire [31:0] _GEN_2295 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2289; // @[ivncontrol4.scala 452:143 457:22]
  wire [31:0] _GEN_2296 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2290; // @[ivncontrol4.scala 452:143 458:22]
  wire [31:0] _GEN_2297 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2291; // @[ivncontrol4.scala 452:143 459:22]
  wire [31:0] _GEN_2298 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_1710; // @[ivncontrol4.scala 443:140 444:22]
  wire [31:0] _GEN_2299 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2292; // @[ivncontrol4.scala 443:140 445:21]
  wire [31:0] _GEN_2300 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2293; // @[ivncontrol4.scala 443:140 446:21]
  wire [31:0] _GEN_2301 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2294; // @[ivncontrol4.scala 443:140 447:22]
  wire [31:0] _GEN_2302 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2295; // @[ivncontrol4.scala 443:140 448:22]
  wire [31:0] _GEN_2303 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2296; // @[ivncontrol4.scala 443:140 449:22]
  wire [31:0] _GEN_2304 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2297; // @[ivncontrol4.scala 443:140 450:22]
  wire [31:0] _GEN_2386 = 4'h1 == _i_vn_1_T_23[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2387 = 4'h2 == _i_vn_1_T_23[3:0] ? rowcount_2 : _GEN_2386; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2388 = 4'h3 == _i_vn_1_T_23[3:0] ? rowcount_3 : _GEN_2387; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2389 = 4'h4 == _i_vn_1_T_23[3:0] ? rowcount_4 : _GEN_2388; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2390 = 4'h5 == _i_vn_1_T_23[3:0] ? rowcount_5 : _GEN_2389; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2391 = 4'h6 == _i_vn_1_T_23[3:0] ? rowcount_6 : _GEN_2390; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2392 = 4'h7 == _i_vn_1_T_23[3:0] ? rowcount_7 : _GEN_2391; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2393 = 4'h8 == _i_vn_1_T_23[3:0] ? rowcount_8 : _GEN_2392; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2394 = 4'h9 == _i_vn_1_T_23[3:0] ? rowcount_9 : _GEN_2393; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2395 = 4'ha == _i_vn_1_T_23[3:0] ? rowcount_10 : _GEN_2394; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2396 = 4'hb == _i_vn_1_T_23[3:0] ? rowcount_11 : _GEN_2395; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2397 = 4'hc == _i_vn_1_T_23[3:0] ? rowcount_12 : _GEN_2396; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2398 = 4'hd == _i_vn_1_T_23[3:0] ? rowcount_13 : _GEN_2397; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2399 = 4'he == _i_vn_1_T_23[3:0] ? rowcount_14 : _GEN_2398; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2400 = 4'hf == _i_vn_1_T_23[3:0] ? rowcount_15 : _GEN_2399; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _T_710 = _T_523 + _GEN_2400; // @[ivncontrol4.scala 494:130]
  wire [31:0] _T_712 = 32'h8 - _T_710; // @[ivncontrol4.scala 494:19]
  wire [31:0] _i_vn_1_T_25 = 32'h6 + pin; // @[ivncontrol4.scala 495:29]
  wire [31:0] _GEN_2977 = _T_712 == 32'h1 ? _i_vn_1_T_25 : _GEN_2304; // @[ivncontrol4.scala 537:166 540:22]
  wire [31:0] _GEN_2978 = _T_712 == 32'h2 ? _i_vn_1_T_25 : _GEN_2303; // @[ivncontrol4.scala 531:166 534:22]
  wire [31:0] _GEN_2979 = _T_712 == 32'h2 ? _i_vn_1_T_25 : _GEN_2977; // @[ivncontrol4.scala 531:166 535:22]
  wire [31:0] _GEN_2980 = _T_712 == 32'h3 ? _i_vn_1_T_25 : _GEN_2302; // @[ivncontrol4.scala 524:168 526:23]
  wire [31:0] _GEN_2981 = _T_712 == 32'h3 ? _i_vn_1_T_25 : _GEN_2978; // @[ivncontrol4.scala 524:168 527:22]
  wire [31:0] _GEN_2982 = _T_712 == 32'h3 ? _i_vn_1_T_25 : _GEN_2979; // @[ivncontrol4.scala 524:168 528:22]
  wire [31:0] _GEN_2983 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2301; // @[ivncontrol4.scala 518:166 520:22]
  wire [31:0] _GEN_2984 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2980; // @[ivncontrol4.scala 518:166 521:22]
  wire [31:0] _GEN_2985 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2981; // @[ivncontrol4.scala 518:166 522:22]
  wire [31:0] _GEN_2986 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2982; // @[ivncontrol4.scala 518:166 523:22]
  wire [31:0] _GEN_2987 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2300; // @[ivncontrol4.scala 511:166 513:23]
  wire [31:0] _GEN_2988 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2983; // @[ivncontrol4.scala 511:166 514:22]
  wire [31:0] _GEN_2989 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2984; // @[ivncontrol4.scala 511:166 515:22]
  wire [31:0] _GEN_2990 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2985; // @[ivncontrol4.scala 511:166 516:22]
  wire [31:0] _GEN_2991 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2986; // @[ivncontrol4.scala 511:166 517:22]
  wire [31:0] _GEN_2992 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2299; // @[ivncontrol4.scala 503:166 505:22]
  wire [31:0] _GEN_2993 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2987; // @[ivncontrol4.scala 503:166 506:21]
  wire [31:0] _GEN_2994 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2988; // @[ivncontrol4.scala 503:166 507:22]
  wire [31:0] _GEN_2995 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2989; // @[ivncontrol4.scala 503:166 508:22]
  wire [31:0] _GEN_2996 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2990; // @[ivncontrol4.scala 503:166 509:22]
  wire [31:0] _GEN_2997 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2991; // @[ivncontrol4.scala 503:166 510:22]
  wire [31:0] _GEN_2998 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2298; // @[ivncontrol4.scala 494:162 495:22]
  wire [31:0] _GEN_2999 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2992; // @[ivncontrol4.scala 494:162 496:21]
  wire [31:0] _GEN_3000 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2993; // @[ivncontrol4.scala 494:162 497:21]
  wire [31:0] _GEN_3001 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2994; // @[ivncontrol4.scala 494:162 498:22]
  wire [31:0] _GEN_3002 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2995; // @[ivncontrol4.scala 494:162 499:22]
  wire [31:0] _GEN_3003 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2996; // @[ivncontrol4.scala 494:162 500:22]
  wire [31:0] _GEN_3004 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2997; // @[ivncontrol4.scala 494:162 501:22]
  wire [31:0] _GEN_3102 = 4'h1 == _i_vn_1_T_25[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3103 = 4'h2 == _i_vn_1_T_25[3:0] ? rowcount_2 : _GEN_3102; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3104 = 4'h3 == _i_vn_1_T_25[3:0] ? rowcount_3 : _GEN_3103; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3105 = 4'h4 == _i_vn_1_T_25[3:0] ? rowcount_4 : _GEN_3104; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3106 = 4'h5 == _i_vn_1_T_25[3:0] ? rowcount_5 : _GEN_3105; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3107 = 4'h6 == _i_vn_1_T_25[3:0] ? rowcount_6 : _GEN_3106; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3108 = 4'h7 == _i_vn_1_T_25[3:0] ? rowcount_7 : _GEN_3107; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3109 = 4'h8 == _i_vn_1_T_25[3:0] ? rowcount_8 : _GEN_3108; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3110 = 4'h9 == _i_vn_1_T_25[3:0] ? rowcount_9 : _GEN_3109; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3111 = 4'ha == _i_vn_1_T_25[3:0] ? rowcount_10 : _GEN_3110; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3112 = 4'hb == _i_vn_1_T_25[3:0] ? rowcount_11 : _GEN_3111; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3113 = 4'hc == _i_vn_1_T_25[3:0] ? rowcount_12 : _GEN_3112; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3114 = 4'hd == _i_vn_1_T_25[3:0] ? rowcount_13 : _GEN_3113; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3115 = 4'he == _i_vn_1_T_25[3:0] ? rowcount_14 : _GEN_3114; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3116 = 4'hf == _i_vn_1_T_25[3:0] ? rowcount_15 : _GEN_3115; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _T_932 = _T_710 + _GEN_3116; // @[ivncontrol4.scala 545:152]
  wire [31:0] _T_934 = 32'h8 - _T_932; // @[ivncontrol4.scala 545:19]
  wire [31:0] _i_vn_1_T_27 = 32'h7 + pin; // @[ivncontrol4.scala 546:29]
  wire [31:0] _GEN_3789 = _T_934 == 32'h1 ? _i_vn_1_T_27 : _GEN_3004; // @[ivncontrol4.scala 588:188 591:22]
  wire [31:0] _GEN_3790 = _T_934 == 32'h2 ? _i_vn_1_T_27 : _GEN_3003; // @[ivncontrol4.scala 582:188 585:22]
  wire [31:0] _GEN_3791 = _T_934 == 32'h2 ? _i_vn_1_T_27 : _GEN_3789; // @[ivncontrol4.scala 582:188 586:22]
  wire [31:0] _GEN_3792 = _T_934 == 32'h3 ? _i_vn_1_T_27 : _GEN_3002; // @[ivncontrol4.scala 575:190 577:23]
  wire [31:0] _GEN_3793 = _T_934 == 32'h3 ? _i_vn_1_T_27 : _GEN_3790; // @[ivncontrol4.scala 575:190 578:22]
  wire [31:0] _GEN_3794 = _T_934 == 32'h3 ? _i_vn_1_T_27 : _GEN_3791; // @[ivncontrol4.scala 575:190 579:22]
  wire [31:0] _GEN_3795 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_3001; // @[ivncontrol4.scala 569:188 571:22]
  wire [31:0] _GEN_3796 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_3792; // @[ivncontrol4.scala 569:188 572:22]
  wire [31:0] _GEN_3797 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_3793; // @[ivncontrol4.scala 569:188 573:22]
  wire [31:0] _GEN_3798 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_3794; // @[ivncontrol4.scala 569:188 574:22]
  wire [31:0] _GEN_3799 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3000; // @[ivncontrol4.scala 562:188 564:23]
  wire [31:0] _GEN_3800 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3795; // @[ivncontrol4.scala 562:188 565:22]
  wire [31:0] _GEN_3801 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3796; // @[ivncontrol4.scala 562:188 566:22]
  wire [31:0] _GEN_3802 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3797; // @[ivncontrol4.scala 562:188 567:22]
  wire [31:0] _GEN_3803 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3798; // @[ivncontrol4.scala 562:188 568:22]
  wire [31:0] _GEN_3804 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_2999; // @[ivncontrol4.scala 554:188 556:22]
  wire [31:0] _GEN_3805 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3799; // @[ivncontrol4.scala 554:188 557:21]
  wire [31:0] _GEN_3806 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3800; // @[ivncontrol4.scala 554:188 558:22]
  wire [31:0] _GEN_3807 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3801; // @[ivncontrol4.scala 554:188 559:22]
  wire [31:0] _GEN_3808 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3802; // @[ivncontrol4.scala 554:188 560:22]
  wire [31:0] _GEN_3809 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3803; // @[ivncontrol4.scala 554:188 561:22]
  wire [31:0] _GEN_3810 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_2998; // @[ivncontrol4.scala 545:184 546:22]
  wire [31:0] _GEN_3811 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3804; // @[ivncontrol4.scala 545:184 547:21]
  wire [31:0] _GEN_3812 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3805; // @[ivncontrol4.scala 545:184 548:21]
  wire [31:0] _GEN_3813 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3806; // @[ivncontrol4.scala 545:184 549:22]
  wire [31:0] _GEN_3814 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3807; // @[ivncontrol4.scala 545:184 550:22]
  wire [31:0] _GEN_3815 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3808; // @[ivncontrol4.scala 545:184 551:22]
  wire [31:0] _GEN_3816 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3809; // @[ivncontrol4.scala 545:184 552:22]
  wire [31:0] _GEN_3817 = _GEN_312 ? _GEN_477 : 32'h10; // @[ivncontrol4.scala 142:17 189:28]
  wire [31:0] _GEN_3818 = _GEN_312 ? _GEN_3810 : 32'h8; // @[ivncontrol4.scala 142:17 189:28]
  wire [31:0] _GEN_3819 = _GEN_312 ? _GEN_3811 : 32'ha; // @[ivncontrol4.scala 142:17 189:28]
  wire [31:0] _GEN_3820 = _GEN_312 ? _GEN_3812 : 32'h5; // @[ivncontrol4.scala 142:17 189:28]
  wire [31:0] _GEN_3821 = _GEN_312 ? _GEN_3813 : 32'h17; // @[ivncontrol4.scala 143:18 189:28]
  wire [31:0] _GEN_3822 = _GEN_312 ? _GEN_3814 : 32'h14; // @[ivncontrol4.scala 143:18 189:28]
  wire [31:0] _GEN_3823 = _GEN_312 ? _GEN_3815 : 32'h1; // @[ivncontrol4.scala 143:18 189:28]
  wire [31:0] _GEN_3824 = _GEN_312 ? _GEN_3816 : 32'hc; // @[ivncontrol4.scala 143:18 189:28]
  wire  valid1 = 1'h0;
  wire [31:0] _GEN_4221 = reset ? 32'h0 : _GEN_3817; // @[ivncontrol4.scala 17:{23,23}]
  wire [31:0] _GEN_4222 = reset ? 32'h0 : _GEN_3818; // @[ivncontrol4.scala 17:{23,23}]
  wire [31:0] _GEN_4223 = reset ? 32'h0 : _GEN_3819; // @[ivncontrol4.scala 17:{23,23}]
  wire [31:0] _GEN_4224 = reset ? 32'h0 : _GEN_3820; // @[ivncontrol4.scala 17:{23,23}]
  wire [31:0] _GEN_4225 = reset ? 32'h0 : _GEN_3821; // @[ivncontrol4.scala 18:{24,24}]
  wire [31:0] _GEN_4226 = reset ? 32'h0 : _GEN_3822; // @[ivncontrol4.scala 18:{24,24}]
  wire [31:0] _GEN_4227 = reset ? 32'h0 : _GEN_3823; // @[ivncontrol4.scala 18:{24,24}]
  wire [31:0] _GEN_4228 = reset ? 32'h0 : _GEN_3824; // @[ivncontrol4.scala 18:{24,24}]
  assign io_o_vn_0 = i_vn_0; // @[ivncontrol4.scala 138:13]
  assign io_o_vn_1 = i_vn_1; // @[ivncontrol4.scala 138:13]
  assign io_o_vn_2 = i_vn_2; // @[ivncontrol4.scala 138:13]
  assign io_o_vn_3 = i_vn_3; // @[ivncontrol4.scala 138:13]
  assign io_o_vn2_0 = i_vn2_0; // @[ivncontrol4.scala 139:14]
  assign io_o_vn2_1 = i_vn2_1; // @[ivncontrol4.scala 139:14]
  assign io_o_vn2_2 = i_vn2_2; // @[ivncontrol4.scala 139:14]
  assign io_o_vn2_3 = i_vn2_3; // @[ivncontrol4.scala 139:14]
  always @(posedge clock) begin
    i_vn_0 <= _GEN_4221[4:0]; // @[ivncontrol4.scala 17:{23,23}]
    i_vn_1 <= _GEN_4222[4:0]; // @[ivncontrol4.scala 17:{23,23}]
    i_vn_2 <= _GEN_4223[4:0]; // @[ivncontrol4.scala 17:{23,23}]
    i_vn_3 <= _GEN_4224[4:0]; // @[ivncontrol4.scala 17:{23,23}]
    i_vn2_0 <= _GEN_4225[4:0]; // @[ivncontrol4.scala 18:{24,24}]
    i_vn2_1 <= _GEN_4226[4:0]; // @[ivncontrol4.scala 18:{24,24}]
    i_vn2_2 <= _GEN_4227[4:0]; // @[ivncontrol4.scala 18:{24,24}]
    i_vn2_3 <= _GEN_4228[4:0]; // @[ivncontrol4.scala 18:{24,24}]
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_0 <= io_Stationary_matrix_0_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_1 <= io_Stationary_matrix_0_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_2 <= io_Stationary_matrix_0_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_3 <= io_Stationary_matrix_0_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_4 <= io_Stationary_matrix_0_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_5 <= io_Stationary_matrix_0_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_6 <= io_Stationary_matrix_0_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_7 <= io_Stationary_matrix_0_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_0 <= io_Stationary_matrix_1_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_1 <= io_Stationary_matrix_1_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_2 <= io_Stationary_matrix_1_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_3 <= io_Stationary_matrix_1_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_4 <= io_Stationary_matrix_1_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_5 <= io_Stationary_matrix_1_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_6 <= io_Stationary_matrix_1_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_7 <= io_Stationary_matrix_1_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_0 <= io_Stationary_matrix_2_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_1 <= io_Stationary_matrix_2_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_2 <= io_Stationary_matrix_2_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_3 <= io_Stationary_matrix_2_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_4 <= io_Stationary_matrix_2_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_5 <= io_Stationary_matrix_2_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_6 <= io_Stationary_matrix_2_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_7 <= io_Stationary_matrix_2_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_0 <= io_Stationary_matrix_3_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_1 <= io_Stationary_matrix_3_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_2 <= io_Stationary_matrix_3_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_3 <= io_Stationary_matrix_3_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_4 <= io_Stationary_matrix_3_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_5 <= io_Stationary_matrix_3_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_6 <= io_Stationary_matrix_3_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_7 <= io_Stationary_matrix_3_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_0 <= io_Stationary_matrix_4_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_1 <= io_Stationary_matrix_4_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_2 <= io_Stationary_matrix_4_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_3 <= io_Stationary_matrix_4_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_4 <= io_Stationary_matrix_4_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_5 <= io_Stationary_matrix_4_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_6 <= io_Stationary_matrix_4_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_7 <= io_Stationary_matrix_4_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_0 <= io_Stationary_matrix_5_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_1 <= io_Stationary_matrix_5_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_2 <= io_Stationary_matrix_5_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_3 <= io_Stationary_matrix_5_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_4 <= io_Stationary_matrix_5_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_5 <= io_Stationary_matrix_5_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_6 <= io_Stationary_matrix_5_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_7 <= io_Stationary_matrix_5_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_0 <= io_Stationary_matrix_6_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_1 <= io_Stationary_matrix_6_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_2 <= io_Stationary_matrix_6_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_3 <= io_Stationary_matrix_6_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_4 <= io_Stationary_matrix_6_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_5 <= io_Stationary_matrix_6_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_6 <= io_Stationary_matrix_6_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_7 <= io_Stationary_matrix_6_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_0 <= io_Stationary_matrix_7_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_1 <= io_Stationary_matrix_7_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_2 <= io_Stationary_matrix_7_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_3 <= io_Stationary_matrix_7_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_4 <= io_Stationary_matrix_7_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_5 <= io_Stationary_matrix_7_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_6 <= io_Stationary_matrix_7_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_7 <= io_Stationary_matrix_7_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_0 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_0 <= count_0; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_1 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_1 <= count_1; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_2 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_2 <= count_2; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_3 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_3 <= count_3; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_4 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_4 <= count_4; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_5 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_5 <= count_5; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_6 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_6 <= count_6; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_7 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_7 <= count_7; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_8 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_8 <= 32'h0; // @[ivncontrol4.scala 87:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_9 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_9 <= 32'h0; // @[ivncontrol4.scala 87:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_10 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_10 <= 32'h0; // @[ivncontrol4.scala 87:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_11 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_11 <= 32'h0; // @[ivncontrol4.scala 87:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_12 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_12 <= 32'h0; // @[ivncontrol4.scala 87:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_13 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_13 <= 32'h0; // @[ivncontrol4.scala 87:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_14 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_14 <= 32'h0; // @[ivncontrol4.scala 87:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_15 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end
    if (reset) begin // @[ivncontrol4.scala 37:22]
      pin <= 32'h0; // @[ivncontrol4.scala 37:22]
    end else if (_T_72 & rowcount_6 == 32'h0 & rowcount_7 != 32'h0) begin // @[ivncontrol4.scala 183:192]
      pin <= 32'h7; // @[ivncontrol4.scala 184:13]
    end else if (_T_59 & rowcount_5 == 32'h0 & rowcount_6 != 32'h0) begin // @[ivncontrol4.scala 180:169]
      pin <= 32'h6; // @[ivncontrol4.scala 181:13]
    end else if (_T_48 & rowcount_4 == 32'h0 & rowcount_5 != 32'h0) begin // @[ivncontrol4.scala 177:146]
      pin <= 32'h5; // @[ivncontrol4.scala 178:13]
    end else begin
      pin <= _GEN_317;
    end
    if (reset) begin // @[ivncontrol4.scala 41:20]
      i <= 32'h0; // @[ivncontrol4.scala 41:20]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
        i <= _GEN_247;
      end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
        i <= _GEN_247;
      end else begin
        i <= _GEN_265;
      end
    end
    if (reset) begin // @[ivncontrol4.scala 42:20]
      j <= 32'h0; // @[ivncontrol4.scala 42:20]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
        j <= 32'h8; // @[ivncontrol4.scala 116:11]
      end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
        j <= _j_T_1; // @[ivncontrol4.scala 118:11]
      end else begin
        j <= {{28'd0}, _GEN_264};
      end
    end
    if (3'h0 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h0 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h0 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h0 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h0 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h0 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h0 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h0 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_0 <= _GEN_224;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_0 <= _GEN_224;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h0 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_0 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_0 <= _GEN_224;
      end
    end else begin
      count_0 <= _GEN_224;
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_1 <= _GEN_225;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_1 <= _GEN_225;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h1 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_1 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_1 <= _GEN_225;
      end
    end else begin
      count_1 <= _GEN_225;
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_2 <= _GEN_226;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_2 <= _GEN_226;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h2 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_2 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_2 <= _GEN_226;
      end
    end else begin
      count_2 <= _GEN_226;
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_3 <= _GEN_227;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_3 <= _GEN_227;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h3 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_3 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_3 <= _GEN_227;
      end
    end else begin
      count_3 <= _GEN_227;
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_4 <= _GEN_228;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_4 <= _GEN_228;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h4 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_4 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_4 <= _GEN_228;
      end
    end else begin
      count_4 <= _GEN_228;
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_5 <= _GEN_229;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_5 <= _GEN_229;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h5 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_5 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_5 <= _GEN_229;
      end
    end else begin
      count_5 <= _GEN_229;
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_6 <= _GEN_230;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_6 <= _GEN_230;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h6 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_6 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_6 <= _GEN_230;
      end
    end else begin
      count_6 <= _GEN_230;
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_7 <= _GEN_231;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_7 <= _GEN_231;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h7 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_7 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_7 <= _GEN_231;
      end
    end else begin
      count_7 <= _GEN_231;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  i_vn_0 = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  i_vn_1 = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  i_vn_2 = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  i_vn_3 = _RAND_3[4:0];
  _RAND_4 = {1{`RANDOM}};
  i_vn2_0 = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  i_vn2_1 = _RAND_5[4:0];
  _RAND_6 = {1{`RANDOM}};
  i_vn2_2 = _RAND_6[4:0];
  _RAND_7 = {1{`RANDOM}};
  i_vn2_3 = _RAND_7[4:0];
  _RAND_8 = {1{`RANDOM}};
  solution_0_0 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  solution_0_1 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  solution_0_2 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  solution_0_3 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  solution_0_4 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  solution_0_5 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  solution_0_6 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  solution_0_7 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  solution_1_0 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  solution_1_1 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  solution_1_2 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  solution_1_3 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  solution_1_4 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  solution_1_5 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  solution_1_6 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  solution_1_7 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  solution_2_0 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  solution_2_1 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  solution_2_2 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  solution_2_3 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  solution_2_4 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  solution_2_5 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  solution_2_6 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  solution_2_7 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  solution_3_0 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  solution_3_1 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  solution_3_2 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  solution_3_3 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  solution_3_4 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  solution_3_5 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  solution_3_6 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  solution_3_7 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  solution_4_0 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  solution_4_1 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  solution_4_2 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  solution_4_3 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  solution_4_4 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  solution_4_5 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  solution_4_6 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  solution_4_7 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  solution_5_0 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  solution_5_1 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  solution_5_2 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  solution_5_3 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  solution_5_4 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  solution_5_5 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  solution_5_6 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  solution_5_7 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  solution_6_0 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  solution_6_1 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  solution_6_2 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  solution_6_3 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  solution_6_4 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  solution_6_5 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  solution_6_6 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  solution_6_7 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  solution_7_0 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  solution_7_1 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  solution_7_2 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  solution_7_3 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  solution_7_4 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  solution_7_5 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  solution_7_6 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  solution_7_7 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  rowcount_0 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  rowcount_1 = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  rowcount_2 = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  rowcount_3 = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  rowcount_4 = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  rowcount_5 = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  rowcount_6 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  rowcount_7 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  rowcount_8 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  rowcount_9 = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  rowcount_10 = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  rowcount_11 = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  rowcount_12 = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  rowcount_13 = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  rowcount_14 = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  rowcount_15 = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  pin = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  i = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  j = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  mat_0_0 = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  mat_0_1 = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  mat_0_2 = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  mat_0_3 = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  mat_0_4 = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  mat_0_5 = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  mat_0_6 = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  mat_0_7 = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  mat_1_0 = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  mat_1_1 = _RAND_100[31:0];
  _RAND_101 = {1{`RANDOM}};
  mat_1_2 = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  mat_1_3 = _RAND_102[31:0];
  _RAND_103 = {1{`RANDOM}};
  mat_1_4 = _RAND_103[31:0];
  _RAND_104 = {1{`RANDOM}};
  mat_1_5 = _RAND_104[31:0];
  _RAND_105 = {1{`RANDOM}};
  mat_1_6 = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  mat_1_7 = _RAND_106[31:0];
  _RAND_107 = {1{`RANDOM}};
  mat_2_0 = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  mat_2_1 = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  mat_2_2 = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  mat_2_3 = _RAND_110[31:0];
  _RAND_111 = {1{`RANDOM}};
  mat_2_4 = _RAND_111[31:0];
  _RAND_112 = {1{`RANDOM}};
  mat_2_5 = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  mat_2_6 = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  mat_2_7 = _RAND_114[31:0];
  _RAND_115 = {1{`RANDOM}};
  mat_3_0 = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  mat_3_1 = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  mat_3_2 = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  mat_3_3 = _RAND_118[31:0];
  _RAND_119 = {1{`RANDOM}};
  mat_3_4 = _RAND_119[31:0];
  _RAND_120 = {1{`RANDOM}};
  mat_3_5 = _RAND_120[31:0];
  _RAND_121 = {1{`RANDOM}};
  mat_3_6 = _RAND_121[31:0];
  _RAND_122 = {1{`RANDOM}};
  mat_3_7 = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  mat_4_0 = _RAND_123[31:0];
  _RAND_124 = {1{`RANDOM}};
  mat_4_1 = _RAND_124[31:0];
  _RAND_125 = {1{`RANDOM}};
  mat_4_2 = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  mat_4_3 = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  mat_4_4 = _RAND_127[31:0];
  _RAND_128 = {1{`RANDOM}};
  mat_4_5 = _RAND_128[31:0];
  _RAND_129 = {1{`RANDOM}};
  mat_4_6 = _RAND_129[31:0];
  _RAND_130 = {1{`RANDOM}};
  mat_4_7 = _RAND_130[31:0];
  _RAND_131 = {1{`RANDOM}};
  mat_5_0 = _RAND_131[31:0];
  _RAND_132 = {1{`RANDOM}};
  mat_5_1 = _RAND_132[31:0];
  _RAND_133 = {1{`RANDOM}};
  mat_5_2 = _RAND_133[31:0];
  _RAND_134 = {1{`RANDOM}};
  mat_5_3 = _RAND_134[31:0];
  _RAND_135 = {1{`RANDOM}};
  mat_5_4 = _RAND_135[31:0];
  _RAND_136 = {1{`RANDOM}};
  mat_5_5 = _RAND_136[31:0];
  _RAND_137 = {1{`RANDOM}};
  mat_5_6 = _RAND_137[31:0];
  _RAND_138 = {1{`RANDOM}};
  mat_5_7 = _RAND_138[31:0];
  _RAND_139 = {1{`RANDOM}};
  mat_6_0 = _RAND_139[31:0];
  _RAND_140 = {1{`RANDOM}};
  mat_6_1 = _RAND_140[31:0];
  _RAND_141 = {1{`RANDOM}};
  mat_6_2 = _RAND_141[31:0];
  _RAND_142 = {1{`RANDOM}};
  mat_6_3 = _RAND_142[31:0];
  _RAND_143 = {1{`RANDOM}};
  mat_6_4 = _RAND_143[31:0];
  _RAND_144 = {1{`RANDOM}};
  mat_6_5 = _RAND_144[31:0];
  _RAND_145 = {1{`RANDOM}};
  mat_6_6 = _RAND_145[31:0];
  _RAND_146 = {1{`RANDOM}};
  mat_6_7 = _RAND_146[31:0];
  _RAND_147 = {1{`RANDOM}};
  mat_7_0 = _RAND_147[31:0];
  _RAND_148 = {1{`RANDOM}};
  mat_7_1 = _RAND_148[31:0];
  _RAND_149 = {1{`RANDOM}};
  mat_7_2 = _RAND_149[31:0];
  _RAND_150 = {1{`RANDOM}};
  mat_7_3 = _RAND_150[31:0];
  _RAND_151 = {1{`RANDOM}};
  mat_7_4 = _RAND_151[31:0];
  _RAND_152 = {1{`RANDOM}};
  mat_7_5 = _RAND_152[31:0];
  _RAND_153 = {1{`RANDOM}};
  mat_7_6 = _RAND_153[31:0];
  _RAND_154 = {1{`RANDOM}};
  mat_7_7 = _RAND_154[31:0];
  _RAND_155 = {1{`RANDOM}};
  count_0 = _RAND_155[31:0];
  _RAND_156 = {1{`RANDOM}};
  count_1 = _RAND_156[31:0];
  _RAND_157 = {1{`RANDOM}};
  count_2 = _RAND_157[31:0];
  _RAND_158 = {1{`RANDOM}};
  count_3 = _RAND_158[31:0];
  _RAND_159 = {1{`RANDOM}};
  count_4 = _RAND_159[31:0];
  _RAND_160 = {1{`RANDOM}};
  count_5 = _RAND_160[31:0];
  _RAND_161 = {1{`RANDOM}};
  count_6 = _RAND_161[31:0];
  _RAND_162 = {1{`RANDOM}};
  count_7 = _RAND_162[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ivncontrol4_2(
  input         clock,
  input         reset,
  input  [15:0] io_Stationary_matrix_0_0,
  input  [15:0] io_Stationary_matrix_0_1,
  input  [15:0] io_Stationary_matrix_0_2,
  input  [15:0] io_Stationary_matrix_0_3,
  input  [15:0] io_Stationary_matrix_0_4,
  input  [15:0] io_Stationary_matrix_0_5,
  input  [15:0] io_Stationary_matrix_0_6,
  input  [15:0] io_Stationary_matrix_0_7,
  input  [15:0] io_Stationary_matrix_1_0,
  input  [15:0] io_Stationary_matrix_1_1,
  input  [15:0] io_Stationary_matrix_1_2,
  input  [15:0] io_Stationary_matrix_1_3,
  input  [15:0] io_Stationary_matrix_1_4,
  input  [15:0] io_Stationary_matrix_1_5,
  input  [15:0] io_Stationary_matrix_1_6,
  input  [15:0] io_Stationary_matrix_1_7,
  input  [15:0] io_Stationary_matrix_2_0,
  input  [15:0] io_Stationary_matrix_2_1,
  input  [15:0] io_Stationary_matrix_2_2,
  input  [15:0] io_Stationary_matrix_2_3,
  input  [15:0] io_Stationary_matrix_2_4,
  input  [15:0] io_Stationary_matrix_2_5,
  input  [15:0] io_Stationary_matrix_2_6,
  input  [15:0] io_Stationary_matrix_2_7,
  input  [15:0] io_Stationary_matrix_3_0,
  input  [15:0] io_Stationary_matrix_3_1,
  input  [15:0] io_Stationary_matrix_3_2,
  input  [15:0] io_Stationary_matrix_3_3,
  input  [15:0] io_Stationary_matrix_3_4,
  input  [15:0] io_Stationary_matrix_3_5,
  input  [15:0] io_Stationary_matrix_3_6,
  input  [15:0] io_Stationary_matrix_3_7,
  input  [15:0] io_Stationary_matrix_4_0,
  input  [15:0] io_Stationary_matrix_4_1,
  input  [15:0] io_Stationary_matrix_4_2,
  input  [15:0] io_Stationary_matrix_4_3,
  input  [15:0] io_Stationary_matrix_4_4,
  input  [15:0] io_Stationary_matrix_4_5,
  input  [15:0] io_Stationary_matrix_4_6,
  input  [15:0] io_Stationary_matrix_4_7,
  input  [15:0] io_Stationary_matrix_5_0,
  input  [15:0] io_Stationary_matrix_5_1,
  input  [15:0] io_Stationary_matrix_5_2,
  input  [15:0] io_Stationary_matrix_5_3,
  input  [15:0] io_Stationary_matrix_5_4,
  input  [15:0] io_Stationary_matrix_5_5,
  input  [15:0] io_Stationary_matrix_5_6,
  input  [15:0] io_Stationary_matrix_5_7,
  input  [15:0] io_Stationary_matrix_6_0,
  input  [15:0] io_Stationary_matrix_6_1,
  input  [15:0] io_Stationary_matrix_6_2,
  input  [15:0] io_Stationary_matrix_6_3,
  input  [15:0] io_Stationary_matrix_6_4,
  input  [15:0] io_Stationary_matrix_6_5,
  input  [15:0] io_Stationary_matrix_6_6,
  input  [15:0] io_Stationary_matrix_6_7,
  input  [15:0] io_Stationary_matrix_7_0,
  input  [15:0] io_Stationary_matrix_7_1,
  input  [15:0] io_Stationary_matrix_7_2,
  input  [15:0] io_Stationary_matrix_7_3,
  input  [15:0] io_Stationary_matrix_7_4,
  input  [15:0] io_Stationary_matrix_7_5,
  input  [15:0] io_Stationary_matrix_7_6,
  input  [15:0] io_Stationary_matrix_7_7,
  output [4:0]  io_o_vn_0,
  output [4:0]  io_o_vn_1,
  output [4:0]  io_o_vn_2,
  output [4:0]  io_o_vn_3,
  output [4:0]  io_o_vn2_0,
  output [4:0]  io_o_vn2_1,
  output [4:0]  io_o_vn2_2,
  output [4:0]  io_o_vn2_3,
  input         io_validpin
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
`endif // RANDOMIZE_REG_INIT
  reg [4:0] i_vn_0; // @[ivncontrol4.scala 17:23]
  reg [4:0] i_vn_1; // @[ivncontrol4.scala 17:23]
  reg [4:0] i_vn_2; // @[ivncontrol4.scala 17:23]
  reg [4:0] i_vn_3; // @[ivncontrol4.scala 17:23]
  reg [4:0] i_vn2_0; // @[ivncontrol4.scala 18:24]
  reg [4:0] i_vn2_1; // @[ivncontrol4.scala 18:24]
  reg [4:0] i_vn2_2; // @[ivncontrol4.scala 18:24]
  reg [4:0] i_vn2_3; // @[ivncontrol4.scala 18:24]
  reg [15:0] solution_0_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_0_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_0_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_0_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_0_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_0_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_0_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_0_7; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_7; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_7; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_7; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_7; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_7; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_7; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_7; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_0; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_1; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_2; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_3; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_4; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_5; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_6; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_7; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_8; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_9; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_10; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_11; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_12; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_13; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_14; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_15; // @[ivncontrol4.scala 27:27]
  reg [31:0] pin; // @[ivncontrol4.scala 37:22]
  reg [31:0] i; // @[ivncontrol4.scala 41:20]
  reg [31:0] j; // @[ivncontrol4.scala 42:20]
  wire  _io_ProcessValid_T = i == 32'h7; // @[ivncontrol4.scala 44:27]
  wire  _io_ProcessValid_T_1 = j == 32'h7; // @[ivncontrol4.scala 44:42]
  wire  _io_ProcessValid_T_2 = i == 32'h7 & j == 32'h7; // @[ivncontrol4.scala 44:36]
  reg [31:0] mat_0_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_0_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_0_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_0_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_0_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_0_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_0_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_0_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] count_0; // @[ivncontrol4.scala 58:20]
  reg [31:0] count_1; // @[ivncontrol4.scala 58:20]
  reg [31:0] count_2; // @[ivncontrol4.scala 58:20]
  reg [31:0] count_3; // @[ivncontrol4.scala 58:20]
  reg [31:0] count_4; // @[ivncontrol4.scala 58:20]
  reg [31:0] count_5; // @[ivncontrol4.scala 58:20]
  reg [31:0] count_6; // @[ivncontrol4.scala 58:20]
  reg [31:0] count_7; // @[ivncontrol4.scala 58:20]
  wire  _GEN_3825 = 3'h0 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_65 = 3'h0 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_0_1 : io_Stationary_matrix_0_0; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_66 = 3'h0 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_0_2 : _GEN_65; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_67 = 3'h0 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_0_3 : _GEN_66; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_68 = 3'h0 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_0_4 : _GEN_67; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_69 = 3'h0 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_0_5 : _GEN_68; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_70 = 3'h0 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_0_6 : _GEN_69; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_71 = 3'h0 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_0_7 : _GEN_70; // @[ivncontrol4.scala 63:{17,17}]
  wire  _GEN_3839 = 3'h1 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_72 = 3'h1 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_1_0 : _GEN_71; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_73 = 3'h1 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_1_1 : _GEN_72; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_74 = 3'h1 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_1_2 : _GEN_73; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_75 = 3'h1 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_1_3 : _GEN_74; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_76 = 3'h1 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_1_4 : _GEN_75; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_77 = 3'h1 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_1_5 : _GEN_76; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_78 = 3'h1 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_1_6 : _GEN_77; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_79 = 3'h1 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_1_7 : _GEN_78; // @[ivncontrol4.scala 63:{17,17}]
  wire  _GEN_3855 = 3'h2 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_80 = 3'h2 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_2_0 : _GEN_79; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_81 = 3'h2 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_2_1 : _GEN_80; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_82 = 3'h2 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_2_2 : _GEN_81; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_83 = 3'h2 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_2_3 : _GEN_82; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_84 = 3'h2 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_2_4 : _GEN_83; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_85 = 3'h2 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_2_5 : _GEN_84; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_86 = 3'h2 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_2_6 : _GEN_85; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_87 = 3'h2 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_2_7 : _GEN_86; // @[ivncontrol4.scala 63:{17,17}]
  wire  _GEN_3871 = 3'h3 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_88 = 3'h3 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_3_0 : _GEN_87; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_89 = 3'h3 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_3_1 : _GEN_88; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_90 = 3'h3 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_3_2 : _GEN_89; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_91 = 3'h3 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_3_3 : _GEN_90; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_92 = 3'h3 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_3_4 : _GEN_91; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_93 = 3'h3 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_3_5 : _GEN_92; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_94 = 3'h3 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_3_6 : _GEN_93; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_95 = 3'h3 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_3_7 : _GEN_94; // @[ivncontrol4.scala 63:{17,17}]
  wire  _GEN_3887 = 3'h4 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_96 = 3'h4 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_4_0 : _GEN_95; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_97 = 3'h4 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_4_1 : _GEN_96; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_98 = 3'h4 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_4_2 : _GEN_97; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_99 = 3'h4 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_4_3 : _GEN_98; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_100 = 3'h4 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_4_4 : _GEN_99; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_101 = 3'h4 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_4_5 : _GEN_100; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_102 = 3'h4 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_4_6 : _GEN_101; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_103 = 3'h4 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_4_7 : _GEN_102; // @[ivncontrol4.scala 63:{17,17}]
  wire  _GEN_3903 = 3'h5 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_104 = 3'h5 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_5_0 : _GEN_103; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_105 = 3'h5 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_5_1 : _GEN_104; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_106 = 3'h5 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_5_2 : _GEN_105; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_107 = 3'h5 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_5_3 : _GEN_106; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_108 = 3'h5 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_5_4 : _GEN_107; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_109 = 3'h5 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_5_5 : _GEN_108; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_110 = 3'h5 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_5_6 : _GEN_109; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_111 = 3'h5 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_5_7 : _GEN_110; // @[ivncontrol4.scala 63:{17,17}]
  wire  _GEN_3919 = 3'h6 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_112 = 3'h6 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_6_0 : _GEN_111; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_113 = 3'h6 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_6_1 : _GEN_112; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_114 = 3'h6 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_6_2 : _GEN_113; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_115 = 3'h6 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_6_3 : _GEN_114; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_116 = 3'h6 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_6_4 : _GEN_115; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_117 = 3'h6 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_6_5 : _GEN_116; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_118 = 3'h6 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_6_6 : _GEN_117; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_119 = 3'h6 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_6_7 : _GEN_118; // @[ivncontrol4.scala 63:{17,17}]
  wire  _GEN_3935 = 3'h7 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_120 = 3'h7 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_7_0 : _GEN_119; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_121 = 3'h7 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_7_1 : _GEN_120; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_122 = 3'h7 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_7_2 : _GEN_121; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_123 = 3'h7 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_7_3 : _GEN_122; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_124 = 3'h7 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_7_4 : _GEN_123; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_125 = 3'h7 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_7_5 : _GEN_124; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_126 = 3'h7 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_7_6 : _GEN_125; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_127 = 3'h7 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_7_7 : _GEN_126; // @[ivncontrol4.scala 63:{17,17}]
  wire [31:0] _mat_T_1_T_2 = {{16'd0}, _GEN_127}; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_129 = _GEN_3825 & 4'h1 == j[3:0] ? solution_0_1 : solution_0_0; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_130 = _GEN_3825 & 4'h2 == j[3:0] ? solution_0_2 : _GEN_129; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_131 = _GEN_3825 & 4'h3 == j[3:0] ? solution_0_3 : _GEN_130; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_132 = _GEN_3825 & 4'h4 == j[3:0] ? solution_0_4 : _GEN_131; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_133 = _GEN_3825 & 4'h5 == j[3:0] ? solution_0_5 : _GEN_132; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_134 = _GEN_3825 & 4'h6 == j[3:0] ? solution_0_6 : _GEN_133; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_135 = _GEN_3825 & 4'h7 == j[3:0] ? solution_0_7 : _GEN_134; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_136 = _GEN_3825 & 4'h8 == j[3:0] ? 16'h0 : _GEN_135; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_137 = _GEN_3839 & 4'h0 == j[3:0] ? solution_1_0 : _GEN_136; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_138 = _GEN_3839 & 4'h1 == j[3:0] ? solution_1_1 : _GEN_137; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_139 = _GEN_3839 & 4'h2 == j[3:0] ? solution_1_2 : _GEN_138; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_140 = _GEN_3839 & 4'h3 == j[3:0] ? solution_1_3 : _GEN_139; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_141 = _GEN_3839 & 4'h4 == j[3:0] ? solution_1_4 : _GEN_140; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_142 = _GEN_3839 & 4'h5 == j[3:0] ? solution_1_5 : _GEN_141; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_143 = _GEN_3839 & 4'h6 == j[3:0] ? solution_1_6 : _GEN_142; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_144 = _GEN_3839 & 4'h7 == j[3:0] ? solution_1_7 : _GEN_143; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_145 = _GEN_3839 & 4'h8 == j[3:0] ? 16'h0 : _GEN_144; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_146 = _GEN_3855 & 4'h0 == j[3:0] ? solution_2_0 : _GEN_145; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_147 = _GEN_3855 & 4'h1 == j[3:0] ? solution_2_1 : _GEN_146; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_148 = _GEN_3855 & 4'h2 == j[3:0] ? solution_2_2 : _GEN_147; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_149 = _GEN_3855 & 4'h3 == j[3:0] ? solution_2_3 : _GEN_148; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_150 = _GEN_3855 & 4'h4 == j[3:0] ? solution_2_4 : _GEN_149; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_151 = _GEN_3855 & 4'h5 == j[3:0] ? solution_2_5 : _GEN_150; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_152 = _GEN_3855 & 4'h6 == j[3:0] ? solution_2_6 : _GEN_151; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_153 = _GEN_3855 & 4'h7 == j[3:0] ? solution_2_7 : _GEN_152; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_154 = _GEN_3855 & 4'h8 == j[3:0] ? 16'h0 : _GEN_153; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_155 = _GEN_3871 & 4'h0 == j[3:0] ? solution_3_0 : _GEN_154; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_156 = _GEN_3871 & 4'h1 == j[3:0] ? solution_3_1 : _GEN_155; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_157 = _GEN_3871 & 4'h2 == j[3:0] ? solution_3_2 : _GEN_156; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_158 = _GEN_3871 & 4'h3 == j[3:0] ? solution_3_3 : _GEN_157; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_159 = _GEN_3871 & 4'h4 == j[3:0] ? solution_3_4 : _GEN_158; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_160 = _GEN_3871 & 4'h5 == j[3:0] ? solution_3_5 : _GEN_159; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_161 = _GEN_3871 & 4'h6 == j[3:0] ? solution_3_6 : _GEN_160; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_162 = _GEN_3871 & 4'h7 == j[3:0] ? solution_3_7 : _GEN_161; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_163 = _GEN_3871 & 4'h8 == j[3:0] ? 16'h0 : _GEN_162; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_164 = _GEN_3887 & 4'h0 == j[3:0] ? solution_4_0 : _GEN_163; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_165 = _GEN_3887 & 4'h1 == j[3:0] ? solution_4_1 : _GEN_164; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_166 = _GEN_3887 & 4'h2 == j[3:0] ? solution_4_2 : _GEN_165; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_167 = _GEN_3887 & 4'h3 == j[3:0] ? solution_4_3 : _GEN_166; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_168 = _GEN_3887 & 4'h4 == j[3:0] ? solution_4_4 : _GEN_167; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_169 = _GEN_3887 & 4'h5 == j[3:0] ? solution_4_5 : _GEN_168; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_170 = _GEN_3887 & 4'h6 == j[3:0] ? solution_4_6 : _GEN_169; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_171 = _GEN_3887 & 4'h7 == j[3:0] ? solution_4_7 : _GEN_170; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_172 = _GEN_3887 & 4'h8 == j[3:0] ? 16'h0 : _GEN_171; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_173 = _GEN_3903 & 4'h0 == j[3:0] ? solution_5_0 : _GEN_172; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_174 = _GEN_3903 & 4'h1 == j[3:0] ? solution_5_1 : _GEN_173; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_175 = _GEN_3903 & 4'h2 == j[3:0] ? solution_5_2 : _GEN_174; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_176 = _GEN_3903 & 4'h3 == j[3:0] ? solution_5_3 : _GEN_175; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_177 = _GEN_3903 & 4'h4 == j[3:0] ? solution_5_4 : _GEN_176; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_178 = _GEN_3903 & 4'h5 == j[3:0] ? solution_5_5 : _GEN_177; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_179 = _GEN_3903 & 4'h6 == j[3:0] ? solution_5_6 : _GEN_178; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_180 = _GEN_3903 & 4'h7 == j[3:0] ? solution_5_7 : _GEN_179; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_181 = _GEN_3903 & 4'h8 == j[3:0] ? 16'h0 : _GEN_180; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_182 = _GEN_3919 & 4'h0 == j[3:0] ? solution_6_0 : _GEN_181; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_183 = _GEN_3919 & 4'h1 == j[3:0] ? solution_6_1 : _GEN_182; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_184 = _GEN_3919 & 4'h2 == j[3:0] ? solution_6_2 : _GEN_183; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_185 = _GEN_3919 & 4'h3 == j[3:0] ? solution_6_3 : _GEN_184; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_186 = _GEN_3919 & 4'h4 == j[3:0] ? solution_6_4 : _GEN_185; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_187 = _GEN_3919 & 4'h5 == j[3:0] ? solution_6_5 : _GEN_186; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_188 = _GEN_3919 & 4'h6 == j[3:0] ? solution_6_6 : _GEN_187; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_189 = _GEN_3919 & 4'h7 == j[3:0] ? solution_6_7 : _GEN_188; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_190 = _GEN_3919 & 4'h8 == j[3:0] ? 16'h0 : _GEN_189; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_191 = _GEN_3935 & 4'h0 == j[3:0] ? solution_7_0 : _GEN_190; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_192 = _GEN_3935 & 4'h1 == j[3:0] ? solution_7_1 : _GEN_191; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_193 = _GEN_3935 & 4'h2 == j[3:0] ? solution_7_2 : _GEN_192; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_194 = _GEN_3935 & 4'h3 == j[3:0] ? solution_7_3 : _GEN_193; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_195 = _GEN_3935 & 4'h4 == j[3:0] ? solution_7_4 : _GEN_194; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_196 = _GEN_3935 & 4'h5 == j[3:0] ? solution_7_5 : _GEN_195; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_197 = _GEN_3935 & 4'h6 == j[3:0] ? solution_7_6 : _GEN_196; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_198 = _GEN_3935 & 4'h7 == j[3:0] ? solution_7_7 : _GEN_197; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_199 = _GEN_3935 & 4'h8 == j[3:0] ? 16'h0 : _GEN_198; // @[ivncontrol4.scala 65:{31,31}]
  wire [31:0] _GEN_201 = 3'h1 == i[2:0] ? count_1 : count_0; // @[ivncontrol4.scala 66:{33,33}]
  wire [31:0] _GEN_202 = 3'h2 == i[2:0] ? count_2 : _GEN_201; // @[ivncontrol4.scala 66:{33,33}]
  wire [31:0] _GEN_203 = 3'h3 == i[2:0] ? count_3 : _GEN_202; // @[ivncontrol4.scala 66:{33,33}]
  wire [31:0] _GEN_204 = 3'h4 == i[2:0] ? count_4 : _GEN_203; // @[ivncontrol4.scala 66:{33,33}]
  wire [31:0] _GEN_205 = 3'h5 == i[2:0] ? count_5 : _GEN_204; // @[ivncontrol4.scala 66:{33,33}]
  wire [31:0] _GEN_206 = 3'h6 == i[2:0] ? count_6 : _GEN_205; // @[ivncontrol4.scala 66:{33,33}]
  wire [31:0] _GEN_207 = 3'h7 == i[2:0] ? count_7 : _GEN_206; // @[ivncontrol4.scala 66:{33,33}]
  wire [31:0] _count_T_2 = _GEN_207 + 32'h1; // @[ivncontrol4.scala 66:33]
  wire [31:0] _GEN_208 = 3'h0 == i[2:0] ? _count_T_2 : count_0; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_209 = 3'h1 == i[2:0] ? _count_T_2 : count_1; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_210 = 3'h2 == i[2:0] ? _count_T_2 : count_2; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_211 = 3'h3 == i[2:0] ? _count_T_2 : count_3; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_212 = 3'h4 == i[2:0] ? _count_T_2 : count_4; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_213 = 3'h5 == i[2:0] ? _count_T_2 : count_5; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_214 = 3'h6 == i[2:0] ? _count_T_2 : count_6; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_215 = 3'h7 == i[2:0] ? _count_T_2 : count_7; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_216 = _GEN_199 != 16'h0 ? _GEN_208 : count_0; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_217 = _GEN_199 != 16'h0 ? _GEN_209 : count_1; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_218 = _GEN_199 != 16'h0 ? _GEN_210 : count_2; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_219 = _GEN_199 != 16'h0 ? _GEN_211 : count_3; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_220 = _GEN_199 != 16'h0 ? _GEN_212 : count_4; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_221 = _GEN_199 != 16'h0 ? _GEN_213 : count_5; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_222 = _GEN_199 != 16'h0 ? _GEN_214 : count_6; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_223 = _GEN_199 != 16'h0 ? _GEN_215 : count_7; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_224 = io_validpin ? _GEN_216 : count_0; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _GEN_225 = io_validpin ? _GEN_217 : count_1; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _GEN_226 = io_validpin ? _GEN_218 : count_2; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _GEN_227 = io_validpin ? _GEN_219 : count_3; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _GEN_228 = io_validpin ? _GEN_220 : count_4; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _GEN_229 = io_validpin ? _GEN_221 : count_5; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _GEN_230 = io_validpin ? _GEN_222 : count_6; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _GEN_231 = io_validpin ? _GEN_223 : count_7; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _i_T_1 = i + 32'h1; // @[ivncontrol4.scala 113:16]
  wire [31:0] _GEN_247 = i < 32'h7 & _io_ProcessValid_T_1 ? _i_T_1 : i; // @[ivncontrol4.scala 112:74 113:11 41:20]
  wire [31:0] _j_T_1 = j + 32'h1; // @[ivncontrol4.scala 118:16]
  wire [3:0] _GEN_264 = _io_ProcessValid_T & j == 32'h8 ? 4'h8 : 4'h0; // @[ivncontrol4.scala 120:77 121:11 129:11]
  wire [31:0] _GEN_265 = _io_ProcessValid_T & j == 32'h8 ? 32'h7 : _GEN_247; // @[ivncontrol4.scala 120:77 122:11]
  wire  _GEN_312 = _io_ProcessValid_T_2; // @[ivncontrol4.scala 153:41]
  wire [31:0] _GEN_313 = rowcount_0 != 32'h0 ? 32'h0 : pin; // @[ivncontrol4.scala 162:30 163:13 37:22]
  wire  _T_27 = rowcount_0 == 32'h0; // @[ivncontrol4.scala 165:23]
  wire [31:0] _GEN_314 = rowcount_0 == 32'h0 & rowcount_1 != 32'h0 ? 32'h1 : _GEN_313; // @[ivncontrol4.scala 165:54 166:13]
  wire  _T_32 = _T_27 & rowcount_1 == 32'h0; // @[ivncontrol4.scala 168:31]
  wire [31:0] _GEN_315 = _T_27 & rowcount_1 == 32'h0 & rowcount_2 != 32'h0 ? 32'h2 : _GEN_314; // @[ivncontrol4.scala 168:77 169:13]
  wire  _T_39 = _T_32 & rowcount_2 == 32'h0; // @[ivncontrol4.scala 171:54]
  wire [31:0] _GEN_316 = _T_32 & rowcount_2 == 32'h0 & rowcount_3 != 32'h0 ? 32'h3 : _GEN_315; // @[ivncontrol4.scala 171:100 172:13]
  wire  _T_48 = _T_39 & rowcount_3 == 32'h0; // @[ivncontrol4.scala 174:77]
  wire [31:0] _GEN_317 = _T_39 & rowcount_3 == 32'h0 & rowcount_4 != 32'h0 ? 32'h4 : _GEN_316; // @[ivncontrol4.scala 174:123 175:13]
  wire  _T_59 = _T_48 & rowcount_4 == 32'h0; // @[ivncontrol4.scala 177:100]
  wire  _T_72 = _T_59 & rowcount_5 == 32'h0; // @[ivncontrol4.scala 180:123]
  wire  valid = _io_ProcessValid_T_2; // @[ivncontrol4.scala 153:41]
  wire [32:0] _T_91 = {{1'd0}, pin}; // @[ivncontrol4.scala 191:27]
  wire [31:0] _GEN_322 = 4'h1 == _T_91[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_323 = 4'h2 == _T_91[3:0] ? rowcount_2 : _GEN_322; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_324 = 4'h3 == _T_91[3:0] ? rowcount_3 : _GEN_323; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_325 = 4'h4 == _T_91[3:0] ? rowcount_4 : _GEN_324; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_326 = 4'h5 == _T_91[3:0] ? rowcount_5 : _GEN_325; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_327 = 4'h6 == _T_91[3:0] ? rowcount_6 : _GEN_326; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_328 = 4'h7 == _T_91[3:0] ? rowcount_7 : _GEN_327; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_329 = 4'h8 == _T_91[3:0] ? rowcount_8 : _GEN_328; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_330 = 4'h9 == _T_91[3:0] ? rowcount_9 : _GEN_329; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_331 = 4'ha == _T_91[3:0] ? rowcount_10 : _GEN_330; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_332 = 4'hb == _T_91[3:0] ? rowcount_11 : _GEN_331; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_333 = 4'hc == _T_91[3:0] ? rowcount_12 : _GEN_332; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_334 = 4'hd == _T_91[3:0] ? rowcount_13 : _GEN_333; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_335 = 4'he == _T_91[3:0] ? rowcount_14 : _GEN_334; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_336 = 4'hf == _T_91[3:0] ? rowcount_15 : _GEN_335; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_449 = _GEN_336 == 32'h1 ? _T_91[31:0] : 32'h19; // @[ivncontrol4.scala 142:17 241:50 242:21]
  wire [31:0] _GEN_450 = _GEN_336 == 32'h2 ? _T_91[31:0] : _GEN_449; // @[ivncontrol4.scala 237:51 238:21]
  wire [31:0] _GEN_451 = _GEN_336 == 32'h2 ? _T_91[31:0] : 32'h3; // @[ivncontrol4.scala 142:17 237:51 239:21]
  wire [31:0] _GEN_452 = _GEN_336 == 32'h3 ? _T_91[31:0] : _GEN_450; // @[ivncontrol4.scala 232:50 233:21]
  wire [31:0] _GEN_453 = _GEN_336 == 32'h3 ? _T_91[31:0] : _GEN_451; // @[ivncontrol4.scala 232:50 234:21]
  wire [31:0] _GEN_454 = _GEN_336 == 32'h3 ? _T_91[31:0] : 32'h1c; // @[ivncontrol4.scala 142:17 232:50 235:21]
  wire [31:0] _GEN_455 = _GEN_336 == 32'h4 ? _T_91[31:0] : _GEN_452; // @[ivncontrol4.scala 224:50 225:21]
  wire [31:0] _GEN_456 = _GEN_336 == 32'h4 ? _T_91[31:0] : _GEN_453; // @[ivncontrol4.scala 224:50 226:21]
  wire [31:0] _GEN_457 = _GEN_336 == 32'h4 ? _T_91[31:0] : _GEN_454; // @[ivncontrol4.scala 224:50 227:21]
  wire [31:0] _GEN_458 = _GEN_336 == 32'h4 ? _T_91[31:0] : 32'h4; // @[ivncontrol4.scala 142:17 224:50 228:21]
  wire [31:0] _GEN_459 = _GEN_336 == 32'h5 ? _T_91[31:0] : _GEN_455; // @[ivncontrol4.scala 217:50 218:21]
  wire [31:0] _GEN_460 = _GEN_336 == 32'h5 ? _T_91[31:0] : _GEN_456; // @[ivncontrol4.scala 217:50 219:21]
  wire [31:0] _GEN_461 = _GEN_336 == 32'h5 ? _T_91[31:0] : _GEN_457; // @[ivncontrol4.scala 217:50 220:21]
  wire [31:0] _GEN_462 = _GEN_336 == 32'h5 ? _T_91[31:0] : _GEN_458; // @[ivncontrol4.scala 217:50 221:21]
  wire [31:0] _GEN_463 = _GEN_336 == 32'h5 ? _T_91[31:0] : 32'h14; // @[ivncontrol4.scala 143:18 217:50 222:22]
  wire [31:0] _GEN_464 = _GEN_336 == 32'h6 ? _T_91[31:0] : _GEN_459; // @[ivncontrol4.scala 209:52 210:21]
  wire [31:0] _GEN_465 = _GEN_336 == 32'h6 ? _T_91[31:0] : _GEN_460; // @[ivncontrol4.scala 209:52 211:21]
  wire [31:0] _GEN_466 = _GEN_336 == 32'h6 ? _T_91[31:0] : _GEN_461; // @[ivncontrol4.scala 209:52 212:21]
  wire [31:0] _GEN_467 = _GEN_336 == 32'h6 ? _T_91[31:0] : _GEN_462; // @[ivncontrol4.scala 209:52 213:21]
  wire [31:0] _GEN_468 = _GEN_336 == 32'h6 ? _T_91[31:0] : _GEN_463; // @[ivncontrol4.scala 209:52 214:22]
  wire [31:0] _GEN_469 = _GEN_336 == 32'h6 ? _T_91[31:0] : 32'h1b; // @[ivncontrol4.scala 143:18 209:52 215:22]
  wire [31:0] _GEN_470 = _GEN_336 == 32'h7 ? _T_91[31:0] : _GEN_464; // @[ivncontrol4.scala 201:52 202:21]
  wire [31:0] _GEN_471 = _GEN_336 == 32'h7 ? _T_91[31:0] : _GEN_465; // @[ivncontrol4.scala 201:52 203:21]
  wire [31:0] _GEN_472 = _GEN_336 == 32'h7 ? _T_91[31:0] : _GEN_466; // @[ivncontrol4.scala 201:52 204:21]
  wire [31:0] _GEN_473 = _GEN_336 == 32'h7 ? _T_91[31:0] : _GEN_467; // @[ivncontrol4.scala 201:52 205:21]
  wire [31:0] _GEN_474 = _GEN_336 == 32'h7 ? _T_91[31:0] : _GEN_468; // @[ivncontrol4.scala 201:52 206:22]
  wire [31:0] _GEN_475 = _GEN_336 == 32'h7 ? _T_91[31:0] : _GEN_469; // @[ivncontrol4.scala 201:52 207:22]
  wire [31:0] _GEN_476 = _GEN_336 == 32'h7 ? _T_91[31:0] : 32'h5; // @[ivncontrol4.scala 143:18 201:52 208:22]
  wire [31:0] _GEN_477 = _GEN_336 >= 32'h8 ? _T_91[31:0] : _GEN_470; // @[ivncontrol4.scala 191:42 192:21]
  wire [31:0] _GEN_478 = _GEN_336 >= 32'h8 ? _T_91[31:0] : _GEN_471; // @[ivncontrol4.scala 191:42 193:21]
  wire [31:0] _GEN_479 = _GEN_336 >= 32'h8 ? _T_91[31:0] : _GEN_472; // @[ivncontrol4.scala 191:42 194:21]
  wire [31:0] _GEN_480 = _GEN_336 >= 32'h8 ? _T_91[31:0] : _GEN_473; // @[ivncontrol4.scala 191:42 195:21]
  wire [31:0] _GEN_481 = _GEN_336 >= 32'h8 ? _T_91[31:0] : _GEN_474; // @[ivncontrol4.scala 191:42 196:22]
  wire [31:0] _GEN_482 = _GEN_336 >= 32'h8 ? _T_91[31:0] : _GEN_475; // @[ivncontrol4.scala 191:42 197:22]
  wire [31:0] _GEN_483 = _GEN_336 >= 32'h8 ? _T_91[31:0] : _GEN_476; // @[ivncontrol4.scala 191:42 198:22]
  wire [31:0] _GEN_484 = _GEN_336 >= 32'h8 ? _T_91[31:0] : 32'h8; // @[ivncontrol4.scala 143:18 191:42 199:22]
  wire [31:0] _T_127 = 32'h8 - _GEN_336; // @[ivncontrol4.scala 245:18]
  wire [31:0] _i_vn_1_T_15 = 32'h1 + pin; // @[ivncontrol4.scala 246:29]
  wire [31:0] _GEN_597 = _T_127 == 32'h1 ? _i_vn_1_T_15 : _GEN_484; // @[ivncontrol4.scala 286:54 289:22]
  wire [31:0] _GEN_598 = _T_127 == 32'h2 ? _i_vn_1_T_15 : _GEN_483; // @[ivncontrol4.scala 281:54 284:22]
  wire [31:0] _GEN_599 = _T_127 == 32'h2 ? _i_vn_1_T_15 : _GEN_597; // @[ivncontrol4.scala 281:54 285:22]
  wire [31:0] _GEN_600 = _T_127 == 32'h3 ? _i_vn_1_T_15 : _GEN_482; // @[ivncontrol4.scala 274:54 276:22]
  wire [31:0] _GEN_601 = _T_127 == 32'h3 ? _i_vn_1_T_15 : _GEN_598; // @[ivncontrol4.scala 274:54 277:22]
  wire [31:0] _GEN_602 = _T_127 == 32'h3 ? _i_vn_1_T_15 : _GEN_599; // @[ivncontrol4.scala 274:54 278:22]
  wire [31:0] _GEN_603 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_481; // @[ivncontrol4.scala 268:54 270:22]
  wire [31:0] _GEN_604 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_600; // @[ivncontrol4.scala 268:54 271:22]
  wire [31:0] _GEN_605 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_601; // @[ivncontrol4.scala 268:54 272:22]
  wire [31:0] _GEN_606 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_602; // @[ivncontrol4.scala 268:54 273:22]
  wire [31:0] _GEN_607 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_480; // @[ivncontrol4.scala 261:54 263:21]
  wire [31:0] _GEN_608 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_603; // @[ivncontrol4.scala 261:54 264:22]
  wire [31:0] _GEN_609 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_604; // @[ivncontrol4.scala 261:54 265:22]
  wire [31:0] _GEN_610 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_605; // @[ivncontrol4.scala 261:54 266:22]
  wire [31:0] _GEN_611 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_606; // @[ivncontrol4.scala 261:54 267:22]
  wire [31:0] _GEN_612 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_479; // @[ivncontrol4.scala 254:54 255:22]
  wire [31:0] _GEN_613 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_607; // @[ivncontrol4.scala 254:54 256:21]
  wire [31:0] _GEN_614 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_608; // @[ivncontrol4.scala 254:54 257:22]
  wire [31:0] _GEN_615 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_609; // @[ivncontrol4.scala 254:54 258:22]
  wire [31:0] _GEN_616 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_610; // @[ivncontrol4.scala 254:54 259:22]
  wire [31:0] _GEN_617 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_611; // @[ivncontrol4.scala 254:54 260:22]
  wire [31:0] _GEN_618 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_478; // @[ivncontrol4.scala 245:49 246:22]
  wire [31:0] _GEN_619 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_612; // @[ivncontrol4.scala 245:49 247:21]
  wire [31:0] _GEN_620 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_613; // @[ivncontrol4.scala 245:49 248:21]
  wire [31:0] _GEN_621 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_614; // @[ivncontrol4.scala 245:49 249:22]
  wire [31:0] _GEN_622 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_615; // @[ivncontrol4.scala 245:49 250:22]
  wire [31:0] _GEN_623 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_616; // @[ivncontrol4.scala 245:49 251:22]
  wire [31:0] _GEN_624 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_617; // @[ivncontrol4.scala 245:49 252:22]
  wire [31:0] _GEN_642 = 4'h1 == _i_vn_1_T_15[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_643 = 4'h2 == _i_vn_1_T_15[3:0] ? rowcount_2 : _GEN_642; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_644 = 4'h3 == _i_vn_1_T_15[3:0] ? rowcount_3 : _GEN_643; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_645 = 4'h4 == _i_vn_1_T_15[3:0] ? rowcount_4 : _GEN_644; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_646 = 4'h5 == _i_vn_1_T_15[3:0] ? rowcount_5 : _GEN_645; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_647 = 4'h6 == _i_vn_1_T_15[3:0] ? rowcount_6 : _GEN_646; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_648 = 4'h7 == _i_vn_1_T_15[3:0] ? rowcount_7 : _GEN_647; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_649 = 4'h8 == _i_vn_1_T_15[3:0] ? rowcount_8 : _GEN_648; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_650 = 4'h9 == _i_vn_1_T_15[3:0] ? rowcount_9 : _GEN_649; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_651 = 4'ha == _i_vn_1_T_15[3:0] ? rowcount_10 : _GEN_650; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_652 = 4'hb == _i_vn_1_T_15[3:0] ? rowcount_11 : _GEN_651; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_653 = 4'hc == _i_vn_1_T_15[3:0] ? rowcount_12 : _GEN_652; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_654 = 4'hd == _i_vn_1_T_15[3:0] ? rowcount_13 : _GEN_653; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_655 = 4'he == _i_vn_1_T_15[3:0] ? rowcount_14 : _GEN_654; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_656 = 4'hf == _i_vn_1_T_15[3:0] ? rowcount_15 : _GEN_655; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _T_172 = _GEN_336 + _GEN_656; // @[ivncontrol4.scala 292:41]
  wire [31:0] _T_174 = 32'h8 - _T_172; // @[ivncontrol4.scala 292:18]
  wire [31:0] _i_vn_1_T_17 = 32'h2 + pin; // @[ivncontrol4.scala 293:29]
  wire [31:0] _GEN_849 = _T_174 == 32'h1 ? _i_vn_1_T_17 : _GEN_624; // @[ivncontrol4.scala 335:78 338:22]
  wire [31:0] _GEN_850 = _T_174 == 32'h2 ? _i_vn_1_T_17 : _GEN_623; // @[ivncontrol4.scala 329:76 332:22]
  wire [31:0] _GEN_851 = _T_174 == 32'h2 ? _i_vn_1_T_17 : _GEN_849; // @[ivncontrol4.scala 329:76 333:22]
  wire [31:0] _GEN_852 = _T_174 == 32'h3 ? _i_vn_1_T_17 : _GEN_622; // @[ivncontrol4.scala 322:78 324:23]
  wire [31:0] _GEN_853 = _T_174 == 32'h3 ? _i_vn_1_T_17 : _GEN_850; // @[ivncontrol4.scala 322:78 325:22]
  wire [31:0] _GEN_854 = _T_174 == 32'h3 ? _i_vn_1_T_17 : _GEN_851; // @[ivncontrol4.scala 322:78 326:22]
  wire [31:0] _GEN_855 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_621; // @[ivncontrol4.scala 316:78 318:22]
  wire [31:0] _GEN_856 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_852; // @[ivncontrol4.scala 316:78 319:22]
  wire [31:0] _GEN_857 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_853; // @[ivncontrol4.scala 316:78 320:22]
  wire [31:0] _GEN_858 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_854; // @[ivncontrol4.scala 316:78 321:22]
  wire [31:0] _GEN_859 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_620; // @[ivncontrol4.scala 309:76 311:23]
  wire [31:0] _GEN_860 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_855; // @[ivncontrol4.scala 309:76 312:22]
  wire [31:0] _GEN_861 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_856; // @[ivncontrol4.scala 309:76 313:22]
  wire [31:0] _GEN_862 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_857; // @[ivncontrol4.scala 309:76 314:22]
  wire [31:0] _GEN_863 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_858; // @[ivncontrol4.scala 309:76 315:22]
  wire [31:0] _GEN_864 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_619; // @[ivncontrol4.scala 301:77 303:22]
  wire [31:0] _GEN_865 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_859; // @[ivncontrol4.scala 301:77 304:21]
  wire [31:0] _GEN_866 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_860; // @[ivncontrol4.scala 301:77 305:22]
  wire [31:0] _GEN_867 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_861; // @[ivncontrol4.scala 301:77 306:22]
  wire [31:0] _GEN_868 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_862; // @[ivncontrol4.scala 301:77 307:22]
  wire [31:0] _GEN_869 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_863; // @[ivncontrol4.scala 301:77 308:22]
  wire [31:0] _GEN_870 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_618; // @[ivncontrol4.scala 292:73 293:22]
  wire [31:0] _GEN_871 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_864; // @[ivncontrol4.scala 292:73 294:21]
  wire [31:0] _GEN_872 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_865; // @[ivncontrol4.scala 292:73 295:21]
  wire [31:0] _GEN_873 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_866; // @[ivncontrol4.scala 292:73 296:22]
  wire [31:0] _GEN_874 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_867; // @[ivncontrol4.scala 292:73 297:22]
  wire [31:0] _GEN_875 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_868; // @[ivncontrol4.scala 292:73 298:22]
  wire [31:0] _GEN_876 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_869; // @[ivncontrol4.scala 292:73 299:22]
  wire [31:0] _GEN_910 = 4'h1 == _i_vn_1_T_17[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_911 = 4'h2 == _i_vn_1_T_17[3:0] ? rowcount_2 : _GEN_910; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_912 = 4'h3 == _i_vn_1_T_17[3:0] ? rowcount_3 : _GEN_911; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_913 = 4'h4 == _i_vn_1_T_17[3:0] ? rowcount_4 : _GEN_912; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_914 = 4'h5 == _i_vn_1_T_17[3:0] ? rowcount_5 : _GEN_913; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_915 = 4'h6 == _i_vn_1_T_17[3:0] ? rowcount_6 : _GEN_914; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_916 = 4'h7 == _i_vn_1_T_17[3:0] ? rowcount_7 : _GEN_915; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_917 = 4'h8 == _i_vn_1_T_17[3:0] ? rowcount_8 : _GEN_916; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_918 = 4'h9 == _i_vn_1_T_17[3:0] ? rowcount_9 : _GEN_917; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_919 = 4'ha == _i_vn_1_T_17[3:0] ? rowcount_10 : _GEN_918; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_920 = 4'hb == _i_vn_1_T_17[3:0] ? rowcount_11 : _GEN_919; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_921 = 4'hc == _i_vn_1_T_17[3:0] ? rowcount_12 : _GEN_920; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_922 = 4'hd == _i_vn_1_T_17[3:0] ? rowcount_13 : _GEN_921; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_923 = 4'he == _i_vn_1_T_17[3:0] ? rowcount_14 : _GEN_922; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_924 = 4'hf == _i_vn_1_T_17[3:0] ? rowcount_15 : _GEN_923; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _T_254 = _T_172 + _GEN_924; // @[ivncontrol4.scala 343:62]
  wire [31:0] _T_256 = 32'h8 - _T_254; // @[ivncontrol4.scala 343:17]
  wire [31:0] _i_vn_1_T_19 = 32'h3 + pin; // @[ivncontrol4.scala 344:29]
  wire [31:0] _GEN_1213 = _T_256 == 32'h1 ? _i_vn_1_T_19 : _GEN_876; // @[ivncontrol4.scala 386:100 389:22]
  wire [31:0] _GEN_1214 = _T_256 == 32'h2 ? _i_vn_1_T_19 : _GEN_875; // @[ivncontrol4.scala 380:98 383:22]
  wire [31:0] _GEN_1215 = _T_256 == 32'h2 ? _i_vn_1_T_19 : _GEN_1213; // @[ivncontrol4.scala 380:98 384:22]
  wire [31:0] _GEN_1216 = _T_256 == 32'h3 ? _i_vn_1_T_19 : _GEN_874; // @[ivncontrol4.scala 373:100 375:23]
  wire [31:0] _GEN_1217 = _T_256 == 32'h3 ? _i_vn_1_T_19 : _GEN_1214; // @[ivncontrol4.scala 373:100 376:22]
  wire [31:0] _GEN_1218 = _T_256 == 32'h3 ? _i_vn_1_T_19 : _GEN_1215; // @[ivncontrol4.scala 373:100 377:22]
  wire [31:0] _GEN_1219 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_873; // @[ivncontrol4.scala 367:100 369:22]
  wire [31:0] _GEN_1220 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_1216; // @[ivncontrol4.scala 367:100 370:22]
  wire [31:0] _GEN_1221 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_1217; // @[ivncontrol4.scala 367:100 371:22]
  wire [31:0] _GEN_1222 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_1218; // @[ivncontrol4.scala 367:100 372:22]
  wire [31:0] _GEN_1223 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_872; // @[ivncontrol4.scala 360:98 362:23]
  wire [31:0] _GEN_1224 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1219; // @[ivncontrol4.scala 360:98 363:22]
  wire [31:0] _GEN_1225 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1220; // @[ivncontrol4.scala 360:98 364:22]
  wire [31:0] _GEN_1226 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1221; // @[ivncontrol4.scala 360:98 365:22]
  wire [31:0] _GEN_1227 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1222; // @[ivncontrol4.scala 360:98 366:22]
  wire [31:0] _GEN_1228 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_871; // @[ivncontrol4.scala 352:99 354:22]
  wire [31:0] _GEN_1229 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1223; // @[ivncontrol4.scala 352:99 355:21]
  wire [31:0] _GEN_1230 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1224; // @[ivncontrol4.scala 352:99 356:22]
  wire [31:0] _GEN_1231 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1225; // @[ivncontrol4.scala 352:99 357:22]
  wire [31:0] _GEN_1232 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1226; // @[ivncontrol4.scala 352:99 358:22]
  wire [31:0] _GEN_1233 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1227; // @[ivncontrol4.scala 352:99 359:22]
  wire [31:0] _GEN_1234 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_870; // @[ivncontrol4.scala 343:94 344:22]
  wire [31:0] _GEN_1235 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1228; // @[ivncontrol4.scala 343:94 345:21]
  wire [31:0] _GEN_1236 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1229; // @[ivncontrol4.scala 343:94 346:21]
  wire [31:0] _GEN_1237 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1230; // @[ivncontrol4.scala 343:94 347:22]
  wire [31:0] _GEN_1238 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1231; // @[ivncontrol4.scala 343:94 348:22]
  wire [31:0] _GEN_1239 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1232; // @[ivncontrol4.scala 343:94 349:22]
  wire [31:0] _GEN_1240 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1233; // @[ivncontrol4.scala 343:94 350:22]
  wire [31:0] _GEN_1290 = 4'h1 == _i_vn_1_T_19[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1291 = 4'h2 == _i_vn_1_T_19[3:0] ? rowcount_2 : _GEN_1290; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1292 = 4'h3 == _i_vn_1_T_19[3:0] ? rowcount_3 : _GEN_1291; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1293 = 4'h4 == _i_vn_1_T_19[3:0] ? rowcount_4 : _GEN_1292; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1294 = 4'h5 == _i_vn_1_T_19[3:0] ? rowcount_5 : _GEN_1293; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1295 = 4'h6 == _i_vn_1_T_19[3:0] ? rowcount_6 : _GEN_1294; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1296 = 4'h7 == _i_vn_1_T_19[3:0] ? rowcount_7 : _GEN_1295; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1297 = 4'h8 == _i_vn_1_T_19[3:0] ? rowcount_8 : _GEN_1296; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1298 = 4'h9 == _i_vn_1_T_19[3:0] ? rowcount_9 : _GEN_1297; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1299 = 4'ha == _i_vn_1_T_19[3:0] ? rowcount_10 : _GEN_1298; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1300 = 4'hb == _i_vn_1_T_19[3:0] ? rowcount_11 : _GEN_1299; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1301 = 4'hc == _i_vn_1_T_19[3:0] ? rowcount_12 : _GEN_1300; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1302 = 4'hd == _i_vn_1_T_19[3:0] ? rowcount_13 : _GEN_1301; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1303 = 4'he == _i_vn_1_T_19[3:0] ? rowcount_14 : _GEN_1302; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1304 = 4'hf == _i_vn_1_T_19[3:0] ? rowcount_15 : _GEN_1303; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _T_371 = _T_254 + _GEN_1304; // @[ivncontrol4.scala 393:86]
  wire [31:0] _T_373 = 32'h8 - _T_371; // @[ivncontrol4.scala 393:19]
  wire [31:0] _i_vn_1_T_21 = 32'h4 + pin; // @[ivncontrol4.scala 394:29]
  wire [31:0] _GEN_1689 = _T_373 == 32'h1 ? _i_vn_1_T_21 : _GEN_1240; // @[ivncontrol4.scala 436:122 439:22]
  wire [31:0] _GEN_1690 = _T_373 == 32'h2 ? _i_vn_1_T_21 : _GEN_1239; // @[ivncontrol4.scala 430:121 433:22]
  wire [31:0] _GEN_1691 = _T_373 == 32'h2 ? _i_vn_1_T_21 : _GEN_1689; // @[ivncontrol4.scala 430:121 434:22]
  wire [31:0] _GEN_1692 = _T_373 == 32'h3 ? _i_vn_1_T_21 : _GEN_1238; // @[ivncontrol4.scala 423:123 425:23]
  wire [31:0] _GEN_1693 = _T_373 == 32'h3 ? _i_vn_1_T_21 : _GEN_1690; // @[ivncontrol4.scala 423:123 426:22]
  wire [31:0] _GEN_1694 = _T_373 == 32'h3 ? _i_vn_1_T_21 : _GEN_1691; // @[ivncontrol4.scala 423:123 427:22]
  wire [31:0] _GEN_1695 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1237; // @[ivncontrol4.scala 417:122 419:22]
  wire [31:0] _GEN_1696 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1692; // @[ivncontrol4.scala 417:122 420:22]
  wire [31:0] _GEN_1697 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1693; // @[ivncontrol4.scala 417:122 421:22]
  wire [31:0] _GEN_1698 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1694; // @[ivncontrol4.scala 417:122 422:22]
  wire [31:0] _GEN_1699 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1236; // @[ivncontrol4.scala 410:121 412:23]
  wire [31:0] _GEN_1700 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1695; // @[ivncontrol4.scala 410:121 413:22]
  wire [31:0] _GEN_1701 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1696; // @[ivncontrol4.scala 410:121 414:22]
  wire [31:0] _GEN_1702 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1697; // @[ivncontrol4.scala 410:121 415:22]
  wire [31:0] _GEN_1703 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1698; // @[ivncontrol4.scala 410:121 416:22]
  wire [31:0] _GEN_1704 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1235; // @[ivncontrol4.scala 402:121 404:22]
  wire [31:0] _GEN_1705 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1699; // @[ivncontrol4.scala 402:121 405:21]
  wire [31:0] _GEN_1706 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1700; // @[ivncontrol4.scala 402:121 406:22]
  wire [31:0] _GEN_1707 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1701; // @[ivncontrol4.scala 402:121 407:22]
  wire [31:0] _GEN_1708 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1702; // @[ivncontrol4.scala 402:121 408:22]
  wire [31:0] _GEN_1709 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1703; // @[ivncontrol4.scala 402:121 409:22]
  wire [31:0] _GEN_1710 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1234; // @[ivncontrol4.scala 393:118 394:22]
  wire [31:0] _GEN_1711 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1704; // @[ivncontrol4.scala 393:118 395:21]
  wire [31:0] _GEN_1712 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1705; // @[ivncontrol4.scala 393:118 396:21]
  wire [31:0] _GEN_1713 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1706; // @[ivncontrol4.scala 393:118 397:22]
  wire [31:0] _GEN_1714 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1707; // @[ivncontrol4.scala 393:118 398:22]
  wire [31:0] _GEN_1715 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1708; // @[ivncontrol4.scala 393:118 399:22]
  wire [31:0] _GEN_1716 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1709; // @[ivncontrol4.scala 393:118 400:22]
  wire [31:0] _GEN_1782 = 4'h1 == _i_vn_1_T_21[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1783 = 4'h2 == _i_vn_1_T_21[3:0] ? rowcount_2 : _GEN_1782; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1784 = 4'h3 == _i_vn_1_T_21[3:0] ? rowcount_3 : _GEN_1783; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1785 = 4'h4 == _i_vn_1_T_21[3:0] ? rowcount_4 : _GEN_1784; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1786 = 4'h5 == _i_vn_1_T_21[3:0] ? rowcount_5 : _GEN_1785; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1787 = 4'h6 == _i_vn_1_T_21[3:0] ? rowcount_6 : _GEN_1786; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1788 = 4'h7 == _i_vn_1_T_21[3:0] ? rowcount_7 : _GEN_1787; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1789 = 4'h8 == _i_vn_1_T_21[3:0] ? rowcount_8 : _GEN_1788; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1790 = 4'h9 == _i_vn_1_T_21[3:0] ? rowcount_9 : _GEN_1789; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1791 = 4'ha == _i_vn_1_T_21[3:0] ? rowcount_10 : _GEN_1790; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1792 = 4'hb == _i_vn_1_T_21[3:0] ? rowcount_11 : _GEN_1791; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1793 = 4'hc == _i_vn_1_T_21[3:0] ? rowcount_12 : _GEN_1792; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1794 = 4'hd == _i_vn_1_T_21[3:0] ? rowcount_13 : _GEN_1793; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1795 = 4'he == _i_vn_1_T_21[3:0] ? rowcount_14 : _GEN_1794; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1796 = 4'hf == _i_vn_1_T_21[3:0] ? rowcount_15 : _GEN_1795; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _T_523 = _T_371 + _GEN_1796; // @[ivncontrol4.scala 443:108]
  wire [31:0] _T_525 = 32'h8 - _T_523; // @[ivncontrol4.scala 443:19]
  wire [31:0] _i_vn_1_T_23 = 32'h5 + pin; // @[ivncontrol4.scala 444:29]
  wire [31:0] _GEN_2277 = _T_525 == 32'h1 ? _i_vn_1_T_23 : _GEN_1716; // @[ivncontrol4.scala 486:144 489:22]
  wire [31:0] _GEN_2278 = _T_525 == 32'h2 ? _i_vn_1_T_23 : _GEN_1715; // @[ivncontrol4.scala 480:143 483:22]
  wire [31:0] _GEN_2279 = _T_525 == 32'h2 ? _i_vn_1_T_23 : _GEN_2277; // @[ivncontrol4.scala 480:143 484:22]
  wire [31:0] _GEN_2280 = _T_525 == 32'h3 ? _i_vn_1_T_23 : _GEN_1714; // @[ivncontrol4.scala 473:145 475:23]
  wire [31:0] _GEN_2281 = _T_525 == 32'h3 ? _i_vn_1_T_23 : _GEN_2278; // @[ivncontrol4.scala 473:145 476:22]
  wire [31:0] _GEN_2282 = _T_525 == 32'h3 ? _i_vn_1_T_23 : _GEN_2279; // @[ivncontrol4.scala 473:145 477:22]
  wire [31:0] _GEN_2283 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_1713; // @[ivncontrol4.scala 467:143 469:22]
  wire [31:0] _GEN_2284 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_2280; // @[ivncontrol4.scala 467:143 470:22]
  wire [31:0] _GEN_2285 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_2281; // @[ivncontrol4.scala 467:143 471:22]
  wire [31:0] _GEN_2286 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_2282; // @[ivncontrol4.scala 467:143 472:22]
  wire [31:0] _GEN_2287 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_1712; // @[ivncontrol4.scala 460:143 462:23]
  wire [31:0] _GEN_2288 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2283; // @[ivncontrol4.scala 460:143 463:22]
  wire [31:0] _GEN_2289 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2284; // @[ivncontrol4.scala 460:143 464:22]
  wire [31:0] _GEN_2290 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2285; // @[ivncontrol4.scala 460:143 465:22]
  wire [31:0] _GEN_2291 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2286; // @[ivncontrol4.scala 460:143 466:22]
  wire [31:0] _GEN_2292 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_1711; // @[ivncontrol4.scala 452:143 454:22]
  wire [31:0] _GEN_2293 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2287; // @[ivncontrol4.scala 452:143 455:21]
  wire [31:0] _GEN_2294 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2288; // @[ivncontrol4.scala 452:143 456:22]
  wire [31:0] _GEN_2295 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2289; // @[ivncontrol4.scala 452:143 457:22]
  wire [31:0] _GEN_2296 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2290; // @[ivncontrol4.scala 452:143 458:22]
  wire [31:0] _GEN_2297 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2291; // @[ivncontrol4.scala 452:143 459:22]
  wire [31:0] _GEN_2298 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_1710; // @[ivncontrol4.scala 443:140 444:22]
  wire [31:0] _GEN_2299 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2292; // @[ivncontrol4.scala 443:140 445:21]
  wire [31:0] _GEN_2300 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2293; // @[ivncontrol4.scala 443:140 446:21]
  wire [31:0] _GEN_2301 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2294; // @[ivncontrol4.scala 443:140 447:22]
  wire [31:0] _GEN_2302 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2295; // @[ivncontrol4.scala 443:140 448:22]
  wire [31:0] _GEN_2303 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2296; // @[ivncontrol4.scala 443:140 449:22]
  wire [31:0] _GEN_2304 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2297; // @[ivncontrol4.scala 443:140 450:22]
  wire [31:0] _GEN_2386 = 4'h1 == _i_vn_1_T_23[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2387 = 4'h2 == _i_vn_1_T_23[3:0] ? rowcount_2 : _GEN_2386; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2388 = 4'h3 == _i_vn_1_T_23[3:0] ? rowcount_3 : _GEN_2387; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2389 = 4'h4 == _i_vn_1_T_23[3:0] ? rowcount_4 : _GEN_2388; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2390 = 4'h5 == _i_vn_1_T_23[3:0] ? rowcount_5 : _GEN_2389; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2391 = 4'h6 == _i_vn_1_T_23[3:0] ? rowcount_6 : _GEN_2390; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2392 = 4'h7 == _i_vn_1_T_23[3:0] ? rowcount_7 : _GEN_2391; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2393 = 4'h8 == _i_vn_1_T_23[3:0] ? rowcount_8 : _GEN_2392; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2394 = 4'h9 == _i_vn_1_T_23[3:0] ? rowcount_9 : _GEN_2393; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2395 = 4'ha == _i_vn_1_T_23[3:0] ? rowcount_10 : _GEN_2394; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2396 = 4'hb == _i_vn_1_T_23[3:0] ? rowcount_11 : _GEN_2395; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2397 = 4'hc == _i_vn_1_T_23[3:0] ? rowcount_12 : _GEN_2396; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2398 = 4'hd == _i_vn_1_T_23[3:0] ? rowcount_13 : _GEN_2397; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2399 = 4'he == _i_vn_1_T_23[3:0] ? rowcount_14 : _GEN_2398; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2400 = 4'hf == _i_vn_1_T_23[3:0] ? rowcount_15 : _GEN_2399; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _T_710 = _T_523 + _GEN_2400; // @[ivncontrol4.scala 494:130]
  wire [31:0] _T_712 = 32'h8 - _T_710; // @[ivncontrol4.scala 494:19]
  wire [31:0] _i_vn_1_T_25 = 32'h6 + pin; // @[ivncontrol4.scala 495:29]
  wire [31:0] _GEN_2977 = _T_712 == 32'h1 ? _i_vn_1_T_25 : _GEN_2304; // @[ivncontrol4.scala 537:166 540:22]
  wire [31:0] _GEN_2978 = _T_712 == 32'h2 ? _i_vn_1_T_25 : _GEN_2303; // @[ivncontrol4.scala 531:166 534:22]
  wire [31:0] _GEN_2979 = _T_712 == 32'h2 ? _i_vn_1_T_25 : _GEN_2977; // @[ivncontrol4.scala 531:166 535:22]
  wire [31:0] _GEN_2980 = _T_712 == 32'h3 ? _i_vn_1_T_25 : _GEN_2302; // @[ivncontrol4.scala 524:168 526:23]
  wire [31:0] _GEN_2981 = _T_712 == 32'h3 ? _i_vn_1_T_25 : _GEN_2978; // @[ivncontrol4.scala 524:168 527:22]
  wire [31:0] _GEN_2982 = _T_712 == 32'h3 ? _i_vn_1_T_25 : _GEN_2979; // @[ivncontrol4.scala 524:168 528:22]
  wire [31:0] _GEN_2983 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2301; // @[ivncontrol4.scala 518:166 520:22]
  wire [31:0] _GEN_2984 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2980; // @[ivncontrol4.scala 518:166 521:22]
  wire [31:0] _GEN_2985 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2981; // @[ivncontrol4.scala 518:166 522:22]
  wire [31:0] _GEN_2986 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2982; // @[ivncontrol4.scala 518:166 523:22]
  wire [31:0] _GEN_2987 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2300; // @[ivncontrol4.scala 511:166 513:23]
  wire [31:0] _GEN_2988 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2983; // @[ivncontrol4.scala 511:166 514:22]
  wire [31:0] _GEN_2989 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2984; // @[ivncontrol4.scala 511:166 515:22]
  wire [31:0] _GEN_2990 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2985; // @[ivncontrol4.scala 511:166 516:22]
  wire [31:0] _GEN_2991 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2986; // @[ivncontrol4.scala 511:166 517:22]
  wire [31:0] _GEN_2992 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2299; // @[ivncontrol4.scala 503:166 505:22]
  wire [31:0] _GEN_2993 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2987; // @[ivncontrol4.scala 503:166 506:21]
  wire [31:0] _GEN_2994 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2988; // @[ivncontrol4.scala 503:166 507:22]
  wire [31:0] _GEN_2995 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2989; // @[ivncontrol4.scala 503:166 508:22]
  wire [31:0] _GEN_2996 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2990; // @[ivncontrol4.scala 503:166 509:22]
  wire [31:0] _GEN_2997 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2991; // @[ivncontrol4.scala 503:166 510:22]
  wire [31:0] _GEN_2998 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2298; // @[ivncontrol4.scala 494:162 495:22]
  wire [31:0] _GEN_2999 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2992; // @[ivncontrol4.scala 494:162 496:21]
  wire [31:0] _GEN_3000 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2993; // @[ivncontrol4.scala 494:162 497:21]
  wire [31:0] _GEN_3001 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2994; // @[ivncontrol4.scala 494:162 498:22]
  wire [31:0] _GEN_3002 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2995; // @[ivncontrol4.scala 494:162 499:22]
  wire [31:0] _GEN_3003 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2996; // @[ivncontrol4.scala 494:162 500:22]
  wire [31:0] _GEN_3004 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2997; // @[ivncontrol4.scala 494:162 501:22]
  wire [31:0] _GEN_3102 = 4'h1 == _i_vn_1_T_25[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3103 = 4'h2 == _i_vn_1_T_25[3:0] ? rowcount_2 : _GEN_3102; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3104 = 4'h3 == _i_vn_1_T_25[3:0] ? rowcount_3 : _GEN_3103; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3105 = 4'h4 == _i_vn_1_T_25[3:0] ? rowcount_4 : _GEN_3104; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3106 = 4'h5 == _i_vn_1_T_25[3:0] ? rowcount_5 : _GEN_3105; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3107 = 4'h6 == _i_vn_1_T_25[3:0] ? rowcount_6 : _GEN_3106; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3108 = 4'h7 == _i_vn_1_T_25[3:0] ? rowcount_7 : _GEN_3107; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3109 = 4'h8 == _i_vn_1_T_25[3:0] ? rowcount_8 : _GEN_3108; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3110 = 4'h9 == _i_vn_1_T_25[3:0] ? rowcount_9 : _GEN_3109; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3111 = 4'ha == _i_vn_1_T_25[3:0] ? rowcount_10 : _GEN_3110; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3112 = 4'hb == _i_vn_1_T_25[3:0] ? rowcount_11 : _GEN_3111; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3113 = 4'hc == _i_vn_1_T_25[3:0] ? rowcount_12 : _GEN_3112; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3114 = 4'hd == _i_vn_1_T_25[3:0] ? rowcount_13 : _GEN_3113; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3115 = 4'he == _i_vn_1_T_25[3:0] ? rowcount_14 : _GEN_3114; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3116 = 4'hf == _i_vn_1_T_25[3:0] ? rowcount_15 : _GEN_3115; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _T_932 = _T_710 + _GEN_3116; // @[ivncontrol4.scala 545:152]
  wire [31:0] _T_934 = 32'h8 - _T_932; // @[ivncontrol4.scala 545:19]
  wire [31:0] _i_vn_1_T_27 = 32'h7 + pin; // @[ivncontrol4.scala 546:29]
  wire [31:0] _GEN_3789 = _T_934 == 32'h1 ? _i_vn_1_T_27 : _GEN_3004; // @[ivncontrol4.scala 588:188 591:22]
  wire [31:0] _GEN_3790 = _T_934 == 32'h2 ? _i_vn_1_T_27 : _GEN_3003; // @[ivncontrol4.scala 582:188 585:22]
  wire [31:0] _GEN_3791 = _T_934 == 32'h2 ? _i_vn_1_T_27 : _GEN_3789; // @[ivncontrol4.scala 582:188 586:22]
  wire [31:0] _GEN_3792 = _T_934 == 32'h3 ? _i_vn_1_T_27 : _GEN_3002; // @[ivncontrol4.scala 575:190 577:23]
  wire [31:0] _GEN_3793 = _T_934 == 32'h3 ? _i_vn_1_T_27 : _GEN_3790; // @[ivncontrol4.scala 575:190 578:22]
  wire [31:0] _GEN_3794 = _T_934 == 32'h3 ? _i_vn_1_T_27 : _GEN_3791; // @[ivncontrol4.scala 575:190 579:22]
  wire [31:0] _GEN_3795 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_3001; // @[ivncontrol4.scala 569:188 571:22]
  wire [31:0] _GEN_3796 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_3792; // @[ivncontrol4.scala 569:188 572:22]
  wire [31:0] _GEN_3797 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_3793; // @[ivncontrol4.scala 569:188 573:22]
  wire [31:0] _GEN_3798 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_3794; // @[ivncontrol4.scala 569:188 574:22]
  wire [31:0] _GEN_3799 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3000; // @[ivncontrol4.scala 562:188 564:23]
  wire [31:0] _GEN_3800 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3795; // @[ivncontrol4.scala 562:188 565:22]
  wire [31:0] _GEN_3801 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3796; // @[ivncontrol4.scala 562:188 566:22]
  wire [31:0] _GEN_3802 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3797; // @[ivncontrol4.scala 562:188 567:22]
  wire [31:0] _GEN_3803 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3798; // @[ivncontrol4.scala 562:188 568:22]
  wire [31:0] _GEN_3804 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_2999; // @[ivncontrol4.scala 554:188 556:22]
  wire [31:0] _GEN_3805 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3799; // @[ivncontrol4.scala 554:188 557:21]
  wire [31:0] _GEN_3806 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3800; // @[ivncontrol4.scala 554:188 558:22]
  wire [31:0] _GEN_3807 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3801; // @[ivncontrol4.scala 554:188 559:22]
  wire [31:0] _GEN_3808 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3802; // @[ivncontrol4.scala 554:188 560:22]
  wire [31:0] _GEN_3809 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3803; // @[ivncontrol4.scala 554:188 561:22]
  wire [31:0] _GEN_3810 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_2998; // @[ivncontrol4.scala 545:184 546:22]
  wire [31:0] _GEN_3811 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3804; // @[ivncontrol4.scala 545:184 547:21]
  wire [31:0] _GEN_3812 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3805; // @[ivncontrol4.scala 545:184 548:21]
  wire [31:0] _GEN_3813 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3806; // @[ivncontrol4.scala 545:184 549:22]
  wire [31:0] _GEN_3814 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3807; // @[ivncontrol4.scala 545:184 550:22]
  wire [31:0] _GEN_3815 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3808; // @[ivncontrol4.scala 545:184 551:22]
  wire [31:0] _GEN_3816 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3809; // @[ivncontrol4.scala 545:184 552:22]
  wire [31:0] _GEN_3817 = _GEN_312 ? _GEN_477 : 32'h19; // @[ivncontrol4.scala 142:17 189:28]
  wire [31:0] _GEN_3818 = _GEN_312 ? _GEN_3810 : 32'h3; // @[ivncontrol4.scala 142:17 189:28]
  wire [31:0] _GEN_3819 = _GEN_312 ? _GEN_3811 : 32'h1c; // @[ivncontrol4.scala 142:17 189:28]
  wire [31:0] _GEN_3820 = _GEN_312 ? _GEN_3812 : 32'h4; // @[ivncontrol4.scala 142:17 189:28]
  wire [31:0] _GEN_3821 = _GEN_312 ? _GEN_3813 : 32'h14; // @[ivncontrol4.scala 143:18 189:28]
  wire [31:0] _GEN_3822 = _GEN_312 ? _GEN_3814 : 32'h1b; // @[ivncontrol4.scala 143:18 189:28]
  wire [31:0] _GEN_3823 = _GEN_312 ? _GEN_3815 : 32'h5; // @[ivncontrol4.scala 143:18 189:28]
  wire [31:0] _GEN_3824 = _GEN_312 ? _GEN_3816 : 32'h8; // @[ivncontrol4.scala 143:18 189:28]
  wire  valid1 = 1'h0;
  wire [31:0] _GEN_4221 = reset ? 32'h0 : _GEN_3817; // @[ivncontrol4.scala 17:{23,23}]
  wire [31:0] _GEN_4222 = reset ? 32'h0 : _GEN_3818; // @[ivncontrol4.scala 17:{23,23}]
  wire [31:0] _GEN_4223 = reset ? 32'h0 : _GEN_3819; // @[ivncontrol4.scala 17:{23,23}]
  wire [31:0] _GEN_4224 = reset ? 32'h0 : _GEN_3820; // @[ivncontrol4.scala 17:{23,23}]
  wire [31:0] _GEN_4225 = reset ? 32'h0 : _GEN_3821; // @[ivncontrol4.scala 18:{24,24}]
  wire [31:0] _GEN_4226 = reset ? 32'h0 : _GEN_3822; // @[ivncontrol4.scala 18:{24,24}]
  wire [31:0] _GEN_4227 = reset ? 32'h0 : _GEN_3823; // @[ivncontrol4.scala 18:{24,24}]
  wire [31:0] _GEN_4228 = reset ? 32'h0 : _GEN_3824; // @[ivncontrol4.scala 18:{24,24}]
  assign io_o_vn_0 = i_vn_0; // @[ivncontrol4.scala 138:13]
  assign io_o_vn_1 = i_vn_1; // @[ivncontrol4.scala 138:13]
  assign io_o_vn_2 = i_vn_2; // @[ivncontrol4.scala 138:13]
  assign io_o_vn_3 = i_vn_3; // @[ivncontrol4.scala 138:13]
  assign io_o_vn2_0 = i_vn2_0; // @[ivncontrol4.scala 139:14]
  assign io_o_vn2_1 = i_vn2_1; // @[ivncontrol4.scala 139:14]
  assign io_o_vn2_2 = i_vn2_2; // @[ivncontrol4.scala 139:14]
  assign io_o_vn2_3 = i_vn2_3; // @[ivncontrol4.scala 139:14]
  always @(posedge clock) begin
    i_vn_0 <= _GEN_4221[4:0]; // @[ivncontrol4.scala 17:{23,23}]
    i_vn_1 <= _GEN_4222[4:0]; // @[ivncontrol4.scala 17:{23,23}]
    i_vn_2 <= _GEN_4223[4:0]; // @[ivncontrol4.scala 17:{23,23}]
    i_vn_3 <= _GEN_4224[4:0]; // @[ivncontrol4.scala 17:{23,23}]
    i_vn2_0 <= _GEN_4225[4:0]; // @[ivncontrol4.scala 18:{24,24}]
    i_vn2_1 <= _GEN_4226[4:0]; // @[ivncontrol4.scala 18:{24,24}]
    i_vn2_2 <= _GEN_4227[4:0]; // @[ivncontrol4.scala 18:{24,24}]
    i_vn2_3 <= _GEN_4228[4:0]; // @[ivncontrol4.scala 18:{24,24}]
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_0 <= io_Stationary_matrix_0_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_1 <= io_Stationary_matrix_0_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_2 <= io_Stationary_matrix_0_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_3 <= io_Stationary_matrix_0_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_4 <= io_Stationary_matrix_0_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_5 <= io_Stationary_matrix_0_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_6 <= io_Stationary_matrix_0_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_7 <= io_Stationary_matrix_0_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_0 <= io_Stationary_matrix_1_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_1 <= io_Stationary_matrix_1_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_2 <= io_Stationary_matrix_1_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_3 <= io_Stationary_matrix_1_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_4 <= io_Stationary_matrix_1_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_5 <= io_Stationary_matrix_1_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_6 <= io_Stationary_matrix_1_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_7 <= io_Stationary_matrix_1_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_0 <= io_Stationary_matrix_2_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_1 <= io_Stationary_matrix_2_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_2 <= io_Stationary_matrix_2_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_3 <= io_Stationary_matrix_2_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_4 <= io_Stationary_matrix_2_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_5 <= io_Stationary_matrix_2_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_6 <= io_Stationary_matrix_2_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_7 <= io_Stationary_matrix_2_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_0 <= io_Stationary_matrix_3_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_1 <= io_Stationary_matrix_3_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_2 <= io_Stationary_matrix_3_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_3 <= io_Stationary_matrix_3_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_4 <= io_Stationary_matrix_3_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_5 <= io_Stationary_matrix_3_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_6 <= io_Stationary_matrix_3_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_7 <= io_Stationary_matrix_3_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_0 <= io_Stationary_matrix_4_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_1 <= io_Stationary_matrix_4_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_2 <= io_Stationary_matrix_4_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_3 <= io_Stationary_matrix_4_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_4 <= io_Stationary_matrix_4_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_5 <= io_Stationary_matrix_4_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_6 <= io_Stationary_matrix_4_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_7 <= io_Stationary_matrix_4_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_0 <= io_Stationary_matrix_5_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_1 <= io_Stationary_matrix_5_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_2 <= io_Stationary_matrix_5_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_3 <= io_Stationary_matrix_5_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_4 <= io_Stationary_matrix_5_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_5 <= io_Stationary_matrix_5_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_6 <= io_Stationary_matrix_5_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_7 <= io_Stationary_matrix_5_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_0 <= io_Stationary_matrix_6_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_1 <= io_Stationary_matrix_6_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_2 <= io_Stationary_matrix_6_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_3 <= io_Stationary_matrix_6_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_4 <= io_Stationary_matrix_6_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_5 <= io_Stationary_matrix_6_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_6 <= io_Stationary_matrix_6_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_7 <= io_Stationary_matrix_6_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_0 <= io_Stationary_matrix_7_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_1 <= io_Stationary_matrix_7_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_2 <= io_Stationary_matrix_7_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_3 <= io_Stationary_matrix_7_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_4 <= io_Stationary_matrix_7_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_5 <= io_Stationary_matrix_7_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_6 <= io_Stationary_matrix_7_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_7 <= io_Stationary_matrix_7_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_0 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_0 <= count_0; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_1 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_1 <= count_1; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_2 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_2 <= count_2; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_3 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_3 <= count_3; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_4 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_4 <= count_4; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_5 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_5 <= count_5; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_6 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_6 <= count_6; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_7 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_7 <= count_7; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_8 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_8 <= 32'h0; // @[ivncontrol4.scala 87:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_9 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_9 <= 32'h0; // @[ivncontrol4.scala 87:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_10 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_10 <= 32'h0; // @[ivncontrol4.scala 87:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_11 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_11 <= 32'h0; // @[ivncontrol4.scala 87:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_12 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_12 <= 32'h0; // @[ivncontrol4.scala 87:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_13 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_13 <= 32'h0; // @[ivncontrol4.scala 87:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_14 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_14 <= 32'h0; // @[ivncontrol4.scala 87:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_15 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end
    if (reset) begin // @[ivncontrol4.scala 37:22]
      pin <= 32'h0; // @[ivncontrol4.scala 37:22]
    end else if (_T_72 & rowcount_6 == 32'h0 & rowcount_7 != 32'h0) begin // @[ivncontrol4.scala 183:192]
      pin <= 32'h7; // @[ivncontrol4.scala 184:13]
    end else if (_T_59 & rowcount_5 == 32'h0 & rowcount_6 != 32'h0) begin // @[ivncontrol4.scala 180:169]
      pin <= 32'h6; // @[ivncontrol4.scala 181:13]
    end else if (_T_48 & rowcount_4 == 32'h0 & rowcount_5 != 32'h0) begin // @[ivncontrol4.scala 177:146]
      pin <= 32'h5; // @[ivncontrol4.scala 178:13]
    end else begin
      pin <= _GEN_317;
    end
    if (reset) begin // @[ivncontrol4.scala 41:20]
      i <= 32'h0; // @[ivncontrol4.scala 41:20]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
        i <= _GEN_247;
      end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
        i <= _GEN_247;
      end else begin
        i <= _GEN_265;
      end
    end
    if (reset) begin // @[ivncontrol4.scala 42:20]
      j <= 32'h0; // @[ivncontrol4.scala 42:20]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
        j <= 32'h8; // @[ivncontrol4.scala 116:11]
      end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
        j <= _j_T_1; // @[ivncontrol4.scala 118:11]
      end else begin
        j <= {{28'd0}, _GEN_264};
      end
    end
    if (3'h0 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h0 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h0 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h0 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h0 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h0 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h0 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h0 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_0 <= _GEN_224;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_0 <= _GEN_224;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h0 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_0 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_0 <= _GEN_224;
      end
    end else begin
      count_0 <= _GEN_224;
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_1 <= _GEN_225;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_1 <= _GEN_225;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h1 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_1 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_1 <= _GEN_225;
      end
    end else begin
      count_1 <= _GEN_225;
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_2 <= _GEN_226;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_2 <= _GEN_226;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h2 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_2 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_2 <= _GEN_226;
      end
    end else begin
      count_2 <= _GEN_226;
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_3 <= _GEN_227;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_3 <= _GEN_227;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h3 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_3 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_3 <= _GEN_227;
      end
    end else begin
      count_3 <= _GEN_227;
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_4 <= _GEN_228;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_4 <= _GEN_228;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h4 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_4 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_4 <= _GEN_228;
      end
    end else begin
      count_4 <= _GEN_228;
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_5 <= _GEN_229;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_5 <= _GEN_229;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h5 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_5 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_5 <= _GEN_229;
      end
    end else begin
      count_5 <= _GEN_229;
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_6 <= _GEN_230;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_6 <= _GEN_230;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h6 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_6 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_6 <= _GEN_230;
      end
    end else begin
      count_6 <= _GEN_230;
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_7 <= _GEN_231;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_7 <= _GEN_231;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h7 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_7 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_7 <= _GEN_231;
      end
    end else begin
      count_7 <= _GEN_231;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  i_vn_0 = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  i_vn_1 = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  i_vn_2 = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  i_vn_3 = _RAND_3[4:0];
  _RAND_4 = {1{`RANDOM}};
  i_vn2_0 = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  i_vn2_1 = _RAND_5[4:0];
  _RAND_6 = {1{`RANDOM}};
  i_vn2_2 = _RAND_6[4:0];
  _RAND_7 = {1{`RANDOM}};
  i_vn2_3 = _RAND_7[4:0];
  _RAND_8 = {1{`RANDOM}};
  solution_0_0 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  solution_0_1 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  solution_0_2 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  solution_0_3 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  solution_0_4 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  solution_0_5 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  solution_0_6 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  solution_0_7 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  solution_1_0 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  solution_1_1 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  solution_1_2 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  solution_1_3 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  solution_1_4 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  solution_1_5 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  solution_1_6 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  solution_1_7 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  solution_2_0 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  solution_2_1 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  solution_2_2 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  solution_2_3 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  solution_2_4 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  solution_2_5 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  solution_2_6 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  solution_2_7 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  solution_3_0 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  solution_3_1 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  solution_3_2 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  solution_3_3 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  solution_3_4 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  solution_3_5 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  solution_3_6 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  solution_3_7 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  solution_4_0 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  solution_4_1 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  solution_4_2 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  solution_4_3 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  solution_4_4 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  solution_4_5 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  solution_4_6 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  solution_4_7 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  solution_5_0 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  solution_5_1 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  solution_5_2 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  solution_5_3 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  solution_5_4 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  solution_5_5 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  solution_5_6 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  solution_5_7 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  solution_6_0 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  solution_6_1 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  solution_6_2 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  solution_6_3 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  solution_6_4 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  solution_6_5 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  solution_6_6 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  solution_6_7 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  solution_7_0 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  solution_7_1 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  solution_7_2 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  solution_7_3 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  solution_7_4 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  solution_7_5 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  solution_7_6 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  solution_7_7 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  rowcount_0 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  rowcount_1 = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  rowcount_2 = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  rowcount_3 = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  rowcount_4 = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  rowcount_5 = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  rowcount_6 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  rowcount_7 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  rowcount_8 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  rowcount_9 = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  rowcount_10 = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  rowcount_11 = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  rowcount_12 = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  rowcount_13 = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  rowcount_14 = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  rowcount_15 = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  pin = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  i = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  j = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  mat_0_0 = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  mat_0_1 = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  mat_0_2 = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  mat_0_3 = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  mat_0_4 = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  mat_0_5 = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  mat_0_6 = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  mat_0_7 = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  mat_1_0 = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  mat_1_1 = _RAND_100[31:0];
  _RAND_101 = {1{`RANDOM}};
  mat_1_2 = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  mat_1_3 = _RAND_102[31:0];
  _RAND_103 = {1{`RANDOM}};
  mat_1_4 = _RAND_103[31:0];
  _RAND_104 = {1{`RANDOM}};
  mat_1_5 = _RAND_104[31:0];
  _RAND_105 = {1{`RANDOM}};
  mat_1_6 = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  mat_1_7 = _RAND_106[31:0];
  _RAND_107 = {1{`RANDOM}};
  mat_2_0 = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  mat_2_1 = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  mat_2_2 = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  mat_2_3 = _RAND_110[31:0];
  _RAND_111 = {1{`RANDOM}};
  mat_2_4 = _RAND_111[31:0];
  _RAND_112 = {1{`RANDOM}};
  mat_2_5 = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  mat_2_6 = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  mat_2_7 = _RAND_114[31:0];
  _RAND_115 = {1{`RANDOM}};
  mat_3_0 = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  mat_3_1 = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  mat_3_2 = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  mat_3_3 = _RAND_118[31:0];
  _RAND_119 = {1{`RANDOM}};
  mat_3_4 = _RAND_119[31:0];
  _RAND_120 = {1{`RANDOM}};
  mat_3_5 = _RAND_120[31:0];
  _RAND_121 = {1{`RANDOM}};
  mat_3_6 = _RAND_121[31:0];
  _RAND_122 = {1{`RANDOM}};
  mat_3_7 = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  mat_4_0 = _RAND_123[31:0];
  _RAND_124 = {1{`RANDOM}};
  mat_4_1 = _RAND_124[31:0];
  _RAND_125 = {1{`RANDOM}};
  mat_4_2 = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  mat_4_3 = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  mat_4_4 = _RAND_127[31:0];
  _RAND_128 = {1{`RANDOM}};
  mat_4_5 = _RAND_128[31:0];
  _RAND_129 = {1{`RANDOM}};
  mat_4_6 = _RAND_129[31:0];
  _RAND_130 = {1{`RANDOM}};
  mat_4_7 = _RAND_130[31:0];
  _RAND_131 = {1{`RANDOM}};
  mat_5_0 = _RAND_131[31:0];
  _RAND_132 = {1{`RANDOM}};
  mat_5_1 = _RAND_132[31:0];
  _RAND_133 = {1{`RANDOM}};
  mat_5_2 = _RAND_133[31:0];
  _RAND_134 = {1{`RANDOM}};
  mat_5_3 = _RAND_134[31:0];
  _RAND_135 = {1{`RANDOM}};
  mat_5_4 = _RAND_135[31:0];
  _RAND_136 = {1{`RANDOM}};
  mat_5_5 = _RAND_136[31:0];
  _RAND_137 = {1{`RANDOM}};
  mat_5_6 = _RAND_137[31:0];
  _RAND_138 = {1{`RANDOM}};
  mat_5_7 = _RAND_138[31:0];
  _RAND_139 = {1{`RANDOM}};
  mat_6_0 = _RAND_139[31:0];
  _RAND_140 = {1{`RANDOM}};
  mat_6_1 = _RAND_140[31:0];
  _RAND_141 = {1{`RANDOM}};
  mat_6_2 = _RAND_141[31:0];
  _RAND_142 = {1{`RANDOM}};
  mat_6_3 = _RAND_142[31:0];
  _RAND_143 = {1{`RANDOM}};
  mat_6_4 = _RAND_143[31:0];
  _RAND_144 = {1{`RANDOM}};
  mat_6_5 = _RAND_144[31:0];
  _RAND_145 = {1{`RANDOM}};
  mat_6_6 = _RAND_145[31:0];
  _RAND_146 = {1{`RANDOM}};
  mat_6_7 = _RAND_146[31:0];
  _RAND_147 = {1{`RANDOM}};
  mat_7_0 = _RAND_147[31:0];
  _RAND_148 = {1{`RANDOM}};
  mat_7_1 = _RAND_148[31:0];
  _RAND_149 = {1{`RANDOM}};
  mat_7_2 = _RAND_149[31:0];
  _RAND_150 = {1{`RANDOM}};
  mat_7_3 = _RAND_150[31:0];
  _RAND_151 = {1{`RANDOM}};
  mat_7_4 = _RAND_151[31:0];
  _RAND_152 = {1{`RANDOM}};
  mat_7_5 = _RAND_152[31:0];
  _RAND_153 = {1{`RANDOM}};
  mat_7_6 = _RAND_153[31:0];
  _RAND_154 = {1{`RANDOM}};
  mat_7_7 = _RAND_154[31:0];
  _RAND_155 = {1{`RANDOM}};
  count_0 = _RAND_155[31:0];
  _RAND_156 = {1{`RANDOM}};
  count_1 = _RAND_156[31:0];
  _RAND_157 = {1{`RANDOM}};
  count_2 = _RAND_157[31:0];
  _RAND_158 = {1{`RANDOM}};
  count_3 = _RAND_158[31:0];
  _RAND_159 = {1{`RANDOM}};
  count_4 = _RAND_159[31:0];
  _RAND_160 = {1{`RANDOM}};
  count_5 = _RAND_160[31:0];
  _RAND_161 = {1{`RANDOM}};
  count_6 = _RAND_161[31:0];
  _RAND_162 = {1{`RANDOM}};
  count_7 = _RAND_162[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ivncontrol4_3(
  input         clock,
  input         reset,
  input  [15:0] io_Stationary_matrix_0_0,
  input  [15:0] io_Stationary_matrix_0_1,
  input  [15:0] io_Stationary_matrix_0_2,
  input  [15:0] io_Stationary_matrix_0_3,
  input  [15:0] io_Stationary_matrix_0_4,
  input  [15:0] io_Stationary_matrix_0_5,
  input  [15:0] io_Stationary_matrix_0_6,
  input  [15:0] io_Stationary_matrix_0_7,
  input  [15:0] io_Stationary_matrix_1_0,
  input  [15:0] io_Stationary_matrix_1_1,
  input  [15:0] io_Stationary_matrix_1_2,
  input  [15:0] io_Stationary_matrix_1_3,
  input  [15:0] io_Stationary_matrix_1_4,
  input  [15:0] io_Stationary_matrix_1_5,
  input  [15:0] io_Stationary_matrix_1_6,
  input  [15:0] io_Stationary_matrix_1_7,
  input  [15:0] io_Stationary_matrix_2_0,
  input  [15:0] io_Stationary_matrix_2_1,
  input  [15:0] io_Stationary_matrix_2_2,
  input  [15:0] io_Stationary_matrix_2_3,
  input  [15:0] io_Stationary_matrix_2_4,
  input  [15:0] io_Stationary_matrix_2_5,
  input  [15:0] io_Stationary_matrix_2_6,
  input  [15:0] io_Stationary_matrix_2_7,
  input  [15:0] io_Stationary_matrix_3_0,
  input  [15:0] io_Stationary_matrix_3_1,
  input  [15:0] io_Stationary_matrix_3_2,
  input  [15:0] io_Stationary_matrix_3_3,
  input  [15:0] io_Stationary_matrix_3_4,
  input  [15:0] io_Stationary_matrix_3_5,
  input  [15:0] io_Stationary_matrix_3_6,
  input  [15:0] io_Stationary_matrix_3_7,
  input  [15:0] io_Stationary_matrix_4_0,
  input  [15:0] io_Stationary_matrix_4_1,
  input  [15:0] io_Stationary_matrix_4_2,
  input  [15:0] io_Stationary_matrix_4_3,
  input  [15:0] io_Stationary_matrix_4_4,
  input  [15:0] io_Stationary_matrix_4_5,
  input  [15:0] io_Stationary_matrix_4_6,
  input  [15:0] io_Stationary_matrix_4_7,
  input  [15:0] io_Stationary_matrix_5_0,
  input  [15:0] io_Stationary_matrix_5_1,
  input  [15:0] io_Stationary_matrix_5_2,
  input  [15:0] io_Stationary_matrix_5_3,
  input  [15:0] io_Stationary_matrix_5_4,
  input  [15:0] io_Stationary_matrix_5_5,
  input  [15:0] io_Stationary_matrix_5_6,
  input  [15:0] io_Stationary_matrix_5_7,
  input  [15:0] io_Stationary_matrix_6_0,
  input  [15:0] io_Stationary_matrix_6_1,
  input  [15:0] io_Stationary_matrix_6_2,
  input  [15:0] io_Stationary_matrix_6_3,
  input  [15:0] io_Stationary_matrix_6_4,
  input  [15:0] io_Stationary_matrix_6_5,
  input  [15:0] io_Stationary_matrix_6_6,
  input  [15:0] io_Stationary_matrix_6_7,
  input  [15:0] io_Stationary_matrix_7_0,
  input  [15:0] io_Stationary_matrix_7_1,
  input  [15:0] io_Stationary_matrix_7_2,
  input  [15:0] io_Stationary_matrix_7_3,
  input  [15:0] io_Stationary_matrix_7_4,
  input  [15:0] io_Stationary_matrix_7_5,
  input  [15:0] io_Stationary_matrix_7_6,
  input  [15:0] io_Stationary_matrix_7_7,
  output [4:0]  io_o_vn_0,
  output [4:0]  io_o_vn_1,
  output [4:0]  io_o_vn_2,
  output [4:0]  io_o_vn_3,
  output [4:0]  io_o_vn2_0,
  output [4:0]  io_o_vn2_1,
  output [4:0]  io_o_vn2_2,
  output [4:0]  io_o_vn2_3,
  input         io_validpin
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
`endif // RANDOMIZE_REG_INIT
  reg [4:0] i_vn_0; // @[ivncontrol4.scala 17:23]
  reg [4:0] i_vn_1; // @[ivncontrol4.scala 17:23]
  reg [4:0] i_vn_2; // @[ivncontrol4.scala 17:23]
  reg [4:0] i_vn_3; // @[ivncontrol4.scala 17:23]
  reg [4:0] i_vn2_0; // @[ivncontrol4.scala 18:24]
  reg [4:0] i_vn2_1; // @[ivncontrol4.scala 18:24]
  reg [4:0] i_vn2_2; // @[ivncontrol4.scala 18:24]
  reg [4:0] i_vn2_3; // @[ivncontrol4.scala 18:24]
  reg [15:0] solution_0_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_0_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_0_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_0_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_0_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_0_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_0_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_0_7; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_7; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_7; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_7; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_7; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_7; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_7; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_7; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_0; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_1; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_2; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_3; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_4; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_5; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_6; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_7; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_8; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_9; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_10; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_11; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_12; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_13; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_14; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_15; // @[ivncontrol4.scala 27:27]
  reg [31:0] pin; // @[ivncontrol4.scala 37:22]
  reg [31:0] i; // @[ivncontrol4.scala 41:20]
  reg [31:0] j; // @[ivncontrol4.scala 42:20]
  wire  _io_ProcessValid_T = i == 32'h7; // @[ivncontrol4.scala 44:27]
  wire  _io_ProcessValid_T_1 = j == 32'h7; // @[ivncontrol4.scala 44:42]
  wire  _io_ProcessValid_T_2 = i == 32'h7 & j == 32'h7; // @[ivncontrol4.scala 44:36]
  reg [31:0] mat_0_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_0_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_0_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_0_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_0_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_0_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_0_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_0_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] count_0; // @[ivncontrol4.scala 58:20]
  reg [31:0] count_1; // @[ivncontrol4.scala 58:20]
  reg [31:0] count_2; // @[ivncontrol4.scala 58:20]
  reg [31:0] count_3; // @[ivncontrol4.scala 58:20]
  reg [31:0] count_4; // @[ivncontrol4.scala 58:20]
  reg [31:0] count_5; // @[ivncontrol4.scala 58:20]
  reg [31:0] count_6; // @[ivncontrol4.scala 58:20]
  reg [31:0] count_7; // @[ivncontrol4.scala 58:20]
  wire  _GEN_3825 = 3'h0 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_65 = 3'h0 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_0_1 : io_Stationary_matrix_0_0; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_66 = 3'h0 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_0_2 : _GEN_65; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_67 = 3'h0 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_0_3 : _GEN_66; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_68 = 3'h0 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_0_4 : _GEN_67; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_69 = 3'h0 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_0_5 : _GEN_68; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_70 = 3'h0 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_0_6 : _GEN_69; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_71 = 3'h0 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_0_7 : _GEN_70; // @[ivncontrol4.scala 63:{17,17}]
  wire  _GEN_3839 = 3'h1 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_72 = 3'h1 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_1_0 : _GEN_71; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_73 = 3'h1 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_1_1 : _GEN_72; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_74 = 3'h1 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_1_2 : _GEN_73; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_75 = 3'h1 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_1_3 : _GEN_74; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_76 = 3'h1 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_1_4 : _GEN_75; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_77 = 3'h1 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_1_5 : _GEN_76; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_78 = 3'h1 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_1_6 : _GEN_77; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_79 = 3'h1 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_1_7 : _GEN_78; // @[ivncontrol4.scala 63:{17,17}]
  wire  _GEN_3855 = 3'h2 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_80 = 3'h2 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_2_0 : _GEN_79; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_81 = 3'h2 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_2_1 : _GEN_80; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_82 = 3'h2 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_2_2 : _GEN_81; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_83 = 3'h2 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_2_3 : _GEN_82; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_84 = 3'h2 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_2_4 : _GEN_83; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_85 = 3'h2 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_2_5 : _GEN_84; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_86 = 3'h2 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_2_6 : _GEN_85; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_87 = 3'h2 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_2_7 : _GEN_86; // @[ivncontrol4.scala 63:{17,17}]
  wire  _GEN_3871 = 3'h3 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_88 = 3'h3 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_3_0 : _GEN_87; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_89 = 3'h3 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_3_1 : _GEN_88; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_90 = 3'h3 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_3_2 : _GEN_89; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_91 = 3'h3 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_3_3 : _GEN_90; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_92 = 3'h3 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_3_4 : _GEN_91; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_93 = 3'h3 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_3_5 : _GEN_92; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_94 = 3'h3 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_3_6 : _GEN_93; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_95 = 3'h3 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_3_7 : _GEN_94; // @[ivncontrol4.scala 63:{17,17}]
  wire  _GEN_3887 = 3'h4 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_96 = 3'h4 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_4_0 : _GEN_95; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_97 = 3'h4 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_4_1 : _GEN_96; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_98 = 3'h4 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_4_2 : _GEN_97; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_99 = 3'h4 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_4_3 : _GEN_98; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_100 = 3'h4 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_4_4 : _GEN_99; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_101 = 3'h4 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_4_5 : _GEN_100; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_102 = 3'h4 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_4_6 : _GEN_101; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_103 = 3'h4 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_4_7 : _GEN_102; // @[ivncontrol4.scala 63:{17,17}]
  wire  _GEN_3903 = 3'h5 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_104 = 3'h5 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_5_0 : _GEN_103; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_105 = 3'h5 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_5_1 : _GEN_104; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_106 = 3'h5 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_5_2 : _GEN_105; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_107 = 3'h5 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_5_3 : _GEN_106; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_108 = 3'h5 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_5_4 : _GEN_107; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_109 = 3'h5 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_5_5 : _GEN_108; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_110 = 3'h5 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_5_6 : _GEN_109; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_111 = 3'h5 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_5_7 : _GEN_110; // @[ivncontrol4.scala 63:{17,17}]
  wire  _GEN_3919 = 3'h6 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_112 = 3'h6 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_6_0 : _GEN_111; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_113 = 3'h6 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_6_1 : _GEN_112; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_114 = 3'h6 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_6_2 : _GEN_113; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_115 = 3'h6 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_6_3 : _GEN_114; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_116 = 3'h6 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_6_4 : _GEN_115; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_117 = 3'h6 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_6_5 : _GEN_116; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_118 = 3'h6 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_6_6 : _GEN_117; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_119 = 3'h6 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_6_7 : _GEN_118; // @[ivncontrol4.scala 63:{17,17}]
  wire  _GEN_3935 = 3'h7 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_120 = 3'h7 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_7_0 : _GEN_119; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_121 = 3'h7 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_7_1 : _GEN_120; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_122 = 3'h7 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_7_2 : _GEN_121; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_123 = 3'h7 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_7_3 : _GEN_122; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_124 = 3'h7 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_7_4 : _GEN_123; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_125 = 3'h7 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_7_5 : _GEN_124; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_126 = 3'h7 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_7_6 : _GEN_125; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_127 = 3'h7 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_7_7 : _GEN_126; // @[ivncontrol4.scala 63:{17,17}]
  wire [31:0] _mat_T_1_T_2 = {{16'd0}, _GEN_127}; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_129 = _GEN_3825 & 4'h1 == j[3:0] ? solution_0_1 : solution_0_0; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_130 = _GEN_3825 & 4'h2 == j[3:0] ? solution_0_2 : _GEN_129; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_131 = _GEN_3825 & 4'h3 == j[3:0] ? solution_0_3 : _GEN_130; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_132 = _GEN_3825 & 4'h4 == j[3:0] ? solution_0_4 : _GEN_131; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_133 = _GEN_3825 & 4'h5 == j[3:0] ? solution_0_5 : _GEN_132; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_134 = _GEN_3825 & 4'h6 == j[3:0] ? solution_0_6 : _GEN_133; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_135 = _GEN_3825 & 4'h7 == j[3:0] ? solution_0_7 : _GEN_134; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_136 = _GEN_3825 & 4'h8 == j[3:0] ? 16'h0 : _GEN_135; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_137 = _GEN_3839 & 4'h0 == j[3:0] ? solution_1_0 : _GEN_136; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_138 = _GEN_3839 & 4'h1 == j[3:0] ? solution_1_1 : _GEN_137; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_139 = _GEN_3839 & 4'h2 == j[3:0] ? solution_1_2 : _GEN_138; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_140 = _GEN_3839 & 4'h3 == j[3:0] ? solution_1_3 : _GEN_139; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_141 = _GEN_3839 & 4'h4 == j[3:0] ? solution_1_4 : _GEN_140; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_142 = _GEN_3839 & 4'h5 == j[3:0] ? solution_1_5 : _GEN_141; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_143 = _GEN_3839 & 4'h6 == j[3:0] ? solution_1_6 : _GEN_142; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_144 = _GEN_3839 & 4'h7 == j[3:0] ? solution_1_7 : _GEN_143; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_145 = _GEN_3839 & 4'h8 == j[3:0] ? 16'h0 : _GEN_144; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_146 = _GEN_3855 & 4'h0 == j[3:0] ? solution_2_0 : _GEN_145; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_147 = _GEN_3855 & 4'h1 == j[3:0] ? solution_2_1 : _GEN_146; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_148 = _GEN_3855 & 4'h2 == j[3:0] ? solution_2_2 : _GEN_147; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_149 = _GEN_3855 & 4'h3 == j[3:0] ? solution_2_3 : _GEN_148; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_150 = _GEN_3855 & 4'h4 == j[3:0] ? solution_2_4 : _GEN_149; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_151 = _GEN_3855 & 4'h5 == j[3:0] ? solution_2_5 : _GEN_150; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_152 = _GEN_3855 & 4'h6 == j[3:0] ? solution_2_6 : _GEN_151; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_153 = _GEN_3855 & 4'h7 == j[3:0] ? solution_2_7 : _GEN_152; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_154 = _GEN_3855 & 4'h8 == j[3:0] ? 16'h0 : _GEN_153; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_155 = _GEN_3871 & 4'h0 == j[3:0] ? solution_3_0 : _GEN_154; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_156 = _GEN_3871 & 4'h1 == j[3:0] ? solution_3_1 : _GEN_155; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_157 = _GEN_3871 & 4'h2 == j[3:0] ? solution_3_2 : _GEN_156; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_158 = _GEN_3871 & 4'h3 == j[3:0] ? solution_3_3 : _GEN_157; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_159 = _GEN_3871 & 4'h4 == j[3:0] ? solution_3_4 : _GEN_158; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_160 = _GEN_3871 & 4'h5 == j[3:0] ? solution_3_5 : _GEN_159; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_161 = _GEN_3871 & 4'h6 == j[3:0] ? solution_3_6 : _GEN_160; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_162 = _GEN_3871 & 4'h7 == j[3:0] ? solution_3_7 : _GEN_161; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_163 = _GEN_3871 & 4'h8 == j[3:0] ? 16'h0 : _GEN_162; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_164 = _GEN_3887 & 4'h0 == j[3:0] ? solution_4_0 : _GEN_163; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_165 = _GEN_3887 & 4'h1 == j[3:0] ? solution_4_1 : _GEN_164; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_166 = _GEN_3887 & 4'h2 == j[3:0] ? solution_4_2 : _GEN_165; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_167 = _GEN_3887 & 4'h3 == j[3:0] ? solution_4_3 : _GEN_166; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_168 = _GEN_3887 & 4'h4 == j[3:0] ? solution_4_4 : _GEN_167; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_169 = _GEN_3887 & 4'h5 == j[3:0] ? solution_4_5 : _GEN_168; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_170 = _GEN_3887 & 4'h6 == j[3:0] ? solution_4_6 : _GEN_169; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_171 = _GEN_3887 & 4'h7 == j[3:0] ? solution_4_7 : _GEN_170; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_172 = _GEN_3887 & 4'h8 == j[3:0] ? 16'h0 : _GEN_171; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_173 = _GEN_3903 & 4'h0 == j[3:0] ? solution_5_0 : _GEN_172; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_174 = _GEN_3903 & 4'h1 == j[3:0] ? solution_5_1 : _GEN_173; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_175 = _GEN_3903 & 4'h2 == j[3:0] ? solution_5_2 : _GEN_174; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_176 = _GEN_3903 & 4'h3 == j[3:0] ? solution_5_3 : _GEN_175; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_177 = _GEN_3903 & 4'h4 == j[3:0] ? solution_5_4 : _GEN_176; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_178 = _GEN_3903 & 4'h5 == j[3:0] ? solution_5_5 : _GEN_177; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_179 = _GEN_3903 & 4'h6 == j[3:0] ? solution_5_6 : _GEN_178; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_180 = _GEN_3903 & 4'h7 == j[3:0] ? solution_5_7 : _GEN_179; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_181 = _GEN_3903 & 4'h8 == j[3:0] ? 16'h0 : _GEN_180; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_182 = _GEN_3919 & 4'h0 == j[3:0] ? solution_6_0 : _GEN_181; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_183 = _GEN_3919 & 4'h1 == j[3:0] ? solution_6_1 : _GEN_182; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_184 = _GEN_3919 & 4'h2 == j[3:0] ? solution_6_2 : _GEN_183; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_185 = _GEN_3919 & 4'h3 == j[3:0] ? solution_6_3 : _GEN_184; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_186 = _GEN_3919 & 4'h4 == j[3:0] ? solution_6_4 : _GEN_185; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_187 = _GEN_3919 & 4'h5 == j[3:0] ? solution_6_5 : _GEN_186; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_188 = _GEN_3919 & 4'h6 == j[3:0] ? solution_6_6 : _GEN_187; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_189 = _GEN_3919 & 4'h7 == j[3:0] ? solution_6_7 : _GEN_188; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_190 = _GEN_3919 & 4'h8 == j[3:0] ? 16'h0 : _GEN_189; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_191 = _GEN_3935 & 4'h0 == j[3:0] ? solution_7_0 : _GEN_190; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_192 = _GEN_3935 & 4'h1 == j[3:0] ? solution_7_1 : _GEN_191; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_193 = _GEN_3935 & 4'h2 == j[3:0] ? solution_7_2 : _GEN_192; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_194 = _GEN_3935 & 4'h3 == j[3:0] ? solution_7_3 : _GEN_193; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_195 = _GEN_3935 & 4'h4 == j[3:0] ? solution_7_4 : _GEN_194; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_196 = _GEN_3935 & 4'h5 == j[3:0] ? solution_7_5 : _GEN_195; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_197 = _GEN_3935 & 4'h6 == j[3:0] ? solution_7_6 : _GEN_196; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_198 = _GEN_3935 & 4'h7 == j[3:0] ? solution_7_7 : _GEN_197; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_199 = _GEN_3935 & 4'h8 == j[3:0] ? 16'h0 : _GEN_198; // @[ivncontrol4.scala 65:{31,31}]
  wire [31:0] _GEN_201 = 3'h1 == i[2:0] ? count_1 : count_0; // @[ivncontrol4.scala 66:{33,33}]
  wire [31:0] _GEN_202 = 3'h2 == i[2:0] ? count_2 : _GEN_201; // @[ivncontrol4.scala 66:{33,33}]
  wire [31:0] _GEN_203 = 3'h3 == i[2:0] ? count_3 : _GEN_202; // @[ivncontrol4.scala 66:{33,33}]
  wire [31:0] _GEN_204 = 3'h4 == i[2:0] ? count_4 : _GEN_203; // @[ivncontrol4.scala 66:{33,33}]
  wire [31:0] _GEN_205 = 3'h5 == i[2:0] ? count_5 : _GEN_204; // @[ivncontrol4.scala 66:{33,33}]
  wire [31:0] _GEN_206 = 3'h6 == i[2:0] ? count_6 : _GEN_205; // @[ivncontrol4.scala 66:{33,33}]
  wire [31:0] _GEN_207 = 3'h7 == i[2:0] ? count_7 : _GEN_206; // @[ivncontrol4.scala 66:{33,33}]
  wire [31:0] _count_T_2 = _GEN_207 + 32'h1; // @[ivncontrol4.scala 66:33]
  wire [31:0] _GEN_208 = 3'h0 == i[2:0] ? _count_T_2 : count_0; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_209 = 3'h1 == i[2:0] ? _count_T_2 : count_1; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_210 = 3'h2 == i[2:0] ? _count_T_2 : count_2; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_211 = 3'h3 == i[2:0] ? _count_T_2 : count_3; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_212 = 3'h4 == i[2:0] ? _count_T_2 : count_4; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_213 = 3'h5 == i[2:0] ? _count_T_2 : count_5; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_214 = 3'h6 == i[2:0] ? _count_T_2 : count_6; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_215 = 3'h7 == i[2:0] ? _count_T_2 : count_7; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_216 = _GEN_199 != 16'h0 ? _GEN_208 : count_0; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_217 = _GEN_199 != 16'h0 ? _GEN_209 : count_1; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_218 = _GEN_199 != 16'h0 ? _GEN_210 : count_2; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_219 = _GEN_199 != 16'h0 ? _GEN_211 : count_3; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_220 = _GEN_199 != 16'h0 ? _GEN_212 : count_4; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_221 = _GEN_199 != 16'h0 ? _GEN_213 : count_5; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_222 = _GEN_199 != 16'h0 ? _GEN_214 : count_6; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_223 = _GEN_199 != 16'h0 ? _GEN_215 : count_7; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_224 = io_validpin ? _GEN_216 : count_0; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _GEN_225 = io_validpin ? _GEN_217 : count_1; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _GEN_226 = io_validpin ? _GEN_218 : count_2; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _GEN_227 = io_validpin ? _GEN_219 : count_3; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _GEN_228 = io_validpin ? _GEN_220 : count_4; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _GEN_229 = io_validpin ? _GEN_221 : count_5; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _GEN_230 = io_validpin ? _GEN_222 : count_6; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _GEN_231 = io_validpin ? _GEN_223 : count_7; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _i_T_1 = i + 32'h1; // @[ivncontrol4.scala 113:16]
  wire [31:0] _GEN_247 = i < 32'h7 & _io_ProcessValid_T_1 ? _i_T_1 : i; // @[ivncontrol4.scala 112:74 113:11 41:20]
  wire [31:0] _j_T_1 = j + 32'h1; // @[ivncontrol4.scala 118:16]
  wire [3:0] _GEN_264 = _io_ProcessValid_T & j == 32'h8 ? 4'h8 : 4'h0; // @[ivncontrol4.scala 120:77 121:11 129:11]
  wire [31:0] _GEN_265 = _io_ProcessValid_T & j == 32'h8 ? 32'h7 : _GEN_247; // @[ivncontrol4.scala 120:77 122:11]
  wire  _GEN_312 = _io_ProcessValid_T_2; // @[ivncontrol4.scala 153:41]
  wire [31:0] _GEN_313 = rowcount_0 != 32'h0 ? 32'h0 : pin; // @[ivncontrol4.scala 162:30 163:13 37:22]
  wire  _T_27 = rowcount_0 == 32'h0; // @[ivncontrol4.scala 165:23]
  wire [31:0] _GEN_314 = rowcount_0 == 32'h0 & rowcount_1 != 32'h0 ? 32'h1 : _GEN_313; // @[ivncontrol4.scala 165:54 166:13]
  wire  _T_32 = _T_27 & rowcount_1 == 32'h0; // @[ivncontrol4.scala 168:31]
  wire [31:0] _GEN_315 = _T_27 & rowcount_1 == 32'h0 & rowcount_2 != 32'h0 ? 32'h2 : _GEN_314; // @[ivncontrol4.scala 168:77 169:13]
  wire  _T_39 = _T_32 & rowcount_2 == 32'h0; // @[ivncontrol4.scala 171:54]
  wire [31:0] _GEN_316 = _T_32 & rowcount_2 == 32'h0 & rowcount_3 != 32'h0 ? 32'h3 : _GEN_315; // @[ivncontrol4.scala 171:100 172:13]
  wire  _T_48 = _T_39 & rowcount_3 == 32'h0; // @[ivncontrol4.scala 174:77]
  wire [31:0] _GEN_317 = _T_39 & rowcount_3 == 32'h0 & rowcount_4 != 32'h0 ? 32'h4 : _GEN_316; // @[ivncontrol4.scala 174:123 175:13]
  wire  _T_59 = _T_48 & rowcount_4 == 32'h0; // @[ivncontrol4.scala 177:100]
  wire  _T_72 = _T_59 & rowcount_5 == 32'h0; // @[ivncontrol4.scala 180:123]
  wire  valid = _io_ProcessValid_T_2; // @[ivncontrol4.scala 153:41]
  wire [32:0] _T_91 = {{1'd0}, pin}; // @[ivncontrol4.scala 191:27]
  wire [31:0] _GEN_322 = 4'h1 == _T_91[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_323 = 4'h2 == _T_91[3:0] ? rowcount_2 : _GEN_322; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_324 = 4'h3 == _T_91[3:0] ? rowcount_3 : _GEN_323; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_325 = 4'h4 == _T_91[3:0] ? rowcount_4 : _GEN_324; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_326 = 4'h5 == _T_91[3:0] ? rowcount_5 : _GEN_325; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_327 = 4'h6 == _T_91[3:0] ? rowcount_6 : _GEN_326; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_328 = 4'h7 == _T_91[3:0] ? rowcount_7 : _GEN_327; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_329 = 4'h8 == _T_91[3:0] ? rowcount_8 : _GEN_328; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_330 = 4'h9 == _T_91[3:0] ? rowcount_9 : _GEN_329; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_331 = 4'ha == _T_91[3:0] ? rowcount_10 : _GEN_330; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_332 = 4'hb == _T_91[3:0] ? rowcount_11 : _GEN_331; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_333 = 4'hc == _T_91[3:0] ? rowcount_12 : _GEN_332; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_334 = 4'hd == _T_91[3:0] ? rowcount_13 : _GEN_333; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_335 = 4'he == _T_91[3:0] ? rowcount_14 : _GEN_334; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_336 = 4'hf == _T_91[3:0] ? rowcount_15 : _GEN_335; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_449 = _GEN_336 == 32'h1 ? _T_91[31:0] : 32'h12; // @[ivncontrol4.scala 142:17 241:50 242:21]
  wire [31:0] _GEN_450 = _GEN_336 == 32'h2 ? _T_91[31:0] : _GEN_449; // @[ivncontrol4.scala 237:51 238:21]
  wire [31:0] _GEN_451 = _GEN_336 == 32'h2 ? _T_91[31:0] : 32'h5; // @[ivncontrol4.scala 142:17 237:51 239:21]
  wire [31:0] _GEN_452 = _GEN_336 == 32'h3 ? _T_91[31:0] : _GEN_450; // @[ivncontrol4.scala 232:50 233:21]
  wire [31:0] _GEN_453 = _GEN_336 == 32'h3 ? _T_91[31:0] : _GEN_451; // @[ivncontrol4.scala 232:50 234:21]
  wire [31:0] _GEN_454 = _GEN_336 == 32'h3 ? _T_91[31:0] : 32'h1e; // @[ivncontrol4.scala 142:17 232:50 235:21]
  wire [31:0] _GEN_455 = _GEN_336 == 32'h4 ? _T_91[31:0] : _GEN_452; // @[ivncontrol4.scala 224:50 225:21]
  wire [31:0] _GEN_456 = _GEN_336 == 32'h4 ? _T_91[31:0] : _GEN_453; // @[ivncontrol4.scala 224:50 226:21]
  wire [31:0] _GEN_457 = _GEN_336 == 32'h4 ? _T_91[31:0] : _GEN_454; // @[ivncontrol4.scala 224:50 227:21]
  wire [31:0] _GEN_458 = _GEN_336 == 32'h4 ? _T_91[31:0] : 32'h1f; // @[ivncontrol4.scala 142:17 224:50 228:21]
  wire [31:0] _GEN_459 = _GEN_336 == 32'h5 ? _T_91[31:0] : _GEN_455; // @[ivncontrol4.scala 217:50 218:21]
  wire [31:0] _GEN_460 = _GEN_336 == 32'h5 ? _T_91[31:0] : _GEN_456; // @[ivncontrol4.scala 217:50 219:21]
  wire [31:0] _GEN_461 = _GEN_336 == 32'h5 ? _T_91[31:0] : _GEN_457; // @[ivncontrol4.scala 217:50 220:21]
  wire [31:0] _GEN_462 = _GEN_336 == 32'h5 ? _T_91[31:0] : _GEN_458; // @[ivncontrol4.scala 217:50 221:21]
  wire [31:0] _GEN_463 = _GEN_336 == 32'h5 ? _T_91[31:0] : 32'h17; // @[ivncontrol4.scala 143:18 217:50 222:22]
  wire [31:0] _GEN_464 = _GEN_336 == 32'h6 ? _T_91[31:0] : _GEN_459; // @[ivncontrol4.scala 209:52 210:21]
  wire [31:0] _GEN_465 = _GEN_336 == 32'h6 ? _T_91[31:0] : _GEN_460; // @[ivncontrol4.scala 209:52 211:21]
  wire [31:0] _GEN_466 = _GEN_336 == 32'h6 ? _T_91[31:0] : _GEN_461; // @[ivncontrol4.scala 209:52 212:21]
  wire [31:0] _GEN_467 = _GEN_336 == 32'h6 ? _T_91[31:0] : _GEN_462; // @[ivncontrol4.scala 209:52 213:21]
  wire [31:0] _GEN_468 = _GEN_336 == 32'h6 ? _T_91[31:0] : _GEN_463; // @[ivncontrol4.scala 209:52 214:22]
  wire [31:0] _GEN_469 = _GEN_336 == 32'h6 ? _T_91[31:0] : 32'h1; // @[ivncontrol4.scala 143:18 209:52 215:22]
  wire [31:0] _GEN_470 = _GEN_336 == 32'h7 ? _T_91[31:0] : _GEN_464; // @[ivncontrol4.scala 201:52 202:21]
  wire [31:0] _GEN_471 = _GEN_336 == 32'h7 ? _T_91[31:0] : _GEN_465; // @[ivncontrol4.scala 201:52 203:21]
  wire [31:0] _GEN_472 = _GEN_336 == 32'h7 ? _T_91[31:0] : _GEN_466; // @[ivncontrol4.scala 201:52 204:21]
  wire [31:0] _GEN_473 = _GEN_336 == 32'h7 ? _T_91[31:0] : _GEN_467; // @[ivncontrol4.scala 201:52 205:21]
  wire [31:0] _GEN_474 = _GEN_336 == 32'h7 ? _T_91[31:0] : _GEN_468; // @[ivncontrol4.scala 201:52 206:22]
  wire [31:0] _GEN_475 = _GEN_336 == 32'h7 ? _T_91[31:0] : _GEN_469; // @[ivncontrol4.scala 201:52 207:22]
  wire [31:0] _GEN_476 = _GEN_336 == 32'h7 ? _T_91[31:0] : 32'h1b; // @[ivncontrol4.scala 143:18 201:52 208:22]
  wire [31:0] _GEN_477 = _GEN_336 >= 32'h8 ? _T_91[31:0] : _GEN_470; // @[ivncontrol4.scala 191:42 192:21]
  wire [31:0] _GEN_478 = _GEN_336 >= 32'h8 ? _T_91[31:0] : _GEN_471; // @[ivncontrol4.scala 191:42 193:21]
  wire [31:0] _GEN_479 = _GEN_336 >= 32'h8 ? _T_91[31:0] : _GEN_472; // @[ivncontrol4.scala 191:42 194:21]
  wire [31:0] _GEN_480 = _GEN_336 >= 32'h8 ? _T_91[31:0] : _GEN_473; // @[ivncontrol4.scala 191:42 195:21]
  wire [31:0] _GEN_481 = _GEN_336 >= 32'h8 ? _T_91[31:0] : _GEN_474; // @[ivncontrol4.scala 191:42 196:22]
  wire [31:0] _GEN_482 = _GEN_336 >= 32'h8 ? _T_91[31:0] : _GEN_475; // @[ivncontrol4.scala 191:42 197:22]
  wire [31:0] _GEN_483 = _GEN_336 >= 32'h8 ? _T_91[31:0] : _GEN_476; // @[ivncontrol4.scala 191:42 198:22]
  wire [31:0] _GEN_484 = _GEN_336 >= 32'h8 ? _T_91[31:0] : 32'ha; // @[ivncontrol4.scala 143:18 191:42 199:22]
  wire [31:0] _T_127 = 32'h8 - _GEN_336; // @[ivncontrol4.scala 245:18]
  wire [31:0] _i_vn_1_T_15 = 32'h1 + pin; // @[ivncontrol4.scala 246:29]
  wire [31:0] _GEN_597 = _T_127 == 32'h1 ? _i_vn_1_T_15 : _GEN_484; // @[ivncontrol4.scala 286:54 289:22]
  wire [31:0] _GEN_598 = _T_127 == 32'h2 ? _i_vn_1_T_15 : _GEN_483; // @[ivncontrol4.scala 281:54 284:22]
  wire [31:0] _GEN_599 = _T_127 == 32'h2 ? _i_vn_1_T_15 : _GEN_597; // @[ivncontrol4.scala 281:54 285:22]
  wire [31:0] _GEN_600 = _T_127 == 32'h3 ? _i_vn_1_T_15 : _GEN_482; // @[ivncontrol4.scala 274:54 276:22]
  wire [31:0] _GEN_601 = _T_127 == 32'h3 ? _i_vn_1_T_15 : _GEN_598; // @[ivncontrol4.scala 274:54 277:22]
  wire [31:0] _GEN_602 = _T_127 == 32'h3 ? _i_vn_1_T_15 : _GEN_599; // @[ivncontrol4.scala 274:54 278:22]
  wire [31:0] _GEN_603 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_481; // @[ivncontrol4.scala 268:54 270:22]
  wire [31:0] _GEN_604 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_600; // @[ivncontrol4.scala 268:54 271:22]
  wire [31:0] _GEN_605 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_601; // @[ivncontrol4.scala 268:54 272:22]
  wire [31:0] _GEN_606 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_602; // @[ivncontrol4.scala 268:54 273:22]
  wire [31:0] _GEN_607 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_480; // @[ivncontrol4.scala 261:54 263:21]
  wire [31:0] _GEN_608 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_603; // @[ivncontrol4.scala 261:54 264:22]
  wire [31:0] _GEN_609 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_604; // @[ivncontrol4.scala 261:54 265:22]
  wire [31:0] _GEN_610 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_605; // @[ivncontrol4.scala 261:54 266:22]
  wire [31:0] _GEN_611 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_606; // @[ivncontrol4.scala 261:54 267:22]
  wire [31:0] _GEN_612 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_479; // @[ivncontrol4.scala 254:54 255:22]
  wire [31:0] _GEN_613 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_607; // @[ivncontrol4.scala 254:54 256:21]
  wire [31:0] _GEN_614 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_608; // @[ivncontrol4.scala 254:54 257:22]
  wire [31:0] _GEN_615 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_609; // @[ivncontrol4.scala 254:54 258:22]
  wire [31:0] _GEN_616 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_610; // @[ivncontrol4.scala 254:54 259:22]
  wire [31:0] _GEN_617 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_611; // @[ivncontrol4.scala 254:54 260:22]
  wire [31:0] _GEN_618 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_478; // @[ivncontrol4.scala 245:49 246:22]
  wire [31:0] _GEN_619 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_612; // @[ivncontrol4.scala 245:49 247:21]
  wire [31:0] _GEN_620 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_613; // @[ivncontrol4.scala 245:49 248:21]
  wire [31:0] _GEN_621 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_614; // @[ivncontrol4.scala 245:49 249:22]
  wire [31:0] _GEN_622 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_615; // @[ivncontrol4.scala 245:49 250:22]
  wire [31:0] _GEN_623 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_616; // @[ivncontrol4.scala 245:49 251:22]
  wire [31:0] _GEN_624 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_617; // @[ivncontrol4.scala 245:49 252:22]
  wire [31:0] _GEN_642 = 4'h1 == _i_vn_1_T_15[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_643 = 4'h2 == _i_vn_1_T_15[3:0] ? rowcount_2 : _GEN_642; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_644 = 4'h3 == _i_vn_1_T_15[3:0] ? rowcount_3 : _GEN_643; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_645 = 4'h4 == _i_vn_1_T_15[3:0] ? rowcount_4 : _GEN_644; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_646 = 4'h5 == _i_vn_1_T_15[3:0] ? rowcount_5 : _GEN_645; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_647 = 4'h6 == _i_vn_1_T_15[3:0] ? rowcount_6 : _GEN_646; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_648 = 4'h7 == _i_vn_1_T_15[3:0] ? rowcount_7 : _GEN_647; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_649 = 4'h8 == _i_vn_1_T_15[3:0] ? rowcount_8 : _GEN_648; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_650 = 4'h9 == _i_vn_1_T_15[3:0] ? rowcount_9 : _GEN_649; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_651 = 4'ha == _i_vn_1_T_15[3:0] ? rowcount_10 : _GEN_650; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_652 = 4'hb == _i_vn_1_T_15[3:0] ? rowcount_11 : _GEN_651; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_653 = 4'hc == _i_vn_1_T_15[3:0] ? rowcount_12 : _GEN_652; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_654 = 4'hd == _i_vn_1_T_15[3:0] ? rowcount_13 : _GEN_653; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_655 = 4'he == _i_vn_1_T_15[3:0] ? rowcount_14 : _GEN_654; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_656 = 4'hf == _i_vn_1_T_15[3:0] ? rowcount_15 : _GEN_655; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _T_172 = _GEN_336 + _GEN_656; // @[ivncontrol4.scala 292:41]
  wire [31:0] _T_174 = 32'h8 - _T_172; // @[ivncontrol4.scala 292:18]
  wire [31:0] _i_vn_1_T_17 = 32'h2 + pin; // @[ivncontrol4.scala 293:29]
  wire [31:0] _GEN_849 = _T_174 == 32'h1 ? _i_vn_1_T_17 : _GEN_624; // @[ivncontrol4.scala 335:78 338:22]
  wire [31:0] _GEN_850 = _T_174 == 32'h2 ? _i_vn_1_T_17 : _GEN_623; // @[ivncontrol4.scala 329:76 332:22]
  wire [31:0] _GEN_851 = _T_174 == 32'h2 ? _i_vn_1_T_17 : _GEN_849; // @[ivncontrol4.scala 329:76 333:22]
  wire [31:0] _GEN_852 = _T_174 == 32'h3 ? _i_vn_1_T_17 : _GEN_622; // @[ivncontrol4.scala 322:78 324:23]
  wire [31:0] _GEN_853 = _T_174 == 32'h3 ? _i_vn_1_T_17 : _GEN_850; // @[ivncontrol4.scala 322:78 325:22]
  wire [31:0] _GEN_854 = _T_174 == 32'h3 ? _i_vn_1_T_17 : _GEN_851; // @[ivncontrol4.scala 322:78 326:22]
  wire [31:0] _GEN_855 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_621; // @[ivncontrol4.scala 316:78 318:22]
  wire [31:0] _GEN_856 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_852; // @[ivncontrol4.scala 316:78 319:22]
  wire [31:0] _GEN_857 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_853; // @[ivncontrol4.scala 316:78 320:22]
  wire [31:0] _GEN_858 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_854; // @[ivncontrol4.scala 316:78 321:22]
  wire [31:0] _GEN_859 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_620; // @[ivncontrol4.scala 309:76 311:23]
  wire [31:0] _GEN_860 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_855; // @[ivncontrol4.scala 309:76 312:22]
  wire [31:0] _GEN_861 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_856; // @[ivncontrol4.scala 309:76 313:22]
  wire [31:0] _GEN_862 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_857; // @[ivncontrol4.scala 309:76 314:22]
  wire [31:0] _GEN_863 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_858; // @[ivncontrol4.scala 309:76 315:22]
  wire [31:0] _GEN_864 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_619; // @[ivncontrol4.scala 301:77 303:22]
  wire [31:0] _GEN_865 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_859; // @[ivncontrol4.scala 301:77 304:21]
  wire [31:0] _GEN_866 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_860; // @[ivncontrol4.scala 301:77 305:22]
  wire [31:0] _GEN_867 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_861; // @[ivncontrol4.scala 301:77 306:22]
  wire [31:0] _GEN_868 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_862; // @[ivncontrol4.scala 301:77 307:22]
  wire [31:0] _GEN_869 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_863; // @[ivncontrol4.scala 301:77 308:22]
  wire [31:0] _GEN_870 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_618; // @[ivncontrol4.scala 292:73 293:22]
  wire [31:0] _GEN_871 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_864; // @[ivncontrol4.scala 292:73 294:21]
  wire [31:0] _GEN_872 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_865; // @[ivncontrol4.scala 292:73 295:21]
  wire [31:0] _GEN_873 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_866; // @[ivncontrol4.scala 292:73 296:22]
  wire [31:0] _GEN_874 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_867; // @[ivncontrol4.scala 292:73 297:22]
  wire [31:0] _GEN_875 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_868; // @[ivncontrol4.scala 292:73 298:22]
  wire [31:0] _GEN_876 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_869; // @[ivncontrol4.scala 292:73 299:22]
  wire [31:0] _GEN_910 = 4'h1 == _i_vn_1_T_17[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_911 = 4'h2 == _i_vn_1_T_17[3:0] ? rowcount_2 : _GEN_910; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_912 = 4'h3 == _i_vn_1_T_17[3:0] ? rowcount_3 : _GEN_911; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_913 = 4'h4 == _i_vn_1_T_17[3:0] ? rowcount_4 : _GEN_912; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_914 = 4'h5 == _i_vn_1_T_17[3:0] ? rowcount_5 : _GEN_913; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_915 = 4'h6 == _i_vn_1_T_17[3:0] ? rowcount_6 : _GEN_914; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_916 = 4'h7 == _i_vn_1_T_17[3:0] ? rowcount_7 : _GEN_915; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_917 = 4'h8 == _i_vn_1_T_17[3:0] ? rowcount_8 : _GEN_916; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_918 = 4'h9 == _i_vn_1_T_17[3:0] ? rowcount_9 : _GEN_917; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_919 = 4'ha == _i_vn_1_T_17[3:0] ? rowcount_10 : _GEN_918; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_920 = 4'hb == _i_vn_1_T_17[3:0] ? rowcount_11 : _GEN_919; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_921 = 4'hc == _i_vn_1_T_17[3:0] ? rowcount_12 : _GEN_920; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_922 = 4'hd == _i_vn_1_T_17[3:0] ? rowcount_13 : _GEN_921; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_923 = 4'he == _i_vn_1_T_17[3:0] ? rowcount_14 : _GEN_922; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_924 = 4'hf == _i_vn_1_T_17[3:0] ? rowcount_15 : _GEN_923; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _T_254 = _T_172 + _GEN_924; // @[ivncontrol4.scala 343:62]
  wire [31:0] _T_256 = 32'h8 - _T_254; // @[ivncontrol4.scala 343:17]
  wire [31:0] _i_vn_1_T_19 = 32'h3 + pin; // @[ivncontrol4.scala 344:29]
  wire [31:0] _GEN_1213 = _T_256 == 32'h1 ? _i_vn_1_T_19 : _GEN_876; // @[ivncontrol4.scala 386:100 389:22]
  wire [31:0] _GEN_1214 = _T_256 == 32'h2 ? _i_vn_1_T_19 : _GEN_875; // @[ivncontrol4.scala 380:98 383:22]
  wire [31:0] _GEN_1215 = _T_256 == 32'h2 ? _i_vn_1_T_19 : _GEN_1213; // @[ivncontrol4.scala 380:98 384:22]
  wire [31:0] _GEN_1216 = _T_256 == 32'h3 ? _i_vn_1_T_19 : _GEN_874; // @[ivncontrol4.scala 373:100 375:23]
  wire [31:0] _GEN_1217 = _T_256 == 32'h3 ? _i_vn_1_T_19 : _GEN_1214; // @[ivncontrol4.scala 373:100 376:22]
  wire [31:0] _GEN_1218 = _T_256 == 32'h3 ? _i_vn_1_T_19 : _GEN_1215; // @[ivncontrol4.scala 373:100 377:22]
  wire [31:0] _GEN_1219 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_873; // @[ivncontrol4.scala 367:100 369:22]
  wire [31:0] _GEN_1220 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_1216; // @[ivncontrol4.scala 367:100 370:22]
  wire [31:0] _GEN_1221 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_1217; // @[ivncontrol4.scala 367:100 371:22]
  wire [31:0] _GEN_1222 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_1218; // @[ivncontrol4.scala 367:100 372:22]
  wire [31:0] _GEN_1223 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_872; // @[ivncontrol4.scala 360:98 362:23]
  wire [31:0] _GEN_1224 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1219; // @[ivncontrol4.scala 360:98 363:22]
  wire [31:0] _GEN_1225 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1220; // @[ivncontrol4.scala 360:98 364:22]
  wire [31:0] _GEN_1226 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1221; // @[ivncontrol4.scala 360:98 365:22]
  wire [31:0] _GEN_1227 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1222; // @[ivncontrol4.scala 360:98 366:22]
  wire [31:0] _GEN_1228 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_871; // @[ivncontrol4.scala 352:99 354:22]
  wire [31:0] _GEN_1229 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1223; // @[ivncontrol4.scala 352:99 355:21]
  wire [31:0] _GEN_1230 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1224; // @[ivncontrol4.scala 352:99 356:22]
  wire [31:0] _GEN_1231 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1225; // @[ivncontrol4.scala 352:99 357:22]
  wire [31:0] _GEN_1232 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1226; // @[ivncontrol4.scala 352:99 358:22]
  wire [31:0] _GEN_1233 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1227; // @[ivncontrol4.scala 352:99 359:22]
  wire [31:0] _GEN_1234 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_870; // @[ivncontrol4.scala 343:94 344:22]
  wire [31:0] _GEN_1235 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1228; // @[ivncontrol4.scala 343:94 345:21]
  wire [31:0] _GEN_1236 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1229; // @[ivncontrol4.scala 343:94 346:21]
  wire [31:0] _GEN_1237 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1230; // @[ivncontrol4.scala 343:94 347:22]
  wire [31:0] _GEN_1238 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1231; // @[ivncontrol4.scala 343:94 348:22]
  wire [31:0] _GEN_1239 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1232; // @[ivncontrol4.scala 343:94 349:22]
  wire [31:0] _GEN_1240 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1233; // @[ivncontrol4.scala 343:94 350:22]
  wire [31:0] _GEN_1290 = 4'h1 == _i_vn_1_T_19[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1291 = 4'h2 == _i_vn_1_T_19[3:0] ? rowcount_2 : _GEN_1290; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1292 = 4'h3 == _i_vn_1_T_19[3:0] ? rowcount_3 : _GEN_1291; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1293 = 4'h4 == _i_vn_1_T_19[3:0] ? rowcount_4 : _GEN_1292; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1294 = 4'h5 == _i_vn_1_T_19[3:0] ? rowcount_5 : _GEN_1293; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1295 = 4'h6 == _i_vn_1_T_19[3:0] ? rowcount_6 : _GEN_1294; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1296 = 4'h7 == _i_vn_1_T_19[3:0] ? rowcount_7 : _GEN_1295; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1297 = 4'h8 == _i_vn_1_T_19[3:0] ? rowcount_8 : _GEN_1296; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1298 = 4'h9 == _i_vn_1_T_19[3:0] ? rowcount_9 : _GEN_1297; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1299 = 4'ha == _i_vn_1_T_19[3:0] ? rowcount_10 : _GEN_1298; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1300 = 4'hb == _i_vn_1_T_19[3:0] ? rowcount_11 : _GEN_1299; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1301 = 4'hc == _i_vn_1_T_19[3:0] ? rowcount_12 : _GEN_1300; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1302 = 4'hd == _i_vn_1_T_19[3:0] ? rowcount_13 : _GEN_1301; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1303 = 4'he == _i_vn_1_T_19[3:0] ? rowcount_14 : _GEN_1302; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1304 = 4'hf == _i_vn_1_T_19[3:0] ? rowcount_15 : _GEN_1303; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _T_371 = _T_254 + _GEN_1304; // @[ivncontrol4.scala 393:86]
  wire [31:0] _T_373 = 32'h8 - _T_371; // @[ivncontrol4.scala 393:19]
  wire [31:0] _i_vn_1_T_21 = 32'h4 + pin; // @[ivncontrol4.scala 394:29]
  wire [31:0] _GEN_1689 = _T_373 == 32'h1 ? _i_vn_1_T_21 : _GEN_1240; // @[ivncontrol4.scala 436:122 439:22]
  wire [31:0] _GEN_1690 = _T_373 == 32'h2 ? _i_vn_1_T_21 : _GEN_1239; // @[ivncontrol4.scala 430:121 433:22]
  wire [31:0] _GEN_1691 = _T_373 == 32'h2 ? _i_vn_1_T_21 : _GEN_1689; // @[ivncontrol4.scala 430:121 434:22]
  wire [31:0] _GEN_1692 = _T_373 == 32'h3 ? _i_vn_1_T_21 : _GEN_1238; // @[ivncontrol4.scala 423:123 425:23]
  wire [31:0] _GEN_1693 = _T_373 == 32'h3 ? _i_vn_1_T_21 : _GEN_1690; // @[ivncontrol4.scala 423:123 426:22]
  wire [31:0] _GEN_1694 = _T_373 == 32'h3 ? _i_vn_1_T_21 : _GEN_1691; // @[ivncontrol4.scala 423:123 427:22]
  wire [31:0] _GEN_1695 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1237; // @[ivncontrol4.scala 417:122 419:22]
  wire [31:0] _GEN_1696 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1692; // @[ivncontrol4.scala 417:122 420:22]
  wire [31:0] _GEN_1697 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1693; // @[ivncontrol4.scala 417:122 421:22]
  wire [31:0] _GEN_1698 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1694; // @[ivncontrol4.scala 417:122 422:22]
  wire [31:0] _GEN_1699 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1236; // @[ivncontrol4.scala 410:121 412:23]
  wire [31:0] _GEN_1700 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1695; // @[ivncontrol4.scala 410:121 413:22]
  wire [31:0] _GEN_1701 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1696; // @[ivncontrol4.scala 410:121 414:22]
  wire [31:0] _GEN_1702 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1697; // @[ivncontrol4.scala 410:121 415:22]
  wire [31:0] _GEN_1703 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1698; // @[ivncontrol4.scala 410:121 416:22]
  wire [31:0] _GEN_1704 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1235; // @[ivncontrol4.scala 402:121 404:22]
  wire [31:0] _GEN_1705 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1699; // @[ivncontrol4.scala 402:121 405:21]
  wire [31:0] _GEN_1706 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1700; // @[ivncontrol4.scala 402:121 406:22]
  wire [31:0] _GEN_1707 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1701; // @[ivncontrol4.scala 402:121 407:22]
  wire [31:0] _GEN_1708 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1702; // @[ivncontrol4.scala 402:121 408:22]
  wire [31:0] _GEN_1709 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1703; // @[ivncontrol4.scala 402:121 409:22]
  wire [31:0] _GEN_1710 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1234; // @[ivncontrol4.scala 393:118 394:22]
  wire [31:0] _GEN_1711 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1704; // @[ivncontrol4.scala 393:118 395:21]
  wire [31:0] _GEN_1712 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1705; // @[ivncontrol4.scala 393:118 396:21]
  wire [31:0] _GEN_1713 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1706; // @[ivncontrol4.scala 393:118 397:22]
  wire [31:0] _GEN_1714 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1707; // @[ivncontrol4.scala 393:118 398:22]
  wire [31:0] _GEN_1715 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1708; // @[ivncontrol4.scala 393:118 399:22]
  wire [31:0] _GEN_1716 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1709; // @[ivncontrol4.scala 393:118 400:22]
  wire [31:0] _GEN_1782 = 4'h1 == _i_vn_1_T_21[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1783 = 4'h2 == _i_vn_1_T_21[3:0] ? rowcount_2 : _GEN_1782; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1784 = 4'h3 == _i_vn_1_T_21[3:0] ? rowcount_3 : _GEN_1783; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1785 = 4'h4 == _i_vn_1_T_21[3:0] ? rowcount_4 : _GEN_1784; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1786 = 4'h5 == _i_vn_1_T_21[3:0] ? rowcount_5 : _GEN_1785; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1787 = 4'h6 == _i_vn_1_T_21[3:0] ? rowcount_6 : _GEN_1786; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1788 = 4'h7 == _i_vn_1_T_21[3:0] ? rowcount_7 : _GEN_1787; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1789 = 4'h8 == _i_vn_1_T_21[3:0] ? rowcount_8 : _GEN_1788; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1790 = 4'h9 == _i_vn_1_T_21[3:0] ? rowcount_9 : _GEN_1789; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1791 = 4'ha == _i_vn_1_T_21[3:0] ? rowcount_10 : _GEN_1790; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1792 = 4'hb == _i_vn_1_T_21[3:0] ? rowcount_11 : _GEN_1791; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1793 = 4'hc == _i_vn_1_T_21[3:0] ? rowcount_12 : _GEN_1792; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1794 = 4'hd == _i_vn_1_T_21[3:0] ? rowcount_13 : _GEN_1793; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1795 = 4'he == _i_vn_1_T_21[3:0] ? rowcount_14 : _GEN_1794; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1796 = 4'hf == _i_vn_1_T_21[3:0] ? rowcount_15 : _GEN_1795; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _T_523 = _T_371 + _GEN_1796; // @[ivncontrol4.scala 443:108]
  wire [31:0] _T_525 = 32'h8 - _T_523; // @[ivncontrol4.scala 443:19]
  wire [31:0] _i_vn_1_T_23 = 32'h5 + pin; // @[ivncontrol4.scala 444:29]
  wire [31:0] _GEN_2277 = _T_525 == 32'h1 ? _i_vn_1_T_23 : _GEN_1716; // @[ivncontrol4.scala 486:144 489:22]
  wire [31:0] _GEN_2278 = _T_525 == 32'h2 ? _i_vn_1_T_23 : _GEN_1715; // @[ivncontrol4.scala 480:143 483:22]
  wire [31:0] _GEN_2279 = _T_525 == 32'h2 ? _i_vn_1_T_23 : _GEN_2277; // @[ivncontrol4.scala 480:143 484:22]
  wire [31:0] _GEN_2280 = _T_525 == 32'h3 ? _i_vn_1_T_23 : _GEN_1714; // @[ivncontrol4.scala 473:145 475:23]
  wire [31:0] _GEN_2281 = _T_525 == 32'h3 ? _i_vn_1_T_23 : _GEN_2278; // @[ivncontrol4.scala 473:145 476:22]
  wire [31:0] _GEN_2282 = _T_525 == 32'h3 ? _i_vn_1_T_23 : _GEN_2279; // @[ivncontrol4.scala 473:145 477:22]
  wire [31:0] _GEN_2283 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_1713; // @[ivncontrol4.scala 467:143 469:22]
  wire [31:0] _GEN_2284 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_2280; // @[ivncontrol4.scala 467:143 470:22]
  wire [31:0] _GEN_2285 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_2281; // @[ivncontrol4.scala 467:143 471:22]
  wire [31:0] _GEN_2286 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_2282; // @[ivncontrol4.scala 467:143 472:22]
  wire [31:0] _GEN_2287 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_1712; // @[ivncontrol4.scala 460:143 462:23]
  wire [31:0] _GEN_2288 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2283; // @[ivncontrol4.scala 460:143 463:22]
  wire [31:0] _GEN_2289 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2284; // @[ivncontrol4.scala 460:143 464:22]
  wire [31:0] _GEN_2290 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2285; // @[ivncontrol4.scala 460:143 465:22]
  wire [31:0] _GEN_2291 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2286; // @[ivncontrol4.scala 460:143 466:22]
  wire [31:0] _GEN_2292 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_1711; // @[ivncontrol4.scala 452:143 454:22]
  wire [31:0] _GEN_2293 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2287; // @[ivncontrol4.scala 452:143 455:21]
  wire [31:0] _GEN_2294 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2288; // @[ivncontrol4.scala 452:143 456:22]
  wire [31:0] _GEN_2295 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2289; // @[ivncontrol4.scala 452:143 457:22]
  wire [31:0] _GEN_2296 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2290; // @[ivncontrol4.scala 452:143 458:22]
  wire [31:0] _GEN_2297 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2291; // @[ivncontrol4.scala 452:143 459:22]
  wire [31:0] _GEN_2298 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_1710; // @[ivncontrol4.scala 443:140 444:22]
  wire [31:0] _GEN_2299 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2292; // @[ivncontrol4.scala 443:140 445:21]
  wire [31:0] _GEN_2300 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2293; // @[ivncontrol4.scala 443:140 446:21]
  wire [31:0] _GEN_2301 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2294; // @[ivncontrol4.scala 443:140 447:22]
  wire [31:0] _GEN_2302 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2295; // @[ivncontrol4.scala 443:140 448:22]
  wire [31:0] _GEN_2303 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2296; // @[ivncontrol4.scala 443:140 449:22]
  wire [31:0] _GEN_2304 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2297; // @[ivncontrol4.scala 443:140 450:22]
  wire [31:0] _GEN_2386 = 4'h1 == _i_vn_1_T_23[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2387 = 4'h2 == _i_vn_1_T_23[3:0] ? rowcount_2 : _GEN_2386; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2388 = 4'h3 == _i_vn_1_T_23[3:0] ? rowcount_3 : _GEN_2387; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2389 = 4'h4 == _i_vn_1_T_23[3:0] ? rowcount_4 : _GEN_2388; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2390 = 4'h5 == _i_vn_1_T_23[3:0] ? rowcount_5 : _GEN_2389; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2391 = 4'h6 == _i_vn_1_T_23[3:0] ? rowcount_6 : _GEN_2390; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2392 = 4'h7 == _i_vn_1_T_23[3:0] ? rowcount_7 : _GEN_2391; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2393 = 4'h8 == _i_vn_1_T_23[3:0] ? rowcount_8 : _GEN_2392; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2394 = 4'h9 == _i_vn_1_T_23[3:0] ? rowcount_9 : _GEN_2393; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2395 = 4'ha == _i_vn_1_T_23[3:0] ? rowcount_10 : _GEN_2394; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2396 = 4'hb == _i_vn_1_T_23[3:0] ? rowcount_11 : _GEN_2395; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2397 = 4'hc == _i_vn_1_T_23[3:0] ? rowcount_12 : _GEN_2396; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2398 = 4'hd == _i_vn_1_T_23[3:0] ? rowcount_13 : _GEN_2397; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2399 = 4'he == _i_vn_1_T_23[3:0] ? rowcount_14 : _GEN_2398; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2400 = 4'hf == _i_vn_1_T_23[3:0] ? rowcount_15 : _GEN_2399; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _T_710 = _T_523 + _GEN_2400; // @[ivncontrol4.scala 494:130]
  wire [31:0] _T_712 = 32'h8 - _T_710; // @[ivncontrol4.scala 494:19]
  wire [31:0] _i_vn_1_T_25 = 32'h6 + pin; // @[ivncontrol4.scala 495:29]
  wire [31:0] _GEN_2977 = _T_712 == 32'h1 ? _i_vn_1_T_25 : _GEN_2304; // @[ivncontrol4.scala 537:166 540:22]
  wire [31:0] _GEN_2978 = _T_712 == 32'h2 ? _i_vn_1_T_25 : _GEN_2303; // @[ivncontrol4.scala 531:166 534:22]
  wire [31:0] _GEN_2979 = _T_712 == 32'h2 ? _i_vn_1_T_25 : _GEN_2977; // @[ivncontrol4.scala 531:166 535:22]
  wire [31:0] _GEN_2980 = _T_712 == 32'h3 ? _i_vn_1_T_25 : _GEN_2302; // @[ivncontrol4.scala 524:168 526:23]
  wire [31:0] _GEN_2981 = _T_712 == 32'h3 ? _i_vn_1_T_25 : _GEN_2978; // @[ivncontrol4.scala 524:168 527:22]
  wire [31:0] _GEN_2982 = _T_712 == 32'h3 ? _i_vn_1_T_25 : _GEN_2979; // @[ivncontrol4.scala 524:168 528:22]
  wire [31:0] _GEN_2983 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2301; // @[ivncontrol4.scala 518:166 520:22]
  wire [31:0] _GEN_2984 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2980; // @[ivncontrol4.scala 518:166 521:22]
  wire [31:0] _GEN_2985 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2981; // @[ivncontrol4.scala 518:166 522:22]
  wire [31:0] _GEN_2986 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2982; // @[ivncontrol4.scala 518:166 523:22]
  wire [31:0] _GEN_2987 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2300; // @[ivncontrol4.scala 511:166 513:23]
  wire [31:0] _GEN_2988 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2983; // @[ivncontrol4.scala 511:166 514:22]
  wire [31:0] _GEN_2989 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2984; // @[ivncontrol4.scala 511:166 515:22]
  wire [31:0] _GEN_2990 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2985; // @[ivncontrol4.scala 511:166 516:22]
  wire [31:0] _GEN_2991 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2986; // @[ivncontrol4.scala 511:166 517:22]
  wire [31:0] _GEN_2992 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2299; // @[ivncontrol4.scala 503:166 505:22]
  wire [31:0] _GEN_2993 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2987; // @[ivncontrol4.scala 503:166 506:21]
  wire [31:0] _GEN_2994 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2988; // @[ivncontrol4.scala 503:166 507:22]
  wire [31:0] _GEN_2995 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2989; // @[ivncontrol4.scala 503:166 508:22]
  wire [31:0] _GEN_2996 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2990; // @[ivncontrol4.scala 503:166 509:22]
  wire [31:0] _GEN_2997 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2991; // @[ivncontrol4.scala 503:166 510:22]
  wire [31:0] _GEN_2998 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2298; // @[ivncontrol4.scala 494:162 495:22]
  wire [31:0] _GEN_2999 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2992; // @[ivncontrol4.scala 494:162 496:21]
  wire [31:0] _GEN_3000 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2993; // @[ivncontrol4.scala 494:162 497:21]
  wire [31:0] _GEN_3001 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2994; // @[ivncontrol4.scala 494:162 498:22]
  wire [31:0] _GEN_3002 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2995; // @[ivncontrol4.scala 494:162 499:22]
  wire [31:0] _GEN_3003 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2996; // @[ivncontrol4.scala 494:162 500:22]
  wire [31:0] _GEN_3004 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2997; // @[ivncontrol4.scala 494:162 501:22]
  wire [31:0] _GEN_3102 = 4'h1 == _i_vn_1_T_25[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3103 = 4'h2 == _i_vn_1_T_25[3:0] ? rowcount_2 : _GEN_3102; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3104 = 4'h3 == _i_vn_1_T_25[3:0] ? rowcount_3 : _GEN_3103; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3105 = 4'h4 == _i_vn_1_T_25[3:0] ? rowcount_4 : _GEN_3104; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3106 = 4'h5 == _i_vn_1_T_25[3:0] ? rowcount_5 : _GEN_3105; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3107 = 4'h6 == _i_vn_1_T_25[3:0] ? rowcount_6 : _GEN_3106; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3108 = 4'h7 == _i_vn_1_T_25[3:0] ? rowcount_7 : _GEN_3107; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3109 = 4'h8 == _i_vn_1_T_25[3:0] ? rowcount_8 : _GEN_3108; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3110 = 4'h9 == _i_vn_1_T_25[3:0] ? rowcount_9 : _GEN_3109; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3111 = 4'ha == _i_vn_1_T_25[3:0] ? rowcount_10 : _GEN_3110; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3112 = 4'hb == _i_vn_1_T_25[3:0] ? rowcount_11 : _GEN_3111; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3113 = 4'hc == _i_vn_1_T_25[3:0] ? rowcount_12 : _GEN_3112; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3114 = 4'hd == _i_vn_1_T_25[3:0] ? rowcount_13 : _GEN_3113; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3115 = 4'he == _i_vn_1_T_25[3:0] ? rowcount_14 : _GEN_3114; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3116 = 4'hf == _i_vn_1_T_25[3:0] ? rowcount_15 : _GEN_3115; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _T_932 = _T_710 + _GEN_3116; // @[ivncontrol4.scala 545:152]
  wire [31:0] _T_934 = 32'h8 - _T_932; // @[ivncontrol4.scala 545:19]
  wire [31:0] _i_vn_1_T_27 = 32'h7 + pin; // @[ivncontrol4.scala 546:29]
  wire [31:0] _GEN_3789 = _T_934 == 32'h1 ? _i_vn_1_T_27 : _GEN_3004; // @[ivncontrol4.scala 588:188 591:22]
  wire [31:0] _GEN_3790 = _T_934 == 32'h2 ? _i_vn_1_T_27 : _GEN_3003; // @[ivncontrol4.scala 582:188 585:22]
  wire [31:0] _GEN_3791 = _T_934 == 32'h2 ? _i_vn_1_T_27 : _GEN_3789; // @[ivncontrol4.scala 582:188 586:22]
  wire [31:0] _GEN_3792 = _T_934 == 32'h3 ? _i_vn_1_T_27 : _GEN_3002; // @[ivncontrol4.scala 575:190 577:23]
  wire [31:0] _GEN_3793 = _T_934 == 32'h3 ? _i_vn_1_T_27 : _GEN_3790; // @[ivncontrol4.scala 575:190 578:22]
  wire [31:0] _GEN_3794 = _T_934 == 32'h3 ? _i_vn_1_T_27 : _GEN_3791; // @[ivncontrol4.scala 575:190 579:22]
  wire [31:0] _GEN_3795 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_3001; // @[ivncontrol4.scala 569:188 571:22]
  wire [31:0] _GEN_3796 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_3792; // @[ivncontrol4.scala 569:188 572:22]
  wire [31:0] _GEN_3797 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_3793; // @[ivncontrol4.scala 569:188 573:22]
  wire [31:0] _GEN_3798 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_3794; // @[ivncontrol4.scala 569:188 574:22]
  wire [31:0] _GEN_3799 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3000; // @[ivncontrol4.scala 562:188 564:23]
  wire [31:0] _GEN_3800 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3795; // @[ivncontrol4.scala 562:188 565:22]
  wire [31:0] _GEN_3801 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3796; // @[ivncontrol4.scala 562:188 566:22]
  wire [31:0] _GEN_3802 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3797; // @[ivncontrol4.scala 562:188 567:22]
  wire [31:0] _GEN_3803 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3798; // @[ivncontrol4.scala 562:188 568:22]
  wire [31:0] _GEN_3804 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_2999; // @[ivncontrol4.scala 554:188 556:22]
  wire [31:0] _GEN_3805 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3799; // @[ivncontrol4.scala 554:188 557:21]
  wire [31:0] _GEN_3806 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3800; // @[ivncontrol4.scala 554:188 558:22]
  wire [31:0] _GEN_3807 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3801; // @[ivncontrol4.scala 554:188 559:22]
  wire [31:0] _GEN_3808 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3802; // @[ivncontrol4.scala 554:188 560:22]
  wire [31:0] _GEN_3809 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3803; // @[ivncontrol4.scala 554:188 561:22]
  wire [31:0] _GEN_3810 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_2998; // @[ivncontrol4.scala 545:184 546:22]
  wire [31:0] _GEN_3811 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3804; // @[ivncontrol4.scala 545:184 547:21]
  wire [31:0] _GEN_3812 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3805; // @[ivncontrol4.scala 545:184 548:21]
  wire [31:0] _GEN_3813 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3806; // @[ivncontrol4.scala 545:184 549:22]
  wire [31:0] _GEN_3814 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3807; // @[ivncontrol4.scala 545:184 550:22]
  wire [31:0] _GEN_3815 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3808; // @[ivncontrol4.scala 545:184 551:22]
  wire [31:0] _GEN_3816 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3809; // @[ivncontrol4.scala 545:184 552:22]
  wire [31:0] _GEN_3817 = _GEN_312 ? _GEN_477 : 32'h12; // @[ivncontrol4.scala 142:17 189:28]
  wire [31:0] _GEN_3818 = _GEN_312 ? _GEN_3810 : 32'h5; // @[ivncontrol4.scala 142:17 189:28]
  wire [31:0] _GEN_3819 = _GEN_312 ? _GEN_3811 : 32'h1e; // @[ivncontrol4.scala 142:17 189:28]
  wire [31:0] _GEN_3820 = _GEN_312 ? _GEN_3812 : 32'h1f; // @[ivncontrol4.scala 142:17 189:28]
  wire [31:0] _GEN_3821 = _GEN_312 ? _GEN_3813 : 32'h17; // @[ivncontrol4.scala 143:18 189:28]
  wire [31:0] _GEN_3822 = _GEN_312 ? _GEN_3814 : 32'h1; // @[ivncontrol4.scala 143:18 189:28]
  wire [31:0] _GEN_3823 = _GEN_312 ? _GEN_3815 : 32'h1b; // @[ivncontrol4.scala 143:18 189:28]
  wire [31:0] _GEN_3824 = _GEN_312 ? _GEN_3816 : 32'ha; // @[ivncontrol4.scala 143:18 189:28]
  wire  valid1 = 1'h0;
  wire [31:0] _GEN_4221 = reset ? 32'h0 : _GEN_3817; // @[ivncontrol4.scala 17:{23,23}]
  wire [31:0] _GEN_4222 = reset ? 32'h0 : _GEN_3818; // @[ivncontrol4.scala 17:{23,23}]
  wire [31:0] _GEN_4223 = reset ? 32'h0 : _GEN_3819; // @[ivncontrol4.scala 17:{23,23}]
  wire [31:0] _GEN_4224 = reset ? 32'h0 : _GEN_3820; // @[ivncontrol4.scala 17:{23,23}]
  wire [31:0] _GEN_4225 = reset ? 32'h0 : _GEN_3821; // @[ivncontrol4.scala 18:{24,24}]
  wire [31:0] _GEN_4226 = reset ? 32'h0 : _GEN_3822; // @[ivncontrol4.scala 18:{24,24}]
  wire [31:0] _GEN_4227 = reset ? 32'h0 : _GEN_3823; // @[ivncontrol4.scala 18:{24,24}]
  wire [31:0] _GEN_4228 = reset ? 32'h0 : _GEN_3824; // @[ivncontrol4.scala 18:{24,24}]
  assign io_o_vn_0 = i_vn_0; // @[ivncontrol4.scala 138:13]
  assign io_o_vn_1 = i_vn_1; // @[ivncontrol4.scala 138:13]
  assign io_o_vn_2 = i_vn_2; // @[ivncontrol4.scala 138:13]
  assign io_o_vn_3 = i_vn_3; // @[ivncontrol4.scala 138:13]
  assign io_o_vn2_0 = i_vn2_0; // @[ivncontrol4.scala 139:14]
  assign io_o_vn2_1 = i_vn2_1; // @[ivncontrol4.scala 139:14]
  assign io_o_vn2_2 = i_vn2_2; // @[ivncontrol4.scala 139:14]
  assign io_o_vn2_3 = i_vn2_3; // @[ivncontrol4.scala 139:14]
  always @(posedge clock) begin
    i_vn_0 <= _GEN_4221[4:0]; // @[ivncontrol4.scala 17:{23,23}]
    i_vn_1 <= _GEN_4222[4:0]; // @[ivncontrol4.scala 17:{23,23}]
    i_vn_2 <= _GEN_4223[4:0]; // @[ivncontrol4.scala 17:{23,23}]
    i_vn_3 <= _GEN_4224[4:0]; // @[ivncontrol4.scala 17:{23,23}]
    i_vn2_0 <= _GEN_4225[4:0]; // @[ivncontrol4.scala 18:{24,24}]
    i_vn2_1 <= _GEN_4226[4:0]; // @[ivncontrol4.scala 18:{24,24}]
    i_vn2_2 <= _GEN_4227[4:0]; // @[ivncontrol4.scala 18:{24,24}]
    i_vn2_3 <= _GEN_4228[4:0]; // @[ivncontrol4.scala 18:{24,24}]
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_0 <= io_Stationary_matrix_0_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_1 <= io_Stationary_matrix_0_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_2 <= io_Stationary_matrix_0_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_3 <= io_Stationary_matrix_0_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_4 <= io_Stationary_matrix_0_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_5 <= io_Stationary_matrix_0_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_6 <= io_Stationary_matrix_0_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_7 <= io_Stationary_matrix_0_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_0 <= io_Stationary_matrix_1_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_1 <= io_Stationary_matrix_1_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_2 <= io_Stationary_matrix_1_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_3 <= io_Stationary_matrix_1_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_4 <= io_Stationary_matrix_1_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_5 <= io_Stationary_matrix_1_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_6 <= io_Stationary_matrix_1_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_7 <= io_Stationary_matrix_1_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_0 <= io_Stationary_matrix_2_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_1 <= io_Stationary_matrix_2_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_2 <= io_Stationary_matrix_2_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_3 <= io_Stationary_matrix_2_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_4 <= io_Stationary_matrix_2_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_5 <= io_Stationary_matrix_2_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_6 <= io_Stationary_matrix_2_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_7 <= io_Stationary_matrix_2_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_0 <= io_Stationary_matrix_3_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_1 <= io_Stationary_matrix_3_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_2 <= io_Stationary_matrix_3_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_3 <= io_Stationary_matrix_3_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_4 <= io_Stationary_matrix_3_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_5 <= io_Stationary_matrix_3_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_6 <= io_Stationary_matrix_3_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_7 <= io_Stationary_matrix_3_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_0 <= io_Stationary_matrix_4_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_1 <= io_Stationary_matrix_4_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_2 <= io_Stationary_matrix_4_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_3 <= io_Stationary_matrix_4_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_4 <= io_Stationary_matrix_4_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_5 <= io_Stationary_matrix_4_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_6 <= io_Stationary_matrix_4_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_7 <= io_Stationary_matrix_4_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_0 <= io_Stationary_matrix_5_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_1 <= io_Stationary_matrix_5_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_2 <= io_Stationary_matrix_5_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_3 <= io_Stationary_matrix_5_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_4 <= io_Stationary_matrix_5_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_5 <= io_Stationary_matrix_5_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_6 <= io_Stationary_matrix_5_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_7 <= io_Stationary_matrix_5_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_0 <= io_Stationary_matrix_6_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_1 <= io_Stationary_matrix_6_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_2 <= io_Stationary_matrix_6_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_3 <= io_Stationary_matrix_6_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_4 <= io_Stationary_matrix_6_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_5 <= io_Stationary_matrix_6_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_6 <= io_Stationary_matrix_6_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_7 <= io_Stationary_matrix_6_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_0 <= io_Stationary_matrix_7_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_1 <= io_Stationary_matrix_7_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_2 <= io_Stationary_matrix_7_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_3 <= io_Stationary_matrix_7_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_4 <= io_Stationary_matrix_7_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_5 <= io_Stationary_matrix_7_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_6 <= io_Stationary_matrix_7_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_7 <= io_Stationary_matrix_7_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_0 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_0 <= count_0; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_1 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_1 <= count_1; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_2 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_2 <= count_2; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_3 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_3 <= count_3; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_4 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_4 <= count_4; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_5 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_5 <= count_5; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_6 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_6 <= count_6; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_7 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_7 <= count_7; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_8 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_8 <= 32'h0; // @[ivncontrol4.scala 87:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_9 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_9 <= 32'h0; // @[ivncontrol4.scala 87:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_10 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_10 <= 32'h0; // @[ivncontrol4.scala 87:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_11 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_11 <= 32'h0; // @[ivncontrol4.scala 87:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_12 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_12 <= 32'h0; // @[ivncontrol4.scala 87:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_13 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_13 <= 32'h0; // @[ivncontrol4.scala 87:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_14 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_14 <= 32'h0; // @[ivncontrol4.scala 87:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_15 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end
    if (reset) begin // @[ivncontrol4.scala 37:22]
      pin <= 32'h0; // @[ivncontrol4.scala 37:22]
    end else if (_T_72 & rowcount_6 == 32'h0 & rowcount_7 != 32'h0) begin // @[ivncontrol4.scala 183:192]
      pin <= 32'h7; // @[ivncontrol4.scala 184:13]
    end else if (_T_59 & rowcount_5 == 32'h0 & rowcount_6 != 32'h0) begin // @[ivncontrol4.scala 180:169]
      pin <= 32'h6; // @[ivncontrol4.scala 181:13]
    end else if (_T_48 & rowcount_4 == 32'h0 & rowcount_5 != 32'h0) begin // @[ivncontrol4.scala 177:146]
      pin <= 32'h5; // @[ivncontrol4.scala 178:13]
    end else begin
      pin <= _GEN_317;
    end
    if (reset) begin // @[ivncontrol4.scala 41:20]
      i <= 32'h0; // @[ivncontrol4.scala 41:20]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
        i <= _GEN_247;
      end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
        i <= _GEN_247;
      end else begin
        i <= _GEN_265;
      end
    end
    if (reset) begin // @[ivncontrol4.scala 42:20]
      j <= 32'h0; // @[ivncontrol4.scala 42:20]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
        j <= 32'h8; // @[ivncontrol4.scala 116:11]
      end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
        j <= _j_T_1; // @[ivncontrol4.scala 118:11]
      end else begin
        j <= {{28'd0}, _GEN_264};
      end
    end
    if (3'h0 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h0 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h0 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h0 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h0 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h0 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h0 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h0 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_0 <= _GEN_224;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_0 <= _GEN_224;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h0 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_0 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_0 <= _GEN_224;
      end
    end else begin
      count_0 <= _GEN_224;
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_1 <= _GEN_225;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_1 <= _GEN_225;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h1 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_1 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_1 <= _GEN_225;
      end
    end else begin
      count_1 <= _GEN_225;
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_2 <= _GEN_226;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_2 <= _GEN_226;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h2 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_2 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_2 <= _GEN_226;
      end
    end else begin
      count_2 <= _GEN_226;
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_3 <= _GEN_227;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_3 <= _GEN_227;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h3 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_3 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_3 <= _GEN_227;
      end
    end else begin
      count_3 <= _GEN_227;
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_4 <= _GEN_228;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_4 <= _GEN_228;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h4 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_4 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_4 <= _GEN_228;
      end
    end else begin
      count_4 <= _GEN_228;
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_5 <= _GEN_229;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_5 <= _GEN_229;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h5 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_5 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_5 <= _GEN_229;
      end
    end else begin
      count_5 <= _GEN_229;
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_6 <= _GEN_230;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_6 <= _GEN_230;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h6 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_6 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_6 <= _GEN_230;
      end
    end else begin
      count_6 <= _GEN_230;
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_7 <= _GEN_231;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_7 <= _GEN_231;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h7 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_7 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_7 <= _GEN_231;
      end
    end else begin
      count_7 <= _GEN_231;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  i_vn_0 = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  i_vn_1 = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  i_vn_2 = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  i_vn_3 = _RAND_3[4:0];
  _RAND_4 = {1{`RANDOM}};
  i_vn2_0 = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  i_vn2_1 = _RAND_5[4:0];
  _RAND_6 = {1{`RANDOM}};
  i_vn2_2 = _RAND_6[4:0];
  _RAND_7 = {1{`RANDOM}};
  i_vn2_3 = _RAND_7[4:0];
  _RAND_8 = {1{`RANDOM}};
  solution_0_0 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  solution_0_1 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  solution_0_2 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  solution_0_3 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  solution_0_4 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  solution_0_5 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  solution_0_6 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  solution_0_7 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  solution_1_0 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  solution_1_1 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  solution_1_2 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  solution_1_3 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  solution_1_4 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  solution_1_5 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  solution_1_6 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  solution_1_7 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  solution_2_0 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  solution_2_1 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  solution_2_2 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  solution_2_3 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  solution_2_4 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  solution_2_5 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  solution_2_6 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  solution_2_7 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  solution_3_0 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  solution_3_1 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  solution_3_2 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  solution_3_3 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  solution_3_4 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  solution_3_5 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  solution_3_6 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  solution_3_7 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  solution_4_0 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  solution_4_1 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  solution_4_2 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  solution_4_3 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  solution_4_4 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  solution_4_5 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  solution_4_6 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  solution_4_7 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  solution_5_0 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  solution_5_1 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  solution_5_2 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  solution_5_3 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  solution_5_4 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  solution_5_5 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  solution_5_6 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  solution_5_7 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  solution_6_0 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  solution_6_1 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  solution_6_2 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  solution_6_3 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  solution_6_4 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  solution_6_5 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  solution_6_6 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  solution_6_7 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  solution_7_0 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  solution_7_1 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  solution_7_2 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  solution_7_3 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  solution_7_4 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  solution_7_5 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  solution_7_6 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  solution_7_7 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  rowcount_0 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  rowcount_1 = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  rowcount_2 = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  rowcount_3 = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  rowcount_4 = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  rowcount_5 = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  rowcount_6 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  rowcount_7 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  rowcount_8 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  rowcount_9 = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  rowcount_10 = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  rowcount_11 = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  rowcount_12 = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  rowcount_13 = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  rowcount_14 = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  rowcount_15 = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  pin = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  i = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  j = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  mat_0_0 = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  mat_0_1 = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  mat_0_2 = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  mat_0_3 = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  mat_0_4 = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  mat_0_5 = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  mat_0_6 = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  mat_0_7 = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  mat_1_0 = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  mat_1_1 = _RAND_100[31:0];
  _RAND_101 = {1{`RANDOM}};
  mat_1_2 = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  mat_1_3 = _RAND_102[31:0];
  _RAND_103 = {1{`RANDOM}};
  mat_1_4 = _RAND_103[31:0];
  _RAND_104 = {1{`RANDOM}};
  mat_1_5 = _RAND_104[31:0];
  _RAND_105 = {1{`RANDOM}};
  mat_1_6 = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  mat_1_7 = _RAND_106[31:0];
  _RAND_107 = {1{`RANDOM}};
  mat_2_0 = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  mat_2_1 = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  mat_2_2 = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  mat_2_3 = _RAND_110[31:0];
  _RAND_111 = {1{`RANDOM}};
  mat_2_4 = _RAND_111[31:0];
  _RAND_112 = {1{`RANDOM}};
  mat_2_5 = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  mat_2_6 = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  mat_2_7 = _RAND_114[31:0];
  _RAND_115 = {1{`RANDOM}};
  mat_3_0 = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  mat_3_1 = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  mat_3_2 = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  mat_3_3 = _RAND_118[31:0];
  _RAND_119 = {1{`RANDOM}};
  mat_3_4 = _RAND_119[31:0];
  _RAND_120 = {1{`RANDOM}};
  mat_3_5 = _RAND_120[31:0];
  _RAND_121 = {1{`RANDOM}};
  mat_3_6 = _RAND_121[31:0];
  _RAND_122 = {1{`RANDOM}};
  mat_3_7 = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  mat_4_0 = _RAND_123[31:0];
  _RAND_124 = {1{`RANDOM}};
  mat_4_1 = _RAND_124[31:0];
  _RAND_125 = {1{`RANDOM}};
  mat_4_2 = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  mat_4_3 = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  mat_4_4 = _RAND_127[31:0];
  _RAND_128 = {1{`RANDOM}};
  mat_4_5 = _RAND_128[31:0];
  _RAND_129 = {1{`RANDOM}};
  mat_4_6 = _RAND_129[31:0];
  _RAND_130 = {1{`RANDOM}};
  mat_4_7 = _RAND_130[31:0];
  _RAND_131 = {1{`RANDOM}};
  mat_5_0 = _RAND_131[31:0];
  _RAND_132 = {1{`RANDOM}};
  mat_5_1 = _RAND_132[31:0];
  _RAND_133 = {1{`RANDOM}};
  mat_5_2 = _RAND_133[31:0];
  _RAND_134 = {1{`RANDOM}};
  mat_5_3 = _RAND_134[31:0];
  _RAND_135 = {1{`RANDOM}};
  mat_5_4 = _RAND_135[31:0];
  _RAND_136 = {1{`RANDOM}};
  mat_5_5 = _RAND_136[31:0];
  _RAND_137 = {1{`RANDOM}};
  mat_5_6 = _RAND_137[31:0];
  _RAND_138 = {1{`RANDOM}};
  mat_5_7 = _RAND_138[31:0];
  _RAND_139 = {1{`RANDOM}};
  mat_6_0 = _RAND_139[31:0];
  _RAND_140 = {1{`RANDOM}};
  mat_6_1 = _RAND_140[31:0];
  _RAND_141 = {1{`RANDOM}};
  mat_6_2 = _RAND_141[31:0];
  _RAND_142 = {1{`RANDOM}};
  mat_6_3 = _RAND_142[31:0];
  _RAND_143 = {1{`RANDOM}};
  mat_6_4 = _RAND_143[31:0];
  _RAND_144 = {1{`RANDOM}};
  mat_6_5 = _RAND_144[31:0];
  _RAND_145 = {1{`RANDOM}};
  mat_6_6 = _RAND_145[31:0];
  _RAND_146 = {1{`RANDOM}};
  mat_6_7 = _RAND_146[31:0];
  _RAND_147 = {1{`RANDOM}};
  mat_7_0 = _RAND_147[31:0];
  _RAND_148 = {1{`RANDOM}};
  mat_7_1 = _RAND_148[31:0];
  _RAND_149 = {1{`RANDOM}};
  mat_7_2 = _RAND_149[31:0];
  _RAND_150 = {1{`RANDOM}};
  mat_7_3 = _RAND_150[31:0];
  _RAND_151 = {1{`RANDOM}};
  mat_7_4 = _RAND_151[31:0];
  _RAND_152 = {1{`RANDOM}};
  mat_7_5 = _RAND_152[31:0];
  _RAND_153 = {1{`RANDOM}};
  mat_7_6 = _RAND_153[31:0];
  _RAND_154 = {1{`RANDOM}};
  mat_7_7 = _RAND_154[31:0];
  _RAND_155 = {1{`RANDOM}};
  count_0 = _RAND_155[31:0];
  _RAND_156 = {1{`RANDOM}};
  count_1 = _RAND_156[31:0];
  _RAND_157 = {1{`RANDOM}};
  count_2 = _RAND_157[31:0];
  _RAND_158 = {1{`RANDOM}};
  count_3 = _RAND_158[31:0];
  _RAND_159 = {1{`RANDOM}};
  count_4 = _RAND_159[31:0];
  _RAND_160 = {1{`RANDOM}};
  count_5 = _RAND_160[31:0];
  _RAND_161 = {1{`RANDOM}};
  count_6 = _RAND_161[31:0];
  _RAND_162 = {1{`RANDOM}};
  count_7 = _RAND_162[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ivncontrol4_4(
  input         clock,
  input         reset,
  input  [15:0] io_Stationary_matrix_0_0,
  input  [15:0] io_Stationary_matrix_0_1,
  input  [15:0] io_Stationary_matrix_0_2,
  input  [15:0] io_Stationary_matrix_0_3,
  input  [15:0] io_Stationary_matrix_0_4,
  input  [15:0] io_Stationary_matrix_0_5,
  input  [15:0] io_Stationary_matrix_0_6,
  input  [15:0] io_Stationary_matrix_0_7,
  input  [15:0] io_Stationary_matrix_1_0,
  input  [15:0] io_Stationary_matrix_1_1,
  input  [15:0] io_Stationary_matrix_1_2,
  input  [15:0] io_Stationary_matrix_1_3,
  input  [15:0] io_Stationary_matrix_1_4,
  input  [15:0] io_Stationary_matrix_1_5,
  input  [15:0] io_Stationary_matrix_1_6,
  input  [15:0] io_Stationary_matrix_1_7,
  input  [15:0] io_Stationary_matrix_2_0,
  input  [15:0] io_Stationary_matrix_2_1,
  input  [15:0] io_Stationary_matrix_2_2,
  input  [15:0] io_Stationary_matrix_2_3,
  input  [15:0] io_Stationary_matrix_2_4,
  input  [15:0] io_Stationary_matrix_2_5,
  input  [15:0] io_Stationary_matrix_2_6,
  input  [15:0] io_Stationary_matrix_2_7,
  input  [15:0] io_Stationary_matrix_3_0,
  input  [15:0] io_Stationary_matrix_3_1,
  input  [15:0] io_Stationary_matrix_3_2,
  input  [15:0] io_Stationary_matrix_3_3,
  input  [15:0] io_Stationary_matrix_3_4,
  input  [15:0] io_Stationary_matrix_3_5,
  input  [15:0] io_Stationary_matrix_3_6,
  input  [15:0] io_Stationary_matrix_3_7,
  input  [15:0] io_Stationary_matrix_4_0,
  input  [15:0] io_Stationary_matrix_4_1,
  input  [15:0] io_Stationary_matrix_4_2,
  input  [15:0] io_Stationary_matrix_4_3,
  input  [15:0] io_Stationary_matrix_4_4,
  input  [15:0] io_Stationary_matrix_4_5,
  input  [15:0] io_Stationary_matrix_4_6,
  input  [15:0] io_Stationary_matrix_4_7,
  input  [15:0] io_Stationary_matrix_5_0,
  input  [15:0] io_Stationary_matrix_5_1,
  input  [15:0] io_Stationary_matrix_5_2,
  input  [15:0] io_Stationary_matrix_5_3,
  input  [15:0] io_Stationary_matrix_5_4,
  input  [15:0] io_Stationary_matrix_5_5,
  input  [15:0] io_Stationary_matrix_5_6,
  input  [15:0] io_Stationary_matrix_5_7,
  input  [15:0] io_Stationary_matrix_6_0,
  input  [15:0] io_Stationary_matrix_6_1,
  input  [15:0] io_Stationary_matrix_6_2,
  input  [15:0] io_Stationary_matrix_6_3,
  input  [15:0] io_Stationary_matrix_6_4,
  input  [15:0] io_Stationary_matrix_6_5,
  input  [15:0] io_Stationary_matrix_6_6,
  input  [15:0] io_Stationary_matrix_6_7,
  input  [15:0] io_Stationary_matrix_7_0,
  input  [15:0] io_Stationary_matrix_7_1,
  input  [15:0] io_Stationary_matrix_7_2,
  input  [15:0] io_Stationary_matrix_7_3,
  input  [15:0] io_Stationary_matrix_7_4,
  input  [15:0] io_Stationary_matrix_7_5,
  input  [15:0] io_Stationary_matrix_7_6,
  input  [15:0] io_Stationary_matrix_7_7,
  output [4:0]  io_o_vn_0,
  output [4:0]  io_o_vn_1,
  output [4:0]  io_o_vn_2,
  output [4:0]  io_o_vn_3,
  output [4:0]  io_o_vn2_0,
  output [4:0]  io_o_vn2_1,
  output [4:0]  io_o_vn2_2,
  output [4:0]  io_o_vn2_3,
  input         io_validpin
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
`endif // RANDOMIZE_REG_INIT
  reg [4:0] i_vn_0; // @[ivncontrol4.scala 17:23]
  reg [4:0] i_vn_1; // @[ivncontrol4.scala 17:23]
  reg [4:0] i_vn_2; // @[ivncontrol4.scala 17:23]
  reg [4:0] i_vn_3; // @[ivncontrol4.scala 17:23]
  reg [4:0] i_vn2_0; // @[ivncontrol4.scala 18:24]
  reg [4:0] i_vn2_1; // @[ivncontrol4.scala 18:24]
  reg [4:0] i_vn2_2; // @[ivncontrol4.scala 18:24]
  reg [4:0] i_vn2_3; // @[ivncontrol4.scala 18:24]
  reg [15:0] solution_0_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_0_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_0_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_0_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_0_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_0_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_0_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_0_7; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_7; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_7; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_7; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_7; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_7; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_7; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_7; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_0; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_1; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_2; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_3; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_4; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_5; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_6; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_7; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_8; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_9; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_10; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_11; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_12; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_13; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_14; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_15; // @[ivncontrol4.scala 27:27]
  reg [31:0] pin; // @[ivncontrol4.scala 37:22]
  reg [31:0] i; // @[ivncontrol4.scala 41:20]
  reg [31:0] j; // @[ivncontrol4.scala 42:20]
  wire  _io_ProcessValid_T = i == 32'h7; // @[ivncontrol4.scala 44:27]
  wire  _io_ProcessValid_T_1 = j == 32'h7; // @[ivncontrol4.scala 44:42]
  wire  _io_ProcessValid_T_2 = i == 32'h7 & j == 32'h7; // @[ivncontrol4.scala 44:36]
  reg [31:0] mat_0_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_0_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_0_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_0_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_0_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_0_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_0_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_0_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] count_0; // @[ivncontrol4.scala 58:20]
  reg [31:0] count_1; // @[ivncontrol4.scala 58:20]
  reg [31:0] count_2; // @[ivncontrol4.scala 58:20]
  reg [31:0] count_3; // @[ivncontrol4.scala 58:20]
  reg [31:0] count_4; // @[ivncontrol4.scala 58:20]
  reg [31:0] count_5; // @[ivncontrol4.scala 58:20]
  reg [31:0] count_6; // @[ivncontrol4.scala 58:20]
  reg [31:0] count_7; // @[ivncontrol4.scala 58:20]
  wire  _GEN_3825 = 3'h0 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_65 = 3'h0 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_0_1 : io_Stationary_matrix_0_0; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_66 = 3'h0 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_0_2 : _GEN_65; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_67 = 3'h0 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_0_3 : _GEN_66; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_68 = 3'h0 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_0_4 : _GEN_67; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_69 = 3'h0 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_0_5 : _GEN_68; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_70 = 3'h0 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_0_6 : _GEN_69; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_71 = 3'h0 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_0_7 : _GEN_70; // @[ivncontrol4.scala 63:{17,17}]
  wire  _GEN_3839 = 3'h1 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_72 = 3'h1 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_1_0 : _GEN_71; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_73 = 3'h1 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_1_1 : _GEN_72; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_74 = 3'h1 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_1_2 : _GEN_73; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_75 = 3'h1 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_1_3 : _GEN_74; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_76 = 3'h1 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_1_4 : _GEN_75; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_77 = 3'h1 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_1_5 : _GEN_76; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_78 = 3'h1 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_1_6 : _GEN_77; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_79 = 3'h1 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_1_7 : _GEN_78; // @[ivncontrol4.scala 63:{17,17}]
  wire  _GEN_3855 = 3'h2 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_80 = 3'h2 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_2_0 : _GEN_79; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_81 = 3'h2 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_2_1 : _GEN_80; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_82 = 3'h2 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_2_2 : _GEN_81; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_83 = 3'h2 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_2_3 : _GEN_82; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_84 = 3'h2 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_2_4 : _GEN_83; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_85 = 3'h2 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_2_5 : _GEN_84; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_86 = 3'h2 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_2_6 : _GEN_85; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_87 = 3'h2 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_2_7 : _GEN_86; // @[ivncontrol4.scala 63:{17,17}]
  wire  _GEN_3871 = 3'h3 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_88 = 3'h3 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_3_0 : _GEN_87; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_89 = 3'h3 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_3_1 : _GEN_88; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_90 = 3'h3 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_3_2 : _GEN_89; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_91 = 3'h3 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_3_3 : _GEN_90; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_92 = 3'h3 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_3_4 : _GEN_91; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_93 = 3'h3 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_3_5 : _GEN_92; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_94 = 3'h3 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_3_6 : _GEN_93; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_95 = 3'h3 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_3_7 : _GEN_94; // @[ivncontrol4.scala 63:{17,17}]
  wire  _GEN_3887 = 3'h4 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_96 = 3'h4 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_4_0 : _GEN_95; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_97 = 3'h4 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_4_1 : _GEN_96; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_98 = 3'h4 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_4_2 : _GEN_97; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_99 = 3'h4 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_4_3 : _GEN_98; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_100 = 3'h4 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_4_4 : _GEN_99; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_101 = 3'h4 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_4_5 : _GEN_100; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_102 = 3'h4 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_4_6 : _GEN_101; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_103 = 3'h4 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_4_7 : _GEN_102; // @[ivncontrol4.scala 63:{17,17}]
  wire  _GEN_3903 = 3'h5 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_104 = 3'h5 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_5_0 : _GEN_103; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_105 = 3'h5 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_5_1 : _GEN_104; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_106 = 3'h5 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_5_2 : _GEN_105; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_107 = 3'h5 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_5_3 : _GEN_106; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_108 = 3'h5 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_5_4 : _GEN_107; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_109 = 3'h5 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_5_5 : _GEN_108; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_110 = 3'h5 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_5_6 : _GEN_109; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_111 = 3'h5 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_5_7 : _GEN_110; // @[ivncontrol4.scala 63:{17,17}]
  wire  _GEN_3919 = 3'h6 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_112 = 3'h6 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_6_0 : _GEN_111; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_113 = 3'h6 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_6_1 : _GEN_112; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_114 = 3'h6 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_6_2 : _GEN_113; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_115 = 3'h6 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_6_3 : _GEN_114; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_116 = 3'h6 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_6_4 : _GEN_115; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_117 = 3'h6 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_6_5 : _GEN_116; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_118 = 3'h6 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_6_6 : _GEN_117; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_119 = 3'h6 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_6_7 : _GEN_118; // @[ivncontrol4.scala 63:{17,17}]
  wire  _GEN_3935 = 3'h7 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_120 = 3'h7 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_7_0 : _GEN_119; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_121 = 3'h7 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_7_1 : _GEN_120; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_122 = 3'h7 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_7_2 : _GEN_121; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_123 = 3'h7 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_7_3 : _GEN_122; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_124 = 3'h7 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_7_4 : _GEN_123; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_125 = 3'h7 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_7_5 : _GEN_124; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_126 = 3'h7 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_7_6 : _GEN_125; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_127 = 3'h7 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_7_7 : _GEN_126; // @[ivncontrol4.scala 63:{17,17}]
  wire [31:0] _mat_T_1_T_2 = {{16'd0}, _GEN_127}; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_129 = _GEN_3825 & 4'h1 == j[3:0] ? solution_0_1 : solution_0_0; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_130 = _GEN_3825 & 4'h2 == j[3:0] ? solution_0_2 : _GEN_129; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_131 = _GEN_3825 & 4'h3 == j[3:0] ? solution_0_3 : _GEN_130; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_132 = _GEN_3825 & 4'h4 == j[3:0] ? solution_0_4 : _GEN_131; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_133 = _GEN_3825 & 4'h5 == j[3:0] ? solution_0_5 : _GEN_132; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_134 = _GEN_3825 & 4'h6 == j[3:0] ? solution_0_6 : _GEN_133; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_135 = _GEN_3825 & 4'h7 == j[3:0] ? solution_0_7 : _GEN_134; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_136 = _GEN_3825 & 4'h8 == j[3:0] ? 16'h0 : _GEN_135; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_137 = _GEN_3839 & 4'h0 == j[3:0] ? solution_1_0 : _GEN_136; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_138 = _GEN_3839 & 4'h1 == j[3:0] ? solution_1_1 : _GEN_137; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_139 = _GEN_3839 & 4'h2 == j[3:0] ? solution_1_2 : _GEN_138; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_140 = _GEN_3839 & 4'h3 == j[3:0] ? solution_1_3 : _GEN_139; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_141 = _GEN_3839 & 4'h4 == j[3:0] ? solution_1_4 : _GEN_140; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_142 = _GEN_3839 & 4'h5 == j[3:0] ? solution_1_5 : _GEN_141; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_143 = _GEN_3839 & 4'h6 == j[3:0] ? solution_1_6 : _GEN_142; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_144 = _GEN_3839 & 4'h7 == j[3:0] ? solution_1_7 : _GEN_143; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_145 = _GEN_3839 & 4'h8 == j[3:0] ? 16'h0 : _GEN_144; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_146 = _GEN_3855 & 4'h0 == j[3:0] ? solution_2_0 : _GEN_145; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_147 = _GEN_3855 & 4'h1 == j[3:0] ? solution_2_1 : _GEN_146; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_148 = _GEN_3855 & 4'h2 == j[3:0] ? solution_2_2 : _GEN_147; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_149 = _GEN_3855 & 4'h3 == j[3:0] ? solution_2_3 : _GEN_148; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_150 = _GEN_3855 & 4'h4 == j[3:0] ? solution_2_4 : _GEN_149; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_151 = _GEN_3855 & 4'h5 == j[3:0] ? solution_2_5 : _GEN_150; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_152 = _GEN_3855 & 4'h6 == j[3:0] ? solution_2_6 : _GEN_151; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_153 = _GEN_3855 & 4'h7 == j[3:0] ? solution_2_7 : _GEN_152; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_154 = _GEN_3855 & 4'h8 == j[3:0] ? 16'h0 : _GEN_153; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_155 = _GEN_3871 & 4'h0 == j[3:0] ? solution_3_0 : _GEN_154; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_156 = _GEN_3871 & 4'h1 == j[3:0] ? solution_3_1 : _GEN_155; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_157 = _GEN_3871 & 4'h2 == j[3:0] ? solution_3_2 : _GEN_156; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_158 = _GEN_3871 & 4'h3 == j[3:0] ? solution_3_3 : _GEN_157; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_159 = _GEN_3871 & 4'h4 == j[3:0] ? solution_3_4 : _GEN_158; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_160 = _GEN_3871 & 4'h5 == j[3:0] ? solution_3_5 : _GEN_159; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_161 = _GEN_3871 & 4'h6 == j[3:0] ? solution_3_6 : _GEN_160; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_162 = _GEN_3871 & 4'h7 == j[3:0] ? solution_3_7 : _GEN_161; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_163 = _GEN_3871 & 4'h8 == j[3:0] ? 16'h0 : _GEN_162; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_164 = _GEN_3887 & 4'h0 == j[3:0] ? solution_4_0 : _GEN_163; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_165 = _GEN_3887 & 4'h1 == j[3:0] ? solution_4_1 : _GEN_164; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_166 = _GEN_3887 & 4'h2 == j[3:0] ? solution_4_2 : _GEN_165; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_167 = _GEN_3887 & 4'h3 == j[3:0] ? solution_4_3 : _GEN_166; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_168 = _GEN_3887 & 4'h4 == j[3:0] ? solution_4_4 : _GEN_167; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_169 = _GEN_3887 & 4'h5 == j[3:0] ? solution_4_5 : _GEN_168; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_170 = _GEN_3887 & 4'h6 == j[3:0] ? solution_4_6 : _GEN_169; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_171 = _GEN_3887 & 4'h7 == j[3:0] ? solution_4_7 : _GEN_170; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_172 = _GEN_3887 & 4'h8 == j[3:0] ? 16'h0 : _GEN_171; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_173 = _GEN_3903 & 4'h0 == j[3:0] ? solution_5_0 : _GEN_172; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_174 = _GEN_3903 & 4'h1 == j[3:0] ? solution_5_1 : _GEN_173; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_175 = _GEN_3903 & 4'h2 == j[3:0] ? solution_5_2 : _GEN_174; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_176 = _GEN_3903 & 4'h3 == j[3:0] ? solution_5_3 : _GEN_175; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_177 = _GEN_3903 & 4'h4 == j[3:0] ? solution_5_4 : _GEN_176; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_178 = _GEN_3903 & 4'h5 == j[3:0] ? solution_5_5 : _GEN_177; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_179 = _GEN_3903 & 4'h6 == j[3:0] ? solution_5_6 : _GEN_178; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_180 = _GEN_3903 & 4'h7 == j[3:0] ? solution_5_7 : _GEN_179; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_181 = _GEN_3903 & 4'h8 == j[3:0] ? 16'h0 : _GEN_180; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_182 = _GEN_3919 & 4'h0 == j[3:0] ? solution_6_0 : _GEN_181; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_183 = _GEN_3919 & 4'h1 == j[3:0] ? solution_6_1 : _GEN_182; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_184 = _GEN_3919 & 4'h2 == j[3:0] ? solution_6_2 : _GEN_183; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_185 = _GEN_3919 & 4'h3 == j[3:0] ? solution_6_3 : _GEN_184; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_186 = _GEN_3919 & 4'h4 == j[3:0] ? solution_6_4 : _GEN_185; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_187 = _GEN_3919 & 4'h5 == j[3:0] ? solution_6_5 : _GEN_186; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_188 = _GEN_3919 & 4'h6 == j[3:0] ? solution_6_6 : _GEN_187; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_189 = _GEN_3919 & 4'h7 == j[3:0] ? solution_6_7 : _GEN_188; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_190 = _GEN_3919 & 4'h8 == j[3:0] ? 16'h0 : _GEN_189; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_191 = _GEN_3935 & 4'h0 == j[3:0] ? solution_7_0 : _GEN_190; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_192 = _GEN_3935 & 4'h1 == j[3:0] ? solution_7_1 : _GEN_191; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_193 = _GEN_3935 & 4'h2 == j[3:0] ? solution_7_2 : _GEN_192; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_194 = _GEN_3935 & 4'h3 == j[3:0] ? solution_7_3 : _GEN_193; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_195 = _GEN_3935 & 4'h4 == j[3:0] ? solution_7_4 : _GEN_194; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_196 = _GEN_3935 & 4'h5 == j[3:0] ? solution_7_5 : _GEN_195; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_197 = _GEN_3935 & 4'h6 == j[3:0] ? solution_7_6 : _GEN_196; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_198 = _GEN_3935 & 4'h7 == j[3:0] ? solution_7_7 : _GEN_197; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_199 = _GEN_3935 & 4'h8 == j[3:0] ? 16'h0 : _GEN_198; // @[ivncontrol4.scala 65:{31,31}]
  wire [31:0] _GEN_201 = 3'h1 == i[2:0] ? count_1 : count_0; // @[ivncontrol4.scala 66:{33,33}]
  wire [31:0] _GEN_202 = 3'h2 == i[2:0] ? count_2 : _GEN_201; // @[ivncontrol4.scala 66:{33,33}]
  wire [31:0] _GEN_203 = 3'h3 == i[2:0] ? count_3 : _GEN_202; // @[ivncontrol4.scala 66:{33,33}]
  wire [31:0] _GEN_204 = 3'h4 == i[2:0] ? count_4 : _GEN_203; // @[ivncontrol4.scala 66:{33,33}]
  wire [31:0] _GEN_205 = 3'h5 == i[2:0] ? count_5 : _GEN_204; // @[ivncontrol4.scala 66:{33,33}]
  wire [31:0] _GEN_206 = 3'h6 == i[2:0] ? count_6 : _GEN_205; // @[ivncontrol4.scala 66:{33,33}]
  wire [31:0] _GEN_207 = 3'h7 == i[2:0] ? count_7 : _GEN_206; // @[ivncontrol4.scala 66:{33,33}]
  wire [31:0] _count_T_2 = _GEN_207 + 32'h1; // @[ivncontrol4.scala 66:33]
  wire [31:0] _GEN_208 = 3'h0 == i[2:0] ? _count_T_2 : count_0; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_209 = 3'h1 == i[2:0] ? _count_T_2 : count_1; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_210 = 3'h2 == i[2:0] ? _count_T_2 : count_2; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_211 = 3'h3 == i[2:0] ? _count_T_2 : count_3; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_212 = 3'h4 == i[2:0] ? _count_T_2 : count_4; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_213 = 3'h5 == i[2:0] ? _count_T_2 : count_5; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_214 = 3'h6 == i[2:0] ? _count_T_2 : count_6; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_215 = 3'h7 == i[2:0] ? _count_T_2 : count_7; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_216 = _GEN_199 != 16'h0 ? _GEN_208 : count_0; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_217 = _GEN_199 != 16'h0 ? _GEN_209 : count_1; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_218 = _GEN_199 != 16'h0 ? _GEN_210 : count_2; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_219 = _GEN_199 != 16'h0 ? _GEN_211 : count_3; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_220 = _GEN_199 != 16'h0 ? _GEN_212 : count_4; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_221 = _GEN_199 != 16'h0 ? _GEN_213 : count_5; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_222 = _GEN_199 != 16'h0 ? _GEN_214 : count_6; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_223 = _GEN_199 != 16'h0 ? _GEN_215 : count_7; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_224 = io_validpin ? _GEN_216 : count_0; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _GEN_225 = io_validpin ? _GEN_217 : count_1; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _GEN_226 = io_validpin ? _GEN_218 : count_2; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _GEN_227 = io_validpin ? _GEN_219 : count_3; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _GEN_228 = io_validpin ? _GEN_220 : count_4; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _GEN_229 = io_validpin ? _GEN_221 : count_5; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _GEN_230 = io_validpin ? _GEN_222 : count_6; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _GEN_231 = io_validpin ? _GEN_223 : count_7; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _i_T_1 = i + 32'h1; // @[ivncontrol4.scala 113:16]
  wire [31:0] _GEN_247 = i < 32'h7 & _io_ProcessValid_T_1 ? _i_T_1 : i; // @[ivncontrol4.scala 112:74 113:11 41:20]
  wire [31:0] _j_T_1 = j + 32'h1; // @[ivncontrol4.scala 118:16]
  wire [3:0] _GEN_264 = _io_ProcessValid_T & j == 32'h8 ? 4'h8 : 4'h0; // @[ivncontrol4.scala 120:77 121:11 129:11]
  wire [31:0] _GEN_265 = _io_ProcessValid_T & j == 32'h8 ? 32'h7 : _GEN_247; // @[ivncontrol4.scala 120:77 122:11]
  wire  _GEN_312 = _io_ProcessValid_T_2; // @[ivncontrol4.scala 153:41]
  wire [31:0] _GEN_313 = rowcount_0 != 32'h0 ? 32'h0 : pin; // @[ivncontrol4.scala 162:30 163:13 37:22]
  wire  _T_27 = rowcount_0 == 32'h0; // @[ivncontrol4.scala 165:23]
  wire [31:0] _GEN_314 = rowcount_0 == 32'h0 & rowcount_1 != 32'h0 ? 32'h1 : _GEN_313; // @[ivncontrol4.scala 165:54 166:13]
  wire  _T_32 = _T_27 & rowcount_1 == 32'h0; // @[ivncontrol4.scala 168:31]
  wire [31:0] _GEN_315 = _T_27 & rowcount_1 == 32'h0 & rowcount_2 != 32'h0 ? 32'h2 : _GEN_314; // @[ivncontrol4.scala 168:77 169:13]
  wire  _T_39 = _T_32 & rowcount_2 == 32'h0; // @[ivncontrol4.scala 171:54]
  wire [31:0] _GEN_316 = _T_32 & rowcount_2 == 32'h0 & rowcount_3 != 32'h0 ? 32'h3 : _GEN_315; // @[ivncontrol4.scala 171:100 172:13]
  wire  _T_48 = _T_39 & rowcount_3 == 32'h0; // @[ivncontrol4.scala 174:77]
  wire [31:0] _GEN_317 = _T_39 & rowcount_3 == 32'h0 & rowcount_4 != 32'h0 ? 32'h4 : _GEN_316; // @[ivncontrol4.scala 174:123 175:13]
  wire  _T_59 = _T_48 & rowcount_4 == 32'h0; // @[ivncontrol4.scala 177:100]
  wire  _T_72 = _T_59 & rowcount_5 == 32'h0; // @[ivncontrol4.scala 180:123]
  wire  valid = _io_ProcessValid_T_2; // @[ivncontrol4.scala 153:41]
  wire [32:0] _T_91 = {{1'd0}, pin}; // @[ivncontrol4.scala 191:27]
  wire [31:0] _GEN_322 = 4'h1 == _T_91[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_323 = 4'h2 == _T_91[3:0] ? rowcount_2 : _GEN_322; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_324 = 4'h3 == _T_91[3:0] ? rowcount_3 : _GEN_323; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_325 = 4'h4 == _T_91[3:0] ? rowcount_4 : _GEN_324; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_326 = 4'h5 == _T_91[3:0] ? rowcount_5 : _GEN_325; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_327 = 4'h6 == _T_91[3:0] ? rowcount_6 : _GEN_326; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_328 = 4'h7 == _T_91[3:0] ? rowcount_7 : _GEN_327; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_329 = 4'h8 == _T_91[3:0] ? rowcount_8 : _GEN_328; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_330 = 4'h9 == _T_91[3:0] ? rowcount_9 : _GEN_329; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_331 = 4'ha == _T_91[3:0] ? rowcount_10 : _GEN_330; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_332 = 4'hb == _T_91[3:0] ? rowcount_11 : _GEN_331; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_333 = 4'hc == _T_91[3:0] ? rowcount_12 : _GEN_332; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_334 = 4'hd == _T_91[3:0] ? rowcount_13 : _GEN_333; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_335 = 4'he == _T_91[3:0] ? rowcount_14 : _GEN_334; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_336 = 4'hf == _T_91[3:0] ? rowcount_15 : _GEN_335; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_449 = _GEN_336 == 32'h1 ? _T_91[31:0] : 32'h3; // @[ivncontrol4.scala 142:17 241:50 242:21]
  wire [31:0] _GEN_450 = _GEN_336 == 32'h2 ? _T_91[31:0] : _GEN_449; // @[ivncontrol4.scala 237:51 238:21]
  wire [31:0] _GEN_451 = _GEN_336 == 32'h2 ? _T_91[31:0] : 32'h1; // @[ivncontrol4.scala 142:17 237:51 239:21]
  wire [31:0] _GEN_452 = _GEN_336 == 32'h3 ? _T_91[31:0] : _GEN_450; // @[ivncontrol4.scala 232:50 233:21]
  wire [31:0] _GEN_453 = _GEN_336 == 32'h3 ? _T_91[31:0] : _GEN_451; // @[ivncontrol4.scala 232:50 234:21]
  wire [31:0] _GEN_454 = _GEN_336 == 32'h3 ? _T_91[31:0] : 32'h19; // @[ivncontrol4.scala 142:17 232:50 235:21]
  wire [31:0] _GEN_455 = _GEN_336 == 32'h4 ? _T_91[31:0] : _GEN_452; // @[ivncontrol4.scala 224:50 225:21]
  wire [31:0] _GEN_456 = _GEN_336 == 32'h4 ? _T_91[31:0] : _GEN_453; // @[ivncontrol4.scala 224:50 226:21]
  wire [31:0] _GEN_457 = _GEN_336 == 32'h4 ? _T_91[31:0] : _GEN_454; // @[ivncontrol4.scala 224:50 227:21]
  wire [31:0] _GEN_458 = _GEN_336 == 32'h4 ? _T_91[31:0] : 32'hf; // @[ivncontrol4.scala 142:17 224:50 228:21]
  wire [31:0] _GEN_459 = _GEN_336 == 32'h5 ? _T_91[31:0] : _GEN_455; // @[ivncontrol4.scala 217:50 218:21]
  wire [31:0] _GEN_460 = _GEN_336 == 32'h5 ? _T_91[31:0] : _GEN_456; // @[ivncontrol4.scala 217:50 219:21]
  wire [31:0] _GEN_461 = _GEN_336 == 32'h5 ? _T_91[31:0] : _GEN_457; // @[ivncontrol4.scala 217:50 220:21]
  wire [31:0] _GEN_462 = _GEN_336 == 32'h5 ? _T_91[31:0] : _GEN_458; // @[ivncontrol4.scala 217:50 221:21]
  wire [31:0] _GEN_463 = _GEN_336 == 32'h5 ? _T_91[31:0] : 32'h10; // @[ivncontrol4.scala 143:18 217:50 222:22]
  wire [31:0] _GEN_464 = _GEN_336 == 32'h6 ? _T_91[31:0] : _GEN_459; // @[ivncontrol4.scala 209:52 210:21]
  wire [31:0] _GEN_465 = _GEN_336 == 32'h6 ? _T_91[31:0] : _GEN_460; // @[ivncontrol4.scala 209:52 211:21]
  wire [31:0] _GEN_466 = _GEN_336 == 32'h6 ? _T_91[31:0] : _GEN_461; // @[ivncontrol4.scala 209:52 212:21]
  wire [31:0] _GEN_467 = _GEN_336 == 32'h6 ? _T_91[31:0] : _GEN_462; // @[ivncontrol4.scala 209:52 213:21]
  wire [31:0] _GEN_468 = _GEN_336 == 32'h6 ? _T_91[31:0] : _GEN_463; // @[ivncontrol4.scala 209:52 214:22]
  wire [31:0] _GEN_469 = _GEN_336 == 32'h6 ? _T_91[31:0] : 32'h4; // @[ivncontrol4.scala 143:18 209:52 215:22]
  wire [31:0] _GEN_470 = _GEN_336 == 32'h7 ? _T_91[31:0] : _GEN_464; // @[ivncontrol4.scala 201:52 202:21]
  wire [31:0] _GEN_471 = _GEN_336 == 32'h7 ? _T_91[31:0] : _GEN_465; // @[ivncontrol4.scala 201:52 203:21]
  wire [31:0] _GEN_472 = _GEN_336 == 32'h7 ? _T_91[31:0] : _GEN_466; // @[ivncontrol4.scala 201:52 204:21]
  wire [31:0] _GEN_473 = _GEN_336 == 32'h7 ? _T_91[31:0] : _GEN_467; // @[ivncontrol4.scala 201:52 205:21]
  wire [31:0] _GEN_474 = _GEN_336 == 32'h7 ? _T_91[31:0] : _GEN_468; // @[ivncontrol4.scala 201:52 206:22]
  wire [31:0] _GEN_475 = _GEN_336 == 32'h7 ? _T_91[31:0] : _GEN_469; // @[ivncontrol4.scala 201:52 207:22]
  wire [31:0] _GEN_476 = _GEN_336 == 32'h7 ? _T_91[31:0] : 32'h12; // @[ivncontrol4.scala 143:18 201:52 208:22]
  wire [31:0] _GEN_477 = _GEN_336 >= 32'h8 ? _T_91[31:0] : _GEN_470; // @[ivncontrol4.scala 191:42 192:21]
  wire [31:0] _GEN_478 = _GEN_336 >= 32'h8 ? _T_91[31:0] : _GEN_471; // @[ivncontrol4.scala 191:42 193:21]
  wire [31:0] _GEN_479 = _GEN_336 >= 32'h8 ? _T_91[31:0] : _GEN_472; // @[ivncontrol4.scala 191:42 194:21]
  wire [31:0] _GEN_480 = _GEN_336 >= 32'h8 ? _T_91[31:0] : _GEN_473; // @[ivncontrol4.scala 191:42 195:21]
  wire [31:0] _GEN_481 = _GEN_336 >= 32'h8 ? _T_91[31:0] : _GEN_474; // @[ivncontrol4.scala 191:42 196:22]
  wire [31:0] _GEN_482 = _GEN_336 >= 32'h8 ? _T_91[31:0] : _GEN_475; // @[ivncontrol4.scala 191:42 197:22]
  wire [31:0] _GEN_483 = _GEN_336 >= 32'h8 ? _T_91[31:0] : _GEN_476; // @[ivncontrol4.scala 191:42 198:22]
  wire [31:0] _GEN_484 = _GEN_336 >= 32'h8 ? _T_91[31:0] : 32'h6; // @[ivncontrol4.scala 143:18 191:42 199:22]
  wire [31:0] _T_127 = 32'h8 - _GEN_336; // @[ivncontrol4.scala 245:18]
  wire [31:0] _i_vn_1_T_15 = 32'h1 + pin; // @[ivncontrol4.scala 246:29]
  wire [31:0] _GEN_597 = _T_127 == 32'h1 ? _i_vn_1_T_15 : _GEN_484; // @[ivncontrol4.scala 286:54 289:22]
  wire [31:0] _GEN_598 = _T_127 == 32'h2 ? _i_vn_1_T_15 : _GEN_483; // @[ivncontrol4.scala 281:54 284:22]
  wire [31:0] _GEN_599 = _T_127 == 32'h2 ? _i_vn_1_T_15 : _GEN_597; // @[ivncontrol4.scala 281:54 285:22]
  wire [31:0] _GEN_600 = _T_127 == 32'h3 ? _i_vn_1_T_15 : _GEN_482; // @[ivncontrol4.scala 274:54 276:22]
  wire [31:0] _GEN_601 = _T_127 == 32'h3 ? _i_vn_1_T_15 : _GEN_598; // @[ivncontrol4.scala 274:54 277:22]
  wire [31:0] _GEN_602 = _T_127 == 32'h3 ? _i_vn_1_T_15 : _GEN_599; // @[ivncontrol4.scala 274:54 278:22]
  wire [31:0] _GEN_603 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_481; // @[ivncontrol4.scala 268:54 270:22]
  wire [31:0] _GEN_604 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_600; // @[ivncontrol4.scala 268:54 271:22]
  wire [31:0] _GEN_605 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_601; // @[ivncontrol4.scala 268:54 272:22]
  wire [31:0] _GEN_606 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_602; // @[ivncontrol4.scala 268:54 273:22]
  wire [31:0] _GEN_607 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_480; // @[ivncontrol4.scala 261:54 263:21]
  wire [31:0] _GEN_608 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_603; // @[ivncontrol4.scala 261:54 264:22]
  wire [31:0] _GEN_609 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_604; // @[ivncontrol4.scala 261:54 265:22]
  wire [31:0] _GEN_610 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_605; // @[ivncontrol4.scala 261:54 266:22]
  wire [31:0] _GEN_611 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_606; // @[ivncontrol4.scala 261:54 267:22]
  wire [31:0] _GEN_612 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_479; // @[ivncontrol4.scala 254:54 255:22]
  wire [31:0] _GEN_613 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_607; // @[ivncontrol4.scala 254:54 256:21]
  wire [31:0] _GEN_614 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_608; // @[ivncontrol4.scala 254:54 257:22]
  wire [31:0] _GEN_615 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_609; // @[ivncontrol4.scala 254:54 258:22]
  wire [31:0] _GEN_616 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_610; // @[ivncontrol4.scala 254:54 259:22]
  wire [31:0] _GEN_617 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_611; // @[ivncontrol4.scala 254:54 260:22]
  wire [31:0] _GEN_618 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_478; // @[ivncontrol4.scala 245:49 246:22]
  wire [31:0] _GEN_619 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_612; // @[ivncontrol4.scala 245:49 247:21]
  wire [31:0] _GEN_620 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_613; // @[ivncontrol4.scala 245:49 248:21]
  wire [31:0] _GEN_621 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_614; // @[ivncontrol4.scala 245:49 249:22]
  wire [31:0] _GEN_622 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_615; // @[ivncontrol4.scala 245:49 250:22]
  wire [31:0] _GEN_623 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_616; // @[ivncontrol4.scala 245:49 251:22]
  wire [31:0] _GEN_624 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_617; // @[ivncontrol4.scala 245:49 252:22]
  wire [31:0] _GEN_642 = 4'h1 == _i_vn_1_T_15[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_643 = 4'h2 == _i_vn_1_T_15[3:0] ? rowcount_2 : _GEN_642; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_644 = 4'h3 == _i_vn_1_T_15[3:0] ? rowcount_3 : _GEN_643; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_645 = 4'h4 == _i_vn_1_T_15[3:0] ? rowcount_4 : _GEN_644; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_646 = 4'h5 == _i_vn_1_T_15[3:0] ? rowcount_5 : _GEN_645; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_647 = 4'h6 == _i_vn_1_T_15[3:0] ? rowcount_6 : _GEN_646; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_648 = 4'h7 == _i_vn_1_T_15[3:0] ? rowcount_7 : _GEN_647; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_649 = 4'h8 == _i_vn_1_T_15[3:0] ? rowcount_8 : _GEN_648; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_650 = 4'h9 == _i_vn_1_T_15[3:0] ? rowcount_9 : _GEN_649; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_651 = 4'ha == _i_vn_1_T_15[3:0] ? rowcount_10 : _GEN_650; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_652 = 4'hb == _i_vn_1_T_15[3:0] ? rowcount_11 : _GEN_651; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_653 = 4'hc == _i_vn_1_T_15[3:0] ? rowcount_12 : _GEN_652; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_654 = 4'hd == _i_vn_1_T_15[3:0] ? rowcount_13 : _GEN_653; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_655 = 4'he == _i_vn_1_T_15[3:0] ? rowcount_14 : _GEN_654; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_656 = 4'hf == _i_vn_1_T_15[3:0] ? rowcount_15 : _GEN_655; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _T_172 = _GEN_336 + _GEN_656; // @[ivncontrol4.scala 292:41]
  wire [31:0] _T_174 = 32'h8 - _T_172; // @[ivncontrol4.scala 292:18]
  wire [31:0] _i_vn_1_T_17 = 32'h2 + pin; // @[ivncontrol4.scala 293:29]
  wire [31:0] _GEN_849 = _T_174 == 32'h1 ? _i_vn_1_T_17 : _GEN_624; // @[ivncontrol4.scala 335:78 338:22]
  wire [31:0] _GEN_850 = _T_174 == 32'h2 ? _i_vn_1_T_17 : _GEN_623; // @[ivncontrol4.scala 329:76 332:22]
  wire [31:0] _GEN_851 = _T_174 == 32'h2 ? _i_vn_1_T_17 : _GEN_849; // @[ivncontrol4.scala 329:76 333:22]
  wire [31:0] _GEN_852 = _T_174 == 32'h3 ? _i_vn_1_T_17 : _GEN_622; // @[ivncontrol4.scala 322:78 324:23]
  wire [31:0] _GEN_853 = _T_174 == 32'h3 ? _i_vn_1_T_17 : _GEN_850; // @[ivncontrol4.scala 322:78 325:22]
  wire [31:0] _GEN_854 = _T_174 == 32'h3 ? _i_vn_1_T_17 : _GEN_851; // @[ivncontrol4.scala 322:78 326:22]
  wire [31:0] _GEN_855 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_621; // @[ivncontrol4.scala 316:78 318:22]
  wire [31:0] _GEN_856 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_852; // @[ivncontrol4.scala 316:78 319:22]
  wire [31:0] _GEN_857 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_853; // @[ivncontrol4.scala 316:78 320:22]
  wire [31:0] _GEN_858 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_854; // @[ivncontrol4.scala 316:78 321:22]
  wire [31:0] _GEN_859 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_620; // @[ivncontrol4.scala 309:76 311:23]
  wire [31:0] _GEN_860 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_855; // @[ivncontrol4.scala 309:76 312:22]
  wire [31:0] _GEN_861 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_856; // @[ivncontrol4.scala 309:76 313:22]
  wire [31:0] _GEN_862 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_857; // @[ivncontrol4.scala 309:76 314:22]
  wire [31:0] _GEN_863 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_858; // @[ivncontrol4.scala 309:76 315:22]
  wire [31:0] _GEN_864 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_619; // @[ivncontrol4.scala 301:77 303:22]
  wire [31:0] _GEN_865 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_859; // @[ivncontrol4.scala 301:77 304:21]
  wire [31:0] _GEN_866 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_860; // @[ivncontrol4.scala 301:77 305:22]
  wire [31:0] _GEN_867 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_861; // @[ivncontrol4.scala 301:77 306:22]
  wire [31:0] _GEN_868 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_862; // @[ivncontrol4.scala 301:77 307:22]
  wire [31:0] _GEN_869 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_863; // @[ivncontrol4.scala 301:77 308:22]
  wire [31:0] _GEN_870 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_618; // @[ivncontrol4.scala 292:73 293:22]
  wire [31:0] _GEN_871 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_864; // @[ivncontrol4.scala 292:73 294:21]
  wire [31:0] _GEN_872 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_865; // @[ivncontrol4.scala 292:73 295:21]
  wire [31:0] _GEN_873 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_866; // @[ivncontrol4.scala 292:73 296:22]
  wire [31:0] _GEN_874 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_867; // @[ivncontrol4.scala 292:73 297:22]
  wire [31:0] _GEN_875 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_868; // @[ivncontrol4.scala 292:73 298:22]
  wire [31:0] _GEN_876 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_869; // @[ivncontrol4.scala 292:73 299:22]
  wire [31:0] _GEN_910 = 4'h1 == _i_vn_1_T_17[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_911 = 4'h2 == _i_vn_1_T_17[3:0] ? rowcount_2 : _GEN_910; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_912 = 4'h3 == _i_vn_1_T_17[3:0] ? rowcount_3 : _GEN_911; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_913 = 4'h4 == _i_vn_1_T_17[3:0] ? rowcount_4 : _GEN_912; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_914 = 4'h5 == _i_vn_1_T_17[3:0] ? rowcount_5 : _GEN_913; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_915 = 4'h6 == _i_vn_1_T_17[3:0] ? rowcount_6 : _GEN_914; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_916 = 4'h7 == _i_vn_1_T_17[3:0] ? rowcount_7 : _GEN_915; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_917 = 4'h8 == _i_vn_1_T_17[3:0] ? rowcount_8 : _GEN_916; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_918 = 4'h9 == _i_vn_1_T_17[3:0] ? rowcount_9 : _GEN_917; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_919 = 4'ha == _i_vn_1_T_17[3:0] ? rowcount_10 : _GEN_918; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_920 = 4'hb == _i_vn_1_T_17[3:0] ? rowcount_11 : _GEN_919; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_921 = 4'hc == _i_vn_1_T_17[3:0] ? rowcount_12 : _GEN_920; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_922 = 4'hd == _i_vn_1_T_17[3:0] ? rowcount_13 : _GEN_921; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_923 = 4'he == _i_vn_1_T_17[3:0] ? rowcount_14 : _GEN_922; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_924 = 4'hf == _i_vn_1_T_17[3:0] ? rowcount_15 : _GEN_923; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _T_254 = _T_172 + _GEN_924; // @[ivncontrol4.scala 343:62]
  wire [31:0] _T_256 = 32'h8 - _T_254; // @[ivncontrol4.scala 343:17]
  wire [31:0] _i_vn_1_T_19 = 32'h3 + pin; // @[ivncontrol4.scala 344:29]
  wire [31:0] _GEN_1213 = _T_256 == 32'h1 ? _i_vn_1_T_19 : _GEN_876; // @[ivncontrol4.scala 386:100 389:22]
  wire [31:0] _GEN_1214 = _T_256 == 32'h2 ? _i_vn_1_T_19 : _GEN_875; // @[ivncontrol4.scala 380:98 383:22]
  wire [31:0] _GEN_1215 = _T_256 == 32'h2 ? _i_vn_1_T_19 : _GEN_1213; // @[ivncontrol4.scala 380:98 384:22]
  wire [31:0] _GEN_1216 = _T_256 == 32'h3 ? _i_vn_1_T_19 : _GEN_874; // @[ivncontrol4.scala 373:100 375:23]
  wire [31:0] _GEN_1217 = _T_256 == 32'h3 ? _i_vn_1_T_19 : _GEN_1214; // @[ivncontrol4.scala 373:100 376:22]
  wire [31:0] _GEN_1218 = _T_256 == 32'h3 ? _i_vn_1_T_19 : _GEN_1215; // @[ivncontrol4.scala 373:100 377:22]
  wire [31:0] _GEN_1219 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_873; // @[ivncontrol4.scala 367:100 369:22]
  wire [31:0] _GEN_1220 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_1216; // @[ivncontrol4.scala 367:100 370:22]
  wire [31:0] _GEN_1221 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_1217; // @[ivncontrol4.scala 367:100 371:22]
  wire [31:0] _GEN_1222 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_1218; // @[ivncontrol4.scala 367:100 372:22]
  wire [31:0] _GEN_1223 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_872; // @[ivncontrol4.scala 360:98 362:23]
  wire [31:0] _GEN_1224 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1219; // @[ivncontrol4.scala 360:98 363:22]
  wire [31:0] _GEN_1225 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1220; // @[ivncontrol4.scala 360:98 364:22]
  wire [31:0] _GEN_1226 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1221; // @[ivncontrol4.scala 360:98 365:22]
  wire [31:0] _GEN_1227 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1222; // @[ivncontrol4.scala 360:98 366:22]
  wire [31:0] _GEN_1228 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_871; // @[ivncontrol4.scala 352:99 354:22]
  wire [31:0] _GEN_1229 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1223; // @[ivncontrol4.scala 352:99 355:21]
  wire [31:0] _GEN_1230 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1224; // @[ivncontrol4.scala 352:99 356:22]
  wire [31:0] _GEN_1231 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1225; // @[ivncontrol4.scala 352:99 357:22]
  wire [31:0] _GEN_1232 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1226; // @[ivncontrol4.scala 352:99 358:22]
  wire [31:0] _GEN_1233 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1227; // @[ivncontrol4.scala 352:99 359:22]
  wire [31:0] _GEN_1234 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_870; // @[ivncontrol4.scala 343:94 344:22]
  wire [31:0] _GEN_1235 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1228; // @[ivncontrol4.scala 343:94 345:21]
  wire [31:0] _GEN_1236 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1229; // @[ivncontrol4.scala 343:94 346:21]
  wire [31:0] _GEN_1237 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1230; // @[ivncontrol4.scala 343:94 347:22]
  wire [31:0] _GEN_1238 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1231; // @[ivncontrol4.scala 343:94 348:22]
  wire [31:0] _GEN_1239 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1232; // @[ivncontrol4.scala 343:94 349:22]
  wire [31:0] _GEN_1240 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1233; // @[ivncontrol4.scala 343:94 350:22]
  wire [31:0] _GEN_1290 = 4'h1 == _i_vn_1_T_19[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1291 = 4'h2 == _i_vn_1_T_19[3:0] ? rowcount_2 : _GEN_1290; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1292 = 4'h3 == _i_vn_1_T_19[3:0] ? rowcount_3 : _GEN_1291; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1293 = 4'h4 == _i_vn_1_T_19[3:0] ? rowcount_4 : _GEN_1292; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1294 = 4'h5 == _i_vn_1_T_19[3:0] ? rowcount_5 : _GEN_1293; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1295 = 4'h6 == _i_vn_1_T_19[3:0] ? rowcount_6 : _GEN_1294; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1296 = 4'h7 == _i_vn_1_T_19[3:0] ? rowcount_7 : _GEN_1295; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1297 = 4'h8 == _i_vn_1_T_19[3:0] ? rowcount_8 : _GEN_1296; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1298 = 4'h9 == _i_vn_1_T_19[3:0] ? rowcount_9 : _GEN_1297; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1299 = 4'ha == _i_vn_1_T_19[3:0] ? rowcount_10 : _GEN_1298; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1300 = 4'hb == _i_vn_1_T_19[3:0] ? rowcount_11 : _GEN_1299; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1301 = 4'hc == _i_vn_1_T_19[3:0] ? rowcount_12 : _GEN_1300; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1302 = 4'hd == _i_vn_1_T_19[3:0] ? rowcount_13 : _GEN_1301; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1303 = 4'he == _i_vn_1_T_19[3:0] ? rowcount_14 : _GEN_1302; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1304 = 4'hf == _i_vn_1_T_19[3:0] ? rowcount_15 : _GEN_1303; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _T_371 = _T_254 + _GEN_1304; // @[ivncontrol4.scala 393:86]
  wire [31:0] _T_373 = 32'h8 - _T_371; // @[ivncontrol4.scala 393:19]
  wire [31:0] _i_vn_1_T_21 = 32'h4 + pin; // @[ivncontrol4.scala 394:29]
  wire [31:0] _GEN_1689 = _T_373 == 32'h1 ? _i_vn_1_T_21 : _GEN_1240; // @[ivncontrol4.scala 436:122 439:22]
  wire [31:0] _GEN_1690 = _T_373 == 32'h2 ? _i_vn_1_T_21 : _GEN_1239; // @[ivncontrol4.scala 430:121 433:22]
  wire [31:0] _GEN_1691 = _T_373 == 32'h2 ? _i_vn_1_T_21 : _GEN_1689; // @[ivncontrol4.scala 430:121 434:22]
  wire [31:0] _GEN_1692 = _T_373 == 32'h3 ? _i_vn_1_T_21 : _GEN_1238; // @[ivncontrol4.scala 423:123 425:23]
  wire [31:0] _GEN_1693 = _T_373 == 32'h3 ? _i_vn_1_T_21 : _GEN_1690; // @[ivncontrol4.scala 423:123 426:22]
  wire [31:0] _GEN_1694 = _T_373 == 32'h3 ? _i_vn_1_T_21 : _GEN_1691; // @[ivncontrol4.scala 423:123 427:22]
  wire [31:0] _GEN_1695 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1237; // @[ivncontrol4.scala 417:122 419:22]
  wire [31:0] _GEN_1696 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1692; // @[ivncontrol4.scala 417:122 420:22]
  wire [31:0] _GEN_1697 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1693; // @[ivncontrol4.scala 417:122 421:22]
  wire [31:0] _GEN_1698 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1694; // @[ivncontrol4.scala 417:122 422:22]
  wire [31:0] _GEN_1699 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1236; // @[ivncontrol4.scala 410:121 412:23]
  wire [31:0] _GEN_1700 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1695; // @[ivncontrol4.scala 410:121 413:22]
  wire [31:0] _GEN_1701 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1696; // @[ivncontrol4.scala 410:121 414:22]
  wire [31:0] _GEN_1702 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1697; // @[ivncontrol4.scala 410:121 415:22]
  wire [31:0] _GEN_1703 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1698; // @[ivncontrol4.scala 410:121 416:22]
  wire [31:0] _GEN_1704 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1235; // @[ivncontrol4.scala 402:121 404:22]
  wire [31:0] _GEN_1705 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1699; // @[ivncontrol4.scala 402:121 405:21]
  wire [31:0] _GEN_1706 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1700; // @[ivncontrol4.scala 402:121 406:22]
  wire [31:0] _GEN_1707 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1701; // @[ivncontrol4.scala 402:121 407:22]
  wire [31:0] _GEN_1708 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1702; // @[ivncontrol4.scala 402:121 408:22]
  wire [31:0] _GEN_1709 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1703; // @[ivncontrol4.scala 402:121 409:22]
  wire [31:0] _GEN_1710 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1234; // @[ivncontrol4.scala 393:118 394:22]
  wire [31:0] _GEN_1711 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1704; // @[ivncontrol4.scala 393:118 395:21]
  wire [31:0] _GEN_1712 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1705; // @[ivncontrol4.scala 393:118 396:21]
  wire [31:0] _GEN_1713 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1706; // @[ivncontrol4.scala 393:118 397:22]
  wire [31:0] _GEN_1714 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1707; // @[ivncontrol4.scala 393:118 398:22]
  wire [31:0] _GEN_1715 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1708; // @[ivncontrol4.scala 393:118 399:22]
  wire [31:0] _GEN_1716 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1709; // @[ivncontrol4.scala 393:118 400:22]
  wire [31:0] _GEN_1782 = 4'h1 == _i_vn_1_T_21[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1783 = 4'h2 == _i_vn_1_T_21[3:0] ? rowcount_2 : _GEN_1782; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1784 = 4'h3 == _i_vn_1_T_21[3:0] ? rowcount_3 : _GEN_1783; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1785 = 4'h4 == _i_vn_1_T_21[3:0] ? rowcount_4 : _GEN_1784; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1786 = 4'h5 == _i_vn_1_T_21[3:0] ? rowcount_5 : _GEN_1785; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1787 = 4'h6 == _i_vn_1_T_21[3:0] ? rowcount_6 : _GEN_1786; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1788 = 4'h7 == _i_vn_1_T_21[3:0] ? rowcount_7 : _GEN_1787; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1789 = 4'h8 == _i_vn_1_T_21[3:0] ? rowcount_8 : _GEN_1788; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1790 = 4'h9 == _i_vn_1_T_21[3:0] ? rowcount_9 : _GEN_1789; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1791 = 4'ha == _i_vn_1_T_21[3:0] ? rowcount_10 : _GEN_1790; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1792 = 4'hb == _i_vn_1_T_21[3:0] ? rowcount_11 : _GEN_1791; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1793 = 4'hc == _i_vn_1_T_21[3:0] ? rowcount_12 : _GEN_1792; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1794 = 4'hd == _i_vn_1_T_21[3:0] ? rowcount_13 : _GEN_1793; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1795 = 4'he == _i_vn_1_T_21[3:0] ? rowcount_14 : _GEN_1794; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1796 = 4'hf == _i_vn_1_T_21[3:0] ? rowcount_15 : _GEN_1795; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _T_523 = _T_371 + _GEN_1796; // @[ivncontrol4.scala 443:108]
  wire [31:0] _T_525 = 32'h8 - _T_523; // @[ivncontrol4.scala 443:19]
  wire [31:0] _i_vn_1_T_23 = 32'h5 + pin; // @[ivncontrol4.scala 444:29]
  wire [31:0] _GEN_2277 = _T_525 == 32'h1 ? _i_vn_1_T_23 : _GEN_1716; // @[ivncontrol4.scala 486:144 489:22]
  wire [31:0] _GEN_2278 = _T_525 == 32'h2 ? _i_vn_1_T_23 : _GEN_1715; // @[ivncontrol4.scala 480:143 483:22]
  wire [31:0] _GEN_2279 = _T_525 == 32'h2 ? _i_vn_1_T_23 : _GEN_2277; // @[ivncontrol4.scala 480:143 484:22]
  wire [31:0] _GEN_2280 = _T_525 == 32'h3 ? _i_vn_1_T_23 : _GEN_1714; // @[ivncontrol4.scala 473:145 475:23]
  wire [31:0] _GEN_2281 = _T_525 == 32'h3 ? _i_vn_1_T_23 : _GEN_2278; // @[ivncontrol4.scala 473:145 476:22]
  wire [31:0] _GEN_2282 = _T_525 == 32'h3 ? _i_vn_1_T_23 : _GEN_2279; // @[ivncontrol4.scala 473:145 477:22]
  wire [31:0] _GEN_2283 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_1713; // @[ivncontrol4.scala 467:143 469:22]
  wire [31:0] _GEN_2284 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_2280; // @[ivncontrol4.scala 467:143 470:22]
  wire [31:0] _GEN_2285 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_2281; // @[ivncontrol4.scala 467:143 471:22]
  wire [31:0] _GEN_2286 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_2282; // @[ivncontrol4.scala 467:143 472:22]
  wire [31:0] _GEN_2287 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_1712; // @[ivncontrol4.scala 460:143 462:23]
  wire [31:0] _GEN_2288 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2283; // @[ivncontrol4.scala 460:143 463:22]
  wire [31:0] _GEN_2289 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2284; // @[ivncontrol4.scala 460:143 464:22]
  wire [31:0] _GEN_2290 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2285; // @[ivncontrol4.scala 460:143 465:22]
  wire [31:0] _GEN_2291 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2286; // @[ivncontrol4.scala 460:143 466:22]
  wire [31:0] _GEN_2292 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_1711; // @[ivncontrol4.scala 452:143 454:22]
  wire [31:0] _GEN_2293 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2287; // @[ivncontrol4.scala 452:143 455:21]
  wire [31:0] _GEN_2294 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2288; // @[ivncontrol4.scala 452:143 456:22]
  wire [31:0] _GEN_2295 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2289; // @[ivncontrol4.scala 452:143 457:22]
  wire [31:0] _GEN_2296 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2290; // @[ivncontrol4.scala 452:143 458:22]
  wire [31:0] _GEN_2297 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2291; // @[ivncontrol4.scala 452:143 459:22]
  wire [31:0] _GEN_2298 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_1710; // @[ivncontrol4.scala 443:140 444:22]
  wire [31:0] _GEN_2299 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2292; // @[ivncontrol4.scala 443:140 445:21]
  wire [31:0] _GEN_2300 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2293; // @[ivncontrol4.scala 443:140 446:21]
  wire [31:0] _GEN_2301 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2294; // @[ivncontrol4.scala 443:140 447:22]
  wire [31:0] _GEN_2302 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2295; // @[ivncontrol4.scala 443:140 448:22]
  wire [31:0] _GEN_2303 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2296; // @[ivncontrol4.scala 443:140 449:22]
  wire [31:0] _GEN_2304 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2297; // @[ivncontrol4.scala 443:140 450:22]
  wire [31:0] _GEN_2386 = 4'h1 == _i_vn_1_T_23[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2387 = 4'h2 == _i_vn_1_T_23[3:0] ? rowcount_2 : _GEN_2386; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2388 = 4'h3 == _i_vn_1_T_23[3:0] ? rowcount_3 : _GEN_2387; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2389 = 4'h4 == _i_vn_1_T_23[3:0] ? rowcount_4 : _GEN_2388; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2390 = 4'h5 == _i_vn_1_T_23[3:0] ? rowcount_5 : _GEN_2389; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2391 = 4'h6 == _i_vn_1_T_23[3:0] ? rowcount_6 : _GEN_2390; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2392 = 4'h7 == _i_vn_1_T_23[3:0] ? rowcount_7 : _GEN_2391; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2393 = 4'h8 == _i_vn_1_T_23[3:0] ? rowcount_8 : _GEN_2392; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2394 = 4'h9 == _i_vn_1_T_23[3:0] ? rowcount_9 : _GEN_2393; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2395 = 4'ha == _i_vn_1_T_23[3:0] ? rowcount_10 : _GEN_2394; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2396 = 4'hb == _i_vn_1_T_23[3:0] ? rowcount_11 : _GEN_2395; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2397 = 4'hc == _i_vn_1_T_23[3:0] ? rowcount_12 : _GEN_2396; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2398 = 4'hd == _i_vn_1_T_23[3:0] ? rowcount_13 : _GEN_2397; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2399 = 4'he == _i_vn_1_T_23[3:0] ? rowcount_14 : _GEN_2398; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2400 = 4'hf == _i_vn_1_T_23[3:0] ? rowcount_15 : _GEN_2399; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _T_710 = _T_523 + _GEN_2400; // @[ivncontrol4.scala 494:130]
  wire [31:0] _T_712 = 32'h8 - _T_710; // @[ivncontrol4.scala 494:19]
  wire [31:0] _i_vn_1_T_25 = 32'h6 + pin; // @[ivncontrol4.scala 495:29]
  wire [31:0] _GEN_2977 = _T_712 == 32'h1 ? _i_vn_1_T_25 : _GEN_2304; // @[ivncontrol4.scala 537:166 540:22]
  wire [31:0] _GEN_2978 = _T_712 == 32'h2 ? _i_vn_1_T_25 : _GEN_2303; // @[ivncontrol4.scala 531:166 534:22]
  wire [31:0] _GEN_2979 = _T_712 == 32'h2 ? _i_vn_1_T_25 : _GEN_2977; // @[ivncontrol4.scala 531:166 535:22]
  wire [31:0] _GEN_2980 = _T_712 == 32'h3 ? _i_vn_1_T_25 : _GEN_2302; // @[ivncontrol4.scala 524:168 526:23]
  wire [31:0] _GEN_2981 = _T_712 == 32'h3 ? _i_vn_1_T_25 : _GEN_2978; // @[ivncontrol4.scala 524:168 527:22]
  wire [31:0] _GEN_2982 = _T_712 == 32'h3 ? _i_vn_1_T_25 : _GEN_2979; // @[ivncontrol4.scala 524:168 528:22]
  wire [31:0] _GEN_2983 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2301; // @[ivncontrol4.scala 518:166 520:22]
  wire [31:0] _GEN_2984 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2980; // @[ivncontrol4.scala 518:166 521:22]
  wire [31:0] _GEN_2985 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2981; // @[ivncontrol4.scala 518:166 522:22]
  wire [31:0] _GEN_2986 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2982; // @[ivncontrol4.scala 518:166 523:22]
  wire [31:0] _GEN_2987 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2300; // @[ivncontrol4.scala 511:166 513:23]
  wire [31:0] _GEN_2988 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2983; // @[ivncontrol4.scala 511:166 514:22]
  wire [31:0] _GEN_2989 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2984; // @[ivncontrol4.scala 511:166 515:22]
  wire [31:0] _GEN_2990 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2985; // @[ivncontrol4.scala 511:166 516:22]
  wire [31:0] _GEN_2991 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2986; // @[ivncontrol4.scala 511:166 517:22]
  wire [31:0] _GEN_2992 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2299; // @[ivncontrol4.scala 503:166 505:22]
  wire [31:0] _GEN_2993 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2987; // @[ivncontrol4.scala 503:166 506:21]
  wire [31:0] _GEN_2994 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2988; // @[ivncontrol4.scala 503:166 507:22]
  wire [31:0] _GEN_2995 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2989; // @[ivncontrol4.scala 503:166 508:22]
  wire [31:0] _GEN_2996 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2990; // @[ivncontrol4.scala 503:166 509:22]
  wire [31:0] _GEN_2997 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2991; // @[ivncontrol4.scala 503:166 510:22]
  wire [31:0] _GEN_2998 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2298; // @[ivncontrol4.scala 494:162 495:22]
  wire [31:0] _GEN_2999 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2992; // @[ivncontrol4.scala 494:162 496:21]
  wire [31:0] _GEN_3000 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2993; // @[ivncontrol4.scala 494:162 497:21]
  wire [31:0] _GEN_3001 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2994; // @[ivncontrol4.scala 494:162 498:22]
  wire [31:0] _GEN_3002 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2995; // @[ivncontrol4.scala 494:162 499:22]
  wire [31:0] _GEN_3003 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2996; // @[ivncontrol4.scala 494:162 500:22]
  wire [31:0] _GEN_3004 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2997; // @[ivncontrol4.scala 494:162 501:22]
  wire [31:0] _GEN_3102 = 4'h1 == _i_vn_1_T_25[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3103 = 4'h2 == _i_vn_1_T_25[3:0] ? rowcount_2 : _GEN_3102; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3104 = 4'h3 == _i_vn_1_T_25[3:0] ? rowcount_3 : _GEN_3103; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3105 = 4'h4 == _i_vn_1_T_25[3:0] ? rowcount_4 : _GEN_3104; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3106 = 4'h5 == _i_vn_1_T_25[3:0] ? rowcount_5 : _GEN_3105; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3107 = 4'h6 == _i_vn_1_T_25[3:0] ? rowcount_6 : _GEN_3106; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3108 = 4'h7 == _i_vn_1_T_25[3:0] ? rowcount_7 : _GEN_3107; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3109 = 4'h8 == _i_vn_1_T_25[3:0] ? rowcount_8 : _GEN_3108; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3110 = 4'h9 == _i_vn_1_T_25[3:0] ? rowcount_9 : _GEN_3109; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3111 = 4'ha == _i_vn_1_T_25[3:0] ? rowcount_10 : _GEN_3110; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3112 = 4'hb == _i_vn_1_T_25[3:0] ? rowcount_11 : _GEN_3111; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3113 = 4'hc == _i_vn_1_T_25[3:0] ? rowcount_12 : _GEN_3112; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3114 = 4'hd == _i_vn_1_T_25[3:0] ? rowcount_13 : _GEN_3113; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3115 = 4'he == _i_vn_1_T_25[3:0] ? rowcount_14 : _GEN_3114; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3116 = 4'hf == _i_vn_1_T_25[3:0] ? rowcount_15 : _GEN_3115; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _T_932 = _T_710 + _GEN_3116; // @[ivncontrol4.scala 545:152]
  wire [31:0] _T_934 = 32'h8 - _T_932; // @[ivncontrol4.scala 545:19]
  wire [31:0] _i_vn_1_T_27 = 32'h7 + pin; // @[ivncontrol4.scala 546:29]
  wire [31:0] _GEN_3789 = _T_934 == 32'h1 ? _i_vn_1_T_27 : _GEN_3004; // @[ivncontrol4.scala 588:188 591:22]
  wire [31:0] _GEN_3790 = _T_934 == 32'h2 ? _i_vn_1_T_27 : _GEN_3003; // @[ivncontrol4.scala 582:188 585:22]
  wire [31:0] _GEN_3791 = _T_934 == 32'h2 ? _i_vn_1_T_27 : _GEN_3789; // @[ivncontrol4.scala 582:188 586:22]
  wire [31:0] _GEN_3792 = _T_934 == 32'h3 ? _i_vn_1_T_27 : _GEN_3002; // @[ivncontrol4.scala 575:190 577:23]
  wire [31:0] _GEN_3793 = _T_934 == 32'h3 ? _i_vn_1_T_27 : _GEN_3790; // @[ivncontrol4.scala 575:190 578:22]
  wire [31:0] _GEN_3794 = _T_934 == 32'h3 ? _i_vn_1_T_27 : _GEN_3791; // @[ivncontrol4.scala 575:190 579:22]
  wire [31:0] _GEN_3795 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_3001; // @[ivncontrol4.scala 569:188 571:22]
  wire [31:0] _GEN_3796 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_3792; // @[ivncontrol4.scala 569:188 572:22]
  wire [31:0] _GEN_3797 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_3793; // @[ivncontrol4.scala 569:188 573:22]
  wire [31:0] _GEN_3798 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_3794; // @[ivncontrol4.scala 569:188 574:22]
  wire [31:0] _GEN_3799 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3000; // @[ivncontrol4.scala 562:188 564:23]
  wire [31:0] _GEN_3800 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3795; // @[ivncontrol4.scala 562:188 565:22]
  wire [31:0] _GEN_3801 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3796; // @[ivncontrol4.scala 562:188 566:22]
  wire [31:0] _GEN_3802 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3797; // @[ivncontrol4.scala 562:188 567:22]
  wire [31:0] _GEN_3803 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3798; // @[ivncontrol4.scala 562:188 568:22]
  wire [31:0] _GEN_3804 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_2999; // @[ivncontrol4.scala 554:188 556:22]
  wire [31:0] _GEN_3805 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3799; // @[ivncontrol4.scala 554:188 557:21]
  wire [31:0] _GEN_3806 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3800; // @[ivncontrol4.scala 554:188 558:22]
  wire [31:0] _GEN_3807 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3801; // @[ivncontrol4.scala 554:188 559:22]
  wire [31:0] _GEN_3808 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3802; // @[ivncontrol4.scala 554:188 560:22]
  wire [31:0] _GEN_3809 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3803; // @[ivncontrol4.scala 554:188 561:22]
  wire [31:0] _GEN_3810 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_2998; // @[ivncontrol4.scala 545:184 546:22]
  wire [31:0] _GEN_3811 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3804; // @[ivncontrol4.scala 545:184 547:21]
  wire [31:0] _GEN_3812 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3805; // @[ivncontrol4.scala 545:184 548:21]
  wire [31:0] _GEN_3813 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3806; // @[ivncontrol4.scala 545:184 549:22]
  wire [31:0] _GEN_3814 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3807; // @[ivncontrol4.scala 545:184 550:22]
  wire [31:0] _GEN_3815 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3808; // @[ivncontrol4.scala 545:184 551:22]
  wire [31:0] _GEN_3816 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3809; // @[ivncontrol4.scala 545:184 552:22]
  wire [31:0] _GEN_3817 = _GEN_312 ? _GEN_477 : 32'h3; // @[ivncontrol4.scala 142:17 189:28]
  wire [31:0] _GEN_3818 = _GEN_312 ? _GEN_3810 : 32'h1; // @[ivncontrol4.scala 142:17 189:28]
  wire [31:0] _GEN_3819 = _GEN_312 ? _GEN_3811 : 32'h19; // @[ivncontrol4.scala 142:17 189:28]
  wire [31:0] _GEN_3820 = _GEN_312 ? _GEN_3812 : 32'hf; // @[ivncontrol4.scala 142:17 189:28]
  wire [31:0] _GEN_3821 = _GEN_312 ? _GEN_3813 : 32'h10; // @[ivncontrol4.scala 143:18 189:28]
  wire [31:0] _GEN_3822 = _GEN_312 ? _GEN_3814 : 32'h4; // @[ivncontrol4.scala 143:18 189:28]
  wire [31:0] _GEN_3823 = _GEN_312 ? _GEN_3815 : 32'h12; // @[ivncontrol4.scala 143:18 189:28]
  wire [31:0] _GEN_3824 = _GEN_312 ? _GEN_3816 : 32'h6; // @[ivncontrol4.scala 143:18 189:28]
  wire  valid1 = 1'h0;
  wire [31:0] _GEN_4221 = reset ? 32'h0 : _GEN_3817; // @[ivncontrol4.scala 17:{23,23}]
  wire [31:0] _GEN_4222 = reset ? 32'h0 : _GEN_3818; // @[ivncontrol4.scala 17:{23,23}]
  wire [31:0] _GEN_4223 = reset ? 32'h0 : _GEN_3819; // @[ivncontrol4.scala 17:{23,23}]
  wire [31:0] _GEN_4224 = reset ? 32'h0 : _GEN_3820; // @[ivncontrol4.scala 17:{23,23}]
  wire [31:0] _GEN_4225 = reset ? 32'h0 : _GEN_3821; // @[ivncontrol4.scala 18:{24,24}]
  wire [31:0] _GEN_4226 = reset ? 32'h0 : _GEN_3822; // @[ivncontrol4.scala 18:{24,24}]
  wire [31:0] _GEN_4227 = reset ? 32'h0 : _GEN_3823; // @[ivncontrol4.scala 18:{24,24}]
  wire [31:0] _GEN_4228 = reset ? 32'h0 : _GEN_3824; // @[ivncontrol4.scala 18:{24,24}]
  assign io_o_vn_0 = i_vn_0; // @[ivncontrol4.scala 138:13]
  assign io_o_vn_1 = i_vn_1; // @[ivncontrol4.scala 138:13]
  assign io_o_vn_2 = i_vn_2; // @[ivncontrol4.scala 138:13]
  assign io_o_vn_3 = i_vn_3; // @[ivncontrol4.scala 138:13]
  assign io_o_vn2_0 = i_vn2_0; // @[ivncontrol4.scala 139:14]
  assign io_o_vn2_1 = i_vn2_1; // @[ivncontrol4.scala 139:14]
  assign io_o_vn2_2 = i_vn2_2; // @[ivncontrol4.scala 139:14]
  assign io_o_vn2_3 = i_vn2_3; // @[ivncontrol4.scala 139:14]
  always @(posedge clock) begin
    i_vn_0 <= _GEN_4221[4:0]; // @[ivncontrol4.scala 17:{23,23}]
    i_vn_1 <= _GEN_4222[4:0]; // @[ivncontrol4.scala 17:{23,23}]
    i_vn_2 <= _GEN_4223[4:0]; // @[ivncontrol4.scala 17:{23,23}]
    i_vn_3 <= _GEN_4224[4:0]; // @[ivncontrol4.scala 17:{23,23}]
    i_vn2_0 <= _GEN_4225[4:0]; // @[ivncontrol4.scala 18:{24,24}]
    i_vn2_1 <= _GEN_4226[4:0]; // @[ivncontrol4.scala 18:{24,24}]
    i_vn2_2 <= _GEN_4227[4:0]; // @[ivncontrol4.scala 18:{24,24}]
    i_vn2_3 <= _GEN_4228[4:0]; // @[ivncontrol4.scala 18:{24,24}]
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_0 <= io_Stationary_matrix_0_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_1 <= io_Stationary_matrix_0_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_2 <= io_Stationary_matrix_0_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_3 <= io_Stationary_matrix_0_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_4 <= io_Stationary_matrix_0_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_5 <= io_Stationary_matrix_0_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_6 <= io_Stationary_matrix_0_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_7 <= io_Stationary_matrix_0_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_0 <= io_Stationary_matrix_1_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_1 <= io_Stationary_matrix_1_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_2 <= io_Stationary_matrix_1_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_3 <= io_Stationary_matrix_1_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_4 <= io_Stationary_matrix_1_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_5 <= io_Stationary_matrix_1_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_6 <= io_Stationary_matrix_1_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_7 <= io_Stationary_matrix_1_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_0 <= io_Stationary_matrix_2_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_1 <= io_Stationary_matrix_2_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_2 <= io_Stationary_matrix_2_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_3 <= io_Stationary_matrix_2_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_4 <= io_Stationary_matrix_2_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_5 <= io_Stationary_matrix_2_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_6 <= io_Stationary_matrix_2_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_7 <= io_Stationary_matrix_2_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_0 <= io_Stationary_matrix_3_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_1 <= io_Stationary_matrix_3_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_2 <= io_Stationary_matrix_3_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_3 <= io_Stationary_matrix_3_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_4 <= io_Stationary_matrix_3_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_5 <= io_Stationary_matrix_3_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_6 <= io_Stationary_matrix_3_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_7 <= io_Stationary_matrix_3_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_0 <= io_Stationary_matrix_4_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_1 <= io_Stationary_matrix_4_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_2 <= io_Stationary_matrix_4_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_3 <= io_Stationary_matrix_4_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_4 <= io_Stationary_matrix_4_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_5 <= io_Stationary_matrix_4_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_6 <= io_Stationary_matrix_4_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_7 <= io_Stationary_matrix_4_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_0 <= io_Stationary_matrix_5_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_1 <= io_Stationary_matrix_5_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_2 <= io_Stationary_matrix_5_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_3 <= io_Stationary_matrix_5_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_4 <= io_Stationary_matrix_5_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_5 <= io_Stationary_matrix_5_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_6 <= io_Stationary_matrix_5_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_7 <= io_Stationary_matrix_5_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_0 <= io_Stationary_matrix_6_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_1 <= io_Stationary_matrix_6_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_2 <= io_Stationary_matrix_6_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_3 <= io_Stationary_matrix_6_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_4 <= io_Stationary_matrix_6_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_5 <= io_Stationary_matrix_6_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_6 <= io_Stationary_matrix_6_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_7 <= io_Stationary_matrix_6_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_0 <= io_Stationary_matrix_7_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_1 <= io_Stationary_matrix_7_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_2 <= io_Stationary_matrix_7_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_3 <= io_Stationary_matrix_7_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_4 <= io_Stationary_matrix_7_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_5 <= io_Stationary_matrix_7_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_6 <= io_Stationary_matrix_7_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_7 <= io_Stationary_matrix_7_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_0 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_0 <= count_0; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_1 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_1 <= count_1; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_2 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_2 <= count_2; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_3 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_3 <= count_3; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_4 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_4 <= count_4; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_5 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_5 <= count_5; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_6 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_6 <= count_6; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_7 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_7 <= count_7; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_8 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_8 <= 32'h0; // @[ivncontrol4.scala 87:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_9 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_9 <= 32'h0; // @[ivncontrol4.scala 87:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_10 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_10 <= 32'h0; // @[ivncontrol4.scala 87:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_11 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_11 <= 32'h0; // @[ivncontrol4.scala 87:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_12 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_12 <= 32'h0; // @[ivncontrol4.scala 87:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_13 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_13 <= 32'h0; // @[ivncontrol4.scala 87:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_14 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_14 <= 32'h0; // @[ivncontrol4.scala 87:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_15 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end
    if (reset) begin // @[ivncontrol4.scala 37:22]
      pin <= 32'h0; // @[ivncontrol4.scala 37:22]
    end else if (_T_72 & rowcount_6 == 32'h0 & rowcount_7 != 32'h0) begin // @[ivncontrol4.scala 183:192]
      pin <= 32'h7; // @[ivncontrol4.scala 184:13]
    end else if (_T_59 & rowcount_5 == 32'h0 & rowcount_6 != 32'h0) begin // @[ivncontrol4.scala 180:169]
      pin <= 32'h6; // @[ivncontrol4.scala 181:13]
    end else if (_T_48 & rowcount_4 == 32'h0 & rowcount_5 != 32'h0) begin // @[ivncontrol4.scala 177:146]
      pin <= 32'h5; // @[ivncontrol4.scala 178:13]
    end else begin
      pin <= _GEN_317;
    end
    if (reset) begin // @[ivncontrol4.scala 41:20]
      i <= 32'h0; // @[ivncontrol4.scala 41:20]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
        i <= _GEN_247;
      end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
        i <= _GEN_247;
      end else begin
        i <= _GEN_265;
      end
    end
    if (reset) begin // @[ivncontrol4.scala 42:20]
      j <= 32'h0; // @[ivncontrol4.scala 42:20]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
        j <= 32'h8; // @[ivncontrol4.scala 116:11]
      end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
        j <= _j_T_1; // @[ivncontrol4.scala 118:11]
      end else begin
        j <= {{28'd0}, _GEN_264};
      end
    end
    if (3'h0 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h0 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h0 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h0 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h0 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h0 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h0 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h0 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_0 <= _GEN_224;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_0 <= _GEN_224;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h0 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_0 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_0 <= _GEN_224;
      end
    end else begin
      count_0 <= _GEN_224;
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_1 <= _GEN_225;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_1 <= _GEN_225;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h1 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_1 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_1 <= _GEN_225;
      end
    end else begin
      count_1 <= _GEN_225;
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_2 <= _GEN_226;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_2 <= _GEN_226;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h2 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_2 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_2 <= _GEN_226;
      end
    end else begin
      count_2 <= _GEN_226;
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_3 <= _GEN_227;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_3 <= _GEN_227;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h3 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_3 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_3 <= _GEN_227;
      end
    end else begin
      count_3 <= _GEN_227;
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_4 <= _GEN_228;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_4 <= _GEN_228;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h4 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_4 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_4 <= _GEN_228;
      end
    end else begin
      count_4 <= _GEN_228;
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_5 <= _GEN_229;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_5 <= _GEN_229;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h5 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_5 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_5 <= _GEN_229;
      end
    end else begin
      count_5 <= _GEN_229;
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_6 <= _GEN_230;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_6 <= _GEN_230;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h6 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_6 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_6 <= _GEN_230;
      end
    end else begin
      count_6 <= _GEN_230;
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_7 <= _GEN_231;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_7 <= _GEN_231;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h7 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_7 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_7 <= _GEN_231;
      end
    end else begin
      count_7 <= _GEN_231;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  i_vn_0 = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  i_vn_1 = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  i_vn_2 = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  i_vn_3 = _RAND_3[4:0];
  _RAND_4 = {1{`RANDOM}};
  i_vn2_0 = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  i_vn2_1 = _RAND_5[4:0];
  _RAND_6 = {1{`RANDOM}};
  i_vn2_2 = _RAND_6[4:0];
  _RAND_7 = {1{`RANDOM}};
  i_vn2_3 = _RAND_7[4:0];
  _RAND_8 = {1{`RANDOM}};
  solution_0_0 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  solution_0_1 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  solution_0_2 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  solution_0_3 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  solution_0_4 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  solution_0_5 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  solution_0_6 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  solution_0_7 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  solution_1_0 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  solution_1_1 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  solution_1_2 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  solution_1_3 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  solution_1_4 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  solution_1_5 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  solution_1_6 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  solution_1_7 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  solution_2_0 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  solution_2_1 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  solution_2_2 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  solution_2_3 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  solution_2_4 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  solution_2_5 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  solution_2_6 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  solution_2_7 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  solution_3_0 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  solution_3_1 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  solution_3_2 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  solution_3_3 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  solution_3_4 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  solution_3_5 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  solution_3_6 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  solution_3_7 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  solution_4_0 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  solution_4_1 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  solution_4_2 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  solution_4_3 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  solution_4_4 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  solution_4_5 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  solution_4_6 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  solution_4_7 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  solution_5_0 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  solution_5_1 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  solution_5_2 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  solution_5_3 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  solution_5_4 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  solution_5_5 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  solution_5_6 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  solution_5_7 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  solution_6_0 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  solution_6_1 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  solution_6_2 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  solution_6_3 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  solution_6_4 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  solution_6_5 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  solution_6_6 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  solution_6_7 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  solution_7_0 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  solution_7_1 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  solution_7_2 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  solution_7_3 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  solution_7_4 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  solution_7_5 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  solution_7_6 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  solution_7_7 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  rowcount_0 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  rowcount_1 = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  rowcount_2 = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  rowcount_3 = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  rowcount_4 = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  rowcount_5 = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  rowcount_6 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  rowcount_7 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  rowcount_8 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  rowcount_9 = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  rowcount_10 = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  rowcount_11 = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  rowcount_12 = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  rowcount_13 = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  rowcount_14 = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  rowcount_15 = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  pin = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  i = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  j = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  mat_0_0 = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  mat_0_1 = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  mat_0_2 = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  mat_0_3 = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  mat_0_4 = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  mat_0_5 = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  mat_0_6 = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  mat_0_7 = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  mat_1_0 = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  mat_1_1 = _RAND_100[31:0];
  _RAND_101 = {1{`RANDOM}};
  mat_1_2 = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  mat_1_3 = _RAND_102[31:0];
  _RAND_103 = {1{`RANDOM}};
  mat_1_4 = _RAND_103[31:0];
  _RAND_104 = {1{`RANDOM}};
  mat_1_5 = _RAND_104[31:0];
  _RAND_105 = {1{`RANDOM}};
  mat_1_6 = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  mat_1_7 = _RAND_106[31:0];
  _RAND_107 = {1{`RANDOM}};
  mat_2_0 = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  mat_2_1 = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  mat_2_2 = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  mat_2_3 = _RAND_110[31:0];
  _RAND_111 = {1{`RANDOM}};
  mat_2_4 = _RAND_111[31:0];
  _RAND_112 = {1{`RANDOM}};
  mat_2_5 = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  mat_2_6 = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  mat_2_7 = _RAND_114[31:0];
  _RAND_115 = {1{`RANDOM}};
  mat_3_0 = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  mat_3_1 = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  mat_3_2 = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  mat_3_3 = _RAND_118[31:0];
  _RAND_119 = {1{`RANDOM}};
  mat_3_4 = _RAND_119[31:0];
  _RAND_120 = {1{`RANDOM}};
  mat_3_5 = _RAND_120[31:0];
  _RAND_121 = {1{`RANDOM}};
  mat_3_6 = _RAND_121[31:0];
  _RAND_122 = {1{`RANDOM}};
  mat_3_7 = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  mat_4_0 = _RAND_123[31:0];
  _RAND_124 = {1{`RANDOM}};
  mat_4_1 = _RAND_124[31:0];
  _RAND_125 = {1{`RANDOM}};
  mat_4_2 = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  mat_4_3 = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  mat_4_4 = _RAND_127[31:0];
  _RAND_128 = {1{`RANDOM}};
  mat_4_5 = _RAND_128[31:0];
  _RAND_129 = {1{`RANDOM}};
  mat_4_6 = _RAND_129[31:0];
  _RAND_130 = {1{`RANDOM}};
  mat_4_7 = _RAND_130[31:0];
  _RAND_131 = {1{`RANDOM}};
  mat_5_0 = _RAND_131[31:0];
  _RAND_132 = {1{`RANDOM}};
  mat_5_1 = _RAND_132[31:0];
  _RAND_133 = {1{`RANDOM}};
  mat_5_2 = _RAND_133[31:0];
  _RAND_134 = {1{`RANDOM}};
  mat_5_3 = _RAND_134[31:0];
  _RAND_135 = {1{`RANDOM}};
  mat_5_4 = _RAND_135[31:0];
  _RAND_136 = {1{`RANDOM}};
  mat_5_5 = _RAND_136[31:0];
  _RAND_137 = {1{`RANDOM}};
  mat_5_6 = _RAND_137[31:0];
  _RAND_138 = {1{`RANDOM}};
  mat_5_7 = _RAND_138[31:0];
  _RAND_139 = {1{`RANDOM}};
  mat_6_0 = _RAND_139[31:0];
  _RAND_140 = {1{`RANDOM}};
  mat_6_1 = _RAND_140[31:0];
  _RAND_141 = {1{`RANDOM}};
  mat_6_2 = _RAND_141[31:0];
  _RAND_142 = {1{`RANDOM}};
  mat_6_3 = _RAND_142[31:0];
  _RAND_143 = {1{`RANDOM}};
  mat_6_4 = _RAND_143[31:0];
  _RAND_144 = {1{`RANDOM}};
  mat_6_5 = _RAND_144[31:0];
  _RAND_145 = {1{`RANDOM}};
  mat_6_6 = _RAND_145[31:0];
  _RAND_146 = {1{`RANDOM}};
  mat_6_7 = _RAND_146[31:0];
  _RAND_147 = {1{`RANDOM}};
  mat_7_0 = _RAND_147[31:0];
  _RAND_148 = {1{`RANDOM}};
  mat_7_1 = _RAND_148[31:0];
  _RAND_149 = {1{`RANDOM}};
  mat_7_2 = _RAND_149[31:0];
  _RAND_150 = {1{`RANDOM}};
  mat_7_3 = _RAND_150[31:0];
  _RAND_151 = {1{`RANDOM}};
  mat_7_4 = _RAND_151[31:0];
  _RAND_152 = {1{`RANDOM}};
  mat_7_5 = _RAND_152[31:0];
  _RAND_153 = {1{`RANDOM}};
  mat_7_6 = _RAND_153[31:0];
  _RAND_154 = {1{`RANDOM}};
  mat_7_7 = _RAND_154[31:0];
  _RAND_155 = {1{`RANDOM}};
  count_0 = _RAND_155[31:0];
  _RAND_156 = {1{`RANDOM}};
  count_1 = _RAND_156[31:0];
  _RAND_157 = {1{`RANDOM}};
  count_2 = _RAND_157[31:0];
  _RAND_158 = {1{`RANDOM}};
  count_3 = _RAND_158[31:0];
  _RAND_159 = {1{`RANDOM}};
  count_4 = _RAND_159[31:0];
  _RAND_160 = {1{`RANDOM}};
  count_5 = _RAND_160[31:0];
  _RAND_161 = {1{`RANDOM}};
  count_6 = _RAND_161[31:0];
  _RAND_162 = {1{`RANDOM}};
  count_7 = _RAND_162[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ivncontrol4_5(
  input         clock,
  input         reset,
  input  [15:0] io_Stationary_matrix_0_0,
  input  [15:0] io_Stationary_matrix_0_1,
  input  [15:0] io_Stationary_matrix_0_2,
  input  [15:0] io_Stationary_matrix_0_3,
  input  [15:0] io_Stationary_matrix_0_4,
  input  [15:0] io_Stationary_matrix_0_5,
  input  [15:0] io_Stationary_matrix_0_6,
  input  [15:0] io_Stationary_matrix_0_7,
  input  [15:0] io_Stationary_matrix_1_0,
  input  [15:0] io_Stationary_matrix_1_1,
  input  [15:0] io_Stationary_matrix_1_2,
  input  [15:0] io_Stationary_matrix_1_3,
  input  [15:0] io_Stationary_matrix_1_4,
  input  [15:0] io_Stationary_matrix_1_5,
  input  [15:0] io_Stationary_matrix_1_6,
  input  [15:0] io_Stationary_matrix_1_7,
  input  [15:0] io_Stationary_matrix_2_0,
  input  [15:0] io_Stationary_matrix_2_1,
  input  [15:0] io_Stationary_matrix_2_2,
  input  [15:0] io_Stationary_matrix_2_3,
  input  [15:0] io_Stationary_matrix_2_4,
  input  [15:0] io_Stationary_matrix_2_5,
  input  [15:0] io_Stationary_matrix_2_6,
  input  [15:0] io_Stationary_matrix_2_7,
  input  [15:0] io_Stationary_matrix_3_0,
  input  [15:0] io_Stationary_matrix_3_1,
  input  [15:0] io_Stationary_matrix_3_2,
  input  [15:0] io_Stationary_matrix_3_3,
  input  [15:0] io_Stationary_matrix_3_4,
  input  [15:0] io_Stationary_matrix_3_5,
  input  [15:0] io_Stationary_matrix_3_6,
  input  [15:0] io_Stationary_matrix_3_7,
  input  [15:0] io_Stationary_matrix_4_0,
  input  [15:0] io_Stationary_matrix_4_1,
  input  [15:0] io_Stationary_matrix_4_2,
  input  [15:0] io_Stationary_matrix_4_3,
  input  [15:0] io_Stationary_matrix_4_4,
  input  [15:0] io_Stationary_matrix_4_5,
  input  [15:0] io_Stationary_matrix_4_6,
  input  [15:0] io_Stationary_matrix_4_7,
  input  [15:0] io_Stationary_matrix_5_0,
  input  [15:0] io_Stationary_matrix_5_1,
  input  [15:0] io_Stationary_matrix_5_2,
  input  [15:0] io_Stationary_matrix_5_3,
  input  [15:0] io_Stationary_matrix_5_4,
  input  [15:0] io_Stationary_matrix_5_5,
  input  [15:0] io_Stationary_matrix_5_6,
  input  [15:0] io_Stationary_matrix_5_7,
  input  [15:0] io_Stationary_matrix_6_0,
  input  [15:0] io_Stationary_matrix_6_1,
  input  [15:0] io_Stationary_matrix_6_2,
  input  [15:0] io_Stationary_matrix_6_3,
  input  [15:0] io_Stationary_matrix_6_4,
  input  [15:0] io_Stationary_matrix_6_5,
  input  [15:0] io_Stationary_matrix_6_6,
  input  [15:0] io_Stationary_matrix_6_7,
  input  [15:0] io_Stationary_matrix_7_0,
  input  [15:0] io_Stationary_matrix_7_1,
  input  [15:0] io_Stationary_matrix_7_2,
  input  [15:0] io_Stationary_matrix_7_3,
  input  [15:0] io_Stationary_matrix_7_4,
  input  [15:0] io_Stationary_matrix_7_5,
  input  [15:0] io_Stationary_matrix_7_6,
  input  [15:0] io_Stationary_matrix_7_7,
  output [4:0]  io_o_vn_0,
  output [4:0]  io_o_vn_1,
  output [4:0]  io_o_vn_2,
  output [4:0]  io_o_vn_3,
  output [4:0]  io_o_vn2_0,
  output [4:0]  io_o_vn2_1,
  output [4:0]  io_o_vn2_2,
  output [4:0]  io_o_vn2_3,
  input         io_validpin
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
`endif // RANDOMIZE_REG_INIT
  reg [4:0] i_vn_0; // @[ivncontrol4.scala 17:23]
  reg [4:0] i_vn_1; // @[ivncontrol4.scala 17:23]
  reg [4:0] i_vn_2; // @[ivncontrol4.scala 17:23]
  reg [4:0] i_vn_3; // @[ivncontrol4.scala 17:23]
  reg [4:0] i_vn2_0; // @[ivncontrol4.scala 18:24]
  reg [4:0] i_vn2_1; // @[ivncontrol4.scala 18:24]
  reg [4:0] i_vn2_2; // @[ivncontrol4.scala 18:24]
  reg [4:0] i_vn2_3; // @[ivncontrol4.scala 18:24]
  reg [15:0] solution_0_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_0_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_0_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_0_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_0_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_0_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_0_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_0_7; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_7; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_7; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_7; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_7; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_7; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_7; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_7; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_0; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_1; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_2; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_3; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_4; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_5; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_6; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_7; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_8; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_9; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_10; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_11; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_12; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_13; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_14; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_15; // @[ivncontrol4.scala 27:27]
  reg [31:0] pin; // @[ivncontrol4.scala 37:22]
  reg [31:0] i; // @[ivncontrol4.scala 41:20]
  reg [31:0] j; // @[ivncontrol4.scala 42:20]
  wire  _io_ProcessValid_T = i == 32'h7; // @[ivncontrol4.scala 44:27]
  wire  _io_ProcessValid_T_1 = j == 32'h7; // @[ivncontrol4.scala 44:42]
  wire  _io_ProcessValid_T_2 = i == 32'h7 & j == 32'h7; // @[ivncontrol4.scala 44:36]
  reg [31:0] mat_0_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_0_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_0_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_0_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_0_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_0_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_0_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_0_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] count_0; // @[ivncontrol4.scala 58:20]
  reg [31:0] count_1; // @[ivncontrol4.scala 58:20]
  reg [31:0] count_2; // @[ivncontrol4.scala 58:20]
  reg [31:0] count_3; // @[ivncontrol4.scala 58:20]
  reg [31:0] count_4; // @[ivncontrol4.scala 58:20]
  reg [31:0] count_5; // @[ivncontrol4.scala 58:20]
  reg [31:0] count_6; // @[ivncontrol4.scala 58:20]
  reg [31:0] count_7; // @[ivncontrol4.scala 58:20]
  wire  _GEN_3825 = 3'h0 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_65 = 3'h0 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_0_1 : io_Stationary_matrix_0_0; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_66 = 3'h0 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_0_2 : _GEN_65; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_67 = 3'h0 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_0_3 : _GEN_66; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_68 = 3'h0 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_0_4 : _GEN_67; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_69 = 3'h0 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_0_5 : _GEN_68; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_70 = 3'h0 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_0_6 : _GEN_69; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_71 = 3'h0 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_0_7 : _GEN_70; // @[ivncontrol4.scala 63:{17,17}]
  wire  _GEN_3839 = 3'h1 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_72 = 3'h1 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_1_0 : _GEN_71; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_73 = 3'h1 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_1_1 : _GEN_72; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_74 = 3'h1 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_1_2 : _GEN_73; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_75 = 3'h1 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_1_3 : _GEN_74; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_76 = 3'h1 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_1_4 : _GEN_75; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_77 = 3'h1 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_1_5 : _GEN_76; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_78 = 3'h1 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_1_6 : _GEN_77; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_79 = 3'h1 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_1_7 : _GEN_78; // @[ivncontrol4.scala 63:{17,17}]
  wire  _GEN_3855 = 3'h2 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_80 = 3'h2 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_2_0 : _GEN_79; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_81 = 3'h2 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_2_1 : _GEN_80; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_82 = 3'h2 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_2_2 : _GEN_81; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_83 = 3'h2 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_2_3 : _GEN_82; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_84 = 3'h2 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_2_4 : _GEN_83; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_85 = 3'h2 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_2_5 : _GEN_84; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_86 = 3'h2 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_2_6 : _GEN_85; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_87 = 3'h2 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_2_7 : _GEN_86; // @[ivncontrol4.scala 63:{17,17}]
  wire  _GEN_3871 = 3'h3 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_88 = 3'h3 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_3_0 : _GEN_87; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_89 = 3'h3 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_3_1 : _GEN_88; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_90 = 3'h3 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_3_2 : _GEN_89; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_91 = 3'h3 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_3_3 : _GEN_90; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_92 = 3'h3 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_3_4 : _GEN_91; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_93 = 3'h3 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_3_5 : _GEN_92; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_94 = 3'h3 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_3_6 : _GEN_93; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_95 = 3'h3 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_3_7 : _GEN_94; // @[ivncontrol4.scala 63:{17,17}]
  wire  _GEN_3887 = 3'h4 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_96 = 3'h4 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_4_0 : _GEN_95; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_97 = 3'h4 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_4_1 : _GEN_96; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_98 = 3'h4 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_4_2 : _GEN_97; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_99 = 3'h4 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_4_3 : _GEN_98; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_100 = 3'h4 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_4_4 : _GEN_99; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_101 = 3'h4 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_4_5 : _GEN_100; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_102 = 3'h4 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_4_6 : _GEN_101; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_103 = 3'h4 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_4_7 : _GEN_102; // @[ivncontrol4.scala 63:{17,17}]
  wire  _GEN_3903 = 3'h5 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_104 = 3'h5 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_5_0 : _GEN_103; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_105 = 3'h5 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_5_1 : _GEN_104; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_106 = 3'h5 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_5_2 : _GEN_105; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_107 = 3'h5 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_5_3 : _GEN_106; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_108 = 3'h5 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_5_4 : _GEN_107; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_109 = 3'h5 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_5_5 : _GEN_108; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_110 = 3'h5 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_5_6 : _GEN_109; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_111 = 3'h5 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_5_7 : _GEN_110; // @[ivncontrol4.scala 63:{17,17}]
  wire  _GEN_3919 = 3'h6 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_112 = 3'h6 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_6_0 : _GEN_111; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_113 = 3'h6 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_6_1 : _GEN_112; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_114 = 3'h6 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_6_2 : _GEN_113; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_115 = 3'h6 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_6_3 : _GEN_114; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_116 = 3'h6 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_6_4 : _GEN_115; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_117 = 3'h6 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_6_5 : _GEN_116; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_118 = 3'h6 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_6_6 : _GEN_117; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_119 = 3'h6 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_6_7 : _GEN_118; // @[ivncontrol4.scala 63:{17,17}]
  wire  _GEN_3935 = 3'h7 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_120 = 3'h7 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_7_0 : _GEN_119; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_121 = 3'h7 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_7_1 : _GEN_120; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_122 = 3'h7 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_7_2 : _GEN_121; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_123 = 3'h7 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_7_3 : _GEN_122; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_124 = 3'h7 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_7_4 : _GEN_123; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_125 = 3'h7 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_7_5 : _GEN_124; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_126 = 3'h7 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_7_6 : _GEN_125; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_127 = 3'h7 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_7_7 : _GEN_126; // @[ivncontrol4.scala 63:{17,17}]
  wire [31:0] _mat_T_1_T_2 = {{16'd0}, _GEN_127}; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_129 = _GEN_3825 & 4'h1 == j[3:0] ? solution_0_1 : solution_0_0; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_130 = _GEN_3825 & 4'h2 == j[3:0] ? solution_0_2 : _GEN_129; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_131 = _GEN_3825 & 4'h3 == j[3:0] ? solution_0_3 : _GEN_130; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_132 = _GEN_3825 & 4'h4 == j[3:0] ? solution_0_4 : _GEN_131; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_133 = _GEN_3825 & 4'h5 == j[3:0] ? solution_0_5 : _GEN_132; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_134 = _GEN_3825 & 4'h6 == j[3:0] ? solution_0_6 : _GEN_133; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_135 = _GEN_3825 & 4'h7 == j[3:0] ? solution_0_7 : _GEN_134; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_136 = _GEN_3825 & 4'h8 == j[3:0] ? 16'h0 : _GEN_135; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_137 = _GEN_3839 & 4'h0 == j[3:0] ? solution_1_0 : _GEN_136; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_138 = _GEN_3839 & 4'h1 == j[3:0] ? solution_1_1 : _GEN_137; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_139 = _GEN_3839 & 4'h2 == j[3:0] ? solution_1_2 : _GEN_138; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_140 = _GEN_3839 & 4'h3 == j[3:0] ? solution_1_3 : _GEN_139; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_141 = _GEN_3839 & 4'h4 == j[3:0] ? solution_1_4 : _GEN_140; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_142 = _GEN_3839 & 4'h5 == j[3:0] ? solution_1_5 : _GEN_141; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_143 = _GEN_3839 & 4'h6 == j[3:0] ? solution_1_6 : _GEN_142; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_144 = _GEN_3839 & 4'h7 == j[3:0] ? solution_1_7 : _GEN_143; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_145 = _GEN_3839 & 4'h8 == j[3:0] ? 16'h0 : _GEN_144; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_146 = _GEN_3855 & 4'h0 == j[3:0] ? solution_2_0 : _GEN_145; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_147 = _GEN_3855 & 4'h1 == j[3:0] ? solution_2_1 : _GEN_146; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_148 = _GEN_3855 & 4'h2 == j[3:0] ? solution_2_2 : _GEN_147; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_149 = _GEN_3855 & 4'h3 == j[3:0] ? solution_2_3 : _GEN_148; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_150 = _GEN_3855 & 4'h4 == j[3:0] ? solution_2_4 : _GEN_149; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_151 = _GEN_3855 & 4'h5 == j[3:0] ? solution_2_5 : _GEN_150; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_152 = _GEN_3855 & 4'h6 == j[3:0] ? solution_2_6 : _GEN_151; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_153 = _GEN_3855 & 4'h7 == j[3:0] ? solution_2_7 : _GEN_152; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_154 = _GEN_3855 & 4'h8 == j[3:0] ? 16'h0 : _GEN_153; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_155 = _GEN_3871 & 4'h0 == j[3:0] ? solution_3_0 : _GEN_154; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_156 = _GEN_3871 & 4'h1 == j[3:0] ? solution_3_1 : _GEN_155; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_157 = _GEN_3871 & 4'h2 == j[3:0] ? solution_3_2 : _GEN_156; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_158 = _GEN_3871 & 4'h3 == j[3:0] ? solution_3_3 : _GEN_157; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_159 = _GEN_3871 & 4'h4 == j[3:0] ? solution_3_4 : _GEN_158; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_160 = _GEN_3871 & 4'h5 == j[3:0] ? solution_3_5 : _GEN_159; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_161 = _GEN_3871 & 4'h6 == j[3:0] ? solution_3_6 : _GEN_160; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_162 = _GEN_3871 & 4'h7 == j[3:0] ? solution_3_7 : _GEN_161; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_163 = _GEN_3871 & 4'h8 == j[3:0] ? 16'h0 : _GEN_162; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_164 = _GEN_3887 & 4'h0 == j[3:0] ? solution_4_0 : _GEN_163; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_165 = _GEN_3887 & 4'h1 == j[3:0] ? solution_4_1 : _GEN_164; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_166 = _GEN_3887 & 4'h2 == j[3:0] ? solution_4_2 : _GEN_165; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_167 = _GEN_3887 & 4'h3 == j[3:0] ? solution_4_3 : _GEN_166; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_168 = _GEN_3887 & 4'h4 == j[3:0] ? solution_4_4 : _GEN_167; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_169 = _GEN_3887 & 4'h5 == j[3:0] ? solution_4_5 : _GEN_168; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_170 = _GEN_3887 & 4'h6 == j[3:0] ? solution_4_6 : _GEN_169; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_171 = _GEN_3887 & 4'h7 == j[3:0] ? solution_4_7 : _GEN_170; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_172 = _GEN_3887 & 4'h8 == j[3:0] ? 16'h0 : _GEN_171; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_173 = _GEN_3903 & 4'h0 == j[3:0] ? solution_5_0 : _GEN_172; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_174 = _GEN_3903 & 4'h1 == j[3:0] ? solution_5_1 : _GEN_173; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_175 = _GEN_3903 & 4'h2 == j[3:0] ? solution_5_2 : _GEN_174; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_176 = _GEN_3903 & 4'h3 == j[3:0] ? solution_5_3 : _GEN_175; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_177 = _GEN_3903 & 4'h4 == j[3:0] ? solution_5_4 : _GEN_176; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_178 = _GEN_3903 & 4'h5 == j[3:0] ? solution_5_5 : _GEN_177; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_179 = _GEN_3903 & 4'h6 == j[3:0] ? solution_5_6 : _GEN_178; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_180 = _GEN_3903 & 4'h7 == j[3:0] ? solution_5_7 : _GEN_179; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_181 = _GEN_3903 & 4'h8 == j[3:0] ? 16'h0 : _GEN_180; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_182 = _GEN_3919 & 4'h0 == j[3:0] ? solution_6_0 : _GEN_181; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_183 = _GEN_3919 & 4'h1 == j[3:0] ? solution_6_1 : _GEN_182; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_184 = _GEN_3919 & 4'h2 == j[3:0] ? solution_6_2 : _GEN_183; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_185 = _GEN_3919 & 4'h3 == j[3:0] ? solution_6_3 : _GEN_184; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_186 = _GEN_3919 & 4'h4 == j[3:0] ? solution_6_4 : _GEN_185; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_187 = _GEN_3919 & 4'h5 == j[3:0] ? solution_6_5 : _GEN_186; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_188 = _GEN_3919 & 4'h6 == j[3:0] ? solution_6_6 : _GEN_187; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_189 = _GEN_3919 & 4'h7 == j[3:0] ? solution_6_7 : _GEN_188; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_190 = _GEN_3919 & 4'h8 == j[3:0] ? 16'h0 : _GEN_189; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_191 = _GEN_3935 & 4'h0 == j[3:0] ? solution_7_0 : _GEN_190; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_192 = _GEN_3935 & 4'h1 == j[3:0] ? solution_7_1 : _GEN_191; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_193 = _GEN_3935 & 4'h2 == j[3:0] ? solution_7_2 : _GEN_192; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_194 = _GEN_3935 & 4'h3 == j[3:0] ? solution_7_3 : _GEN_193; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_195 = _GEN_3935 & 4'h4 == j[3:0] ? solution_7_4 : _GEN_194; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_196 = _GEN_3935 & 4'h5 == j[3:0] ? solution_7_5 : _GEN_195; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_197 = _GEN_3935 & 4'h6 == j[3:0] ? solution_7_6 : _GEN_196; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_198 = _GEN_3935 & 4'h7 == j[3:0] ? solution_7_7 : _GEN_197; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_199 = _GEN_3935 & 4'h8 == j[3:0] ? 16'h0 : _GEN_198; // @[ivncontrol4.scala 65:{31,31}]
  wire [31:0] _GEN_201 = 3'h1 == i[2:0] ? count_1 : count_0; // @[ivncontrol4.scala 66:{33,33}]
  wire [31:0] _GEN_202 = 3'h2 == i[2:0] ? count_2 : _GEN_201; // @[ivncontrol4.scala 66:{33,33}]
  wire [31:0] _GEN_203 = 3'h3 == i[2:0] ? count_3 : _GEN_202; // @[ivncontrol4.scala 66:{33,33}]
  wire [31:0] _GEN_204 = 3'h4 == i[2:0] ? count_4 : _GEN_203; // @[ivncontrol4.scala 66:{33,33}]
  wire [31:0] _GEN_205 = 3'h5 == i[2:0] ? count_5 : _GEN_204; // @[ivncontrol4.scala 66:{33,33}]
  wire [31:0] _GEN_206 = 3'h6 == i[2:0] ? count_6 : _GEN_205; // @[ivncontrol4.scala 66:{33,33}]
  wire [31:0] _GEN_207 = 3'h7 == i[2:0] ? count_7 : _GEN_206; // @[ivncontrol4.scala 66:{33,33}]
  wire [31:0] _count_T_2 = _GEN_207 + 32'h1; // @[ivncontrol4.scala 66:33]
  wire [31:0] _GEN_208 = 3'h0 == i[2:0] ? _count_T_2 : count_0; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_209 = 3'h1 == i[2:0] ? _count_T_2 : count_1; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_210 = 3'h2 == i[2:0] ? _count_T_2 : count_2; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_211 = 3'h3 == i[2:0] ? _count_T_2 : count_3; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_212 = 3'h4 == i[2:0] ? _count_T_2 : count_4; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_213 = 3'h5 == i[2:0] ? _count_T_2 : count_5; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_214 = 3'h6 == i[2:0] ? _count_T_2 : count_6; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_215 = 3'h7 == i[2:0] ? _count_T_2 : count_7; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_216 = _GEN_199 != 16'h0 ? _GEN_208 : count_0; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_217 = _GEN_199 != 16'h0 ? _GEN_209 : count_1; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_218 = _GEN_199 != 16'h0 ? _GEN_210 : count_2; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_219 = _GEN_199 != 16'h0 ? _GEN_211 : count_3; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_220 = _GEN_199 != 16'h0 ? _GEN_212 : count_4; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_221 = _GEN_199 != 16'h0 ? _GEN_213 : count_5; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_222 = _GEN_199 != 16'h0 ? _GEN_214 : count_6; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_223 = _GEN_199 != 16'h0 ? _GEN_215 : count_7; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_224 = io_validpin ? _GEN_216 : count_0; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _GEN_225 = io_validpin ? _GEN_217 : count_1; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _GEN_226 = io_validpin ? _GEN_218 : count_2; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _GEN_227 = io_validpin ? _GEN_219 : count_3; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _GEN_228 = io_validpin ? _GEN_220 : count_4; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _GEN_229 = io_validpin ? _GEN_221 : count_5; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _GEN_230 = io_validpin ? _GEN_222 : count_6; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _GEN_231 = io_validpin ? _GEN_223 : count_7; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _i_T_1 = i + 32'h1; // @[ivncontrol4.scala 113:16]
  wire [31:0] _GEN_247 = i < 32'h7 & _io_ProcessValid_T_1 ? _i_T_1 : i; // @[ivncontrol4.scala 112:74 113:11 41:20]
  wire [31:0] _j_T_1 = j + 32'h1; // @[ivncontrol4.scala 118:16]
  wire [3:0] _GEN_264 = _io_ProcessValid_T & j == 32'h8 ? 4'h8 : 4'h0; // @[ivncontrol4.scala 120:77 121:11 129:11]
  wire [31:0] _GEN_265 = _io_ProcessValid_T & j == 32'h8 ? 32'h7 : _GEN_247; // @[ivncontrol4.scala 120:77 122:11]
  wire  _GEN_312 = _io_ProcessValid_T_2; // @[ivncontrol4.scala 153:41]
  wire [31:0] _GEN_313 = rowcount_0 != 32'h0 ? 32'h0 : pin; // @[ivncontrol4.scala 162:30 163:13 37:22]
  wire  _T_27 = rowcount_0 == 32'h0; // @[ivncontrol4.scala 165:23]
  wire [31:0] _GEN_314 = rowcount_0 == 32'h0 & rowcount_1 != 32'h0 ? 32'h1 : _GEN_313; // @[ivncontrol4.scala 165:54 166:13]
  wire  _T_32 = _T_27 & rowcount_1 == 32'h0; // @[ivncontrol4.scala 168:31]
  wire [31:0] _GEN_315 = _T_27 & rowcount_1 == 32'h0 & rowcount_2 != 32'h0 ? 32'h2 : _GEN_314; // @[ivncontrol4.scala 168:77 169:13]
  wire  _T_39 = _T_32 & rowcount_2 == 32'h0; // @[ivncontrol4.scala 171:54]
  wire [31:0] _GEN_316 = _T_32 & rowcount_2 == 32'h0 & rowcount_3 != 32'h0 ? 32'h3 : _GEN_315; // @[ivncontrol4.scala 171:100 172:13]
  wire  _T_48 = _T_39 & rowcount_3 == 32'h0; // @[ivncontrol4.scala 174:77]
  wire [31:0] _GEN_317 = _T_39 & rowcount_3 == 32'h0 & rowcount_4 != 32'h0 ? 32'h4 : _GEN_316; // @[ivncontrol4.scala 174:123 175:13]
  wire  _T_59 = _T_48 & rowcount_4 == 32'h0; // @[ivncontrol4.scala 177:100]
  wire  _T_72 = _T_59 & rowcount_5 == 32'h0; // @[ivncontrol4.scala 180:123]
  wire  valid = _io_ProcessValid_T_2; // @[ivncontrol4.scala 153:41]
  wire [32:0] _T_91 = {{1'd0}, pin}; // @[ivncontrol4.scala 191:27]
  wire [31:0] _GEN_322 = 4'h1 == _T_91[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_323 = 4'h2 == _T_91[3:0] ? rowcount_2 : _GEN_322; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_324 = 4'h3 == _T_91[3:0] ? rowcount_3 : _GEN_323; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_325 = 4'h4 == _T_91[3:0] ? rowcount_4 : _GEN_324; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_326 = 4'h5 == _T_91[3:0] ? rowcount_5 : _GEN_325; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_327 = 4'h6 == _T_91[3:0] ? rowcount_6 : _GEN_326; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_328 = 4'h7 == _T_91[3:0] ? rowcount_7 : _GEN_327; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_329 = 4'h8 == _T_91[3:0] ? rowcount_8 : _GEN_328; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_330 = 4'h9 == _T_91[3:0] ? rowcount_9 : _GEN_329; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_331 = 4'ha == _T_91[3:0] ? rowcount_10 : _GEN_330; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_332 = 4'hb == _T_91[3:0] ? rowcount_11 : _GEN_331; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_333 = 4'hc == _T_91[3:0] ? rowcount_12 : _GEN_332; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_334 = 4'hd == _T_91[3:0] ? rowcount_13 : _GEN_333; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_335 = 4'he == _T_91[3:0] ? rowcount_14 : _GEN_334; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_336 = 4'hf == _T_91[3:0] ? rowcount_15 : _GEN_335; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_449 = _GEN_336 == 32'h1 ? _T_91[31:0] : 32'ha; // @[ivncontrol4.scala 142:17 241:50 242:21]
  wire [31:0] _GEN_450 = _GEN_336 == 32'h2 ? _T_91[31:0] : _GEN_449; // @[ivncontrol4.scala 237:51 238:21]
  wire [31:0] _GEN_451 = _GEN_336 == 32'h2 ? _T_91[31:0] : 32'h12; // @[ivncontrol4.scala 142:17 237:51 239:21]
  wire [31:0] _GEN_452 = _GEN_336 == 32'h3 ? _T_91[31:0] : _GEN_450; // @[ivncontrol4.scala 232:50 233:21]
  wire [31:0] _GEN_453 = _GEN_336 == 32'h3 ? _T_91[31:0] : _GEN_451; // @[ivncontrol4.scala 232:50 234:21]
  wire [31:0] _GEN_454 = _GEN_336 == 32'h3 ? _T_91[31:0] : 32'hd; // @[ivncontrol4.scala 142:17 232:50 235:21]
  wire [31:0] _GEN_455 = _GEN_336 == 32'h4 ? _T_91[31:0] : _GEN_452; // @[ivncontrol4.scala 224:50 225:21]
  wire [31:0] _GEN_456 = _GEN_336 == 32'h4 ? _T_91[31:0] : _GEN_453; // @[ivncontrol4.scala 224:50 226:21]
  wire [31:0] _GEN_457 = _GEN_336 == 32'h4 ? _T_91[31:0] : _GEN_454; // @[ivncontrol4.scala 224:50 227:21]
  wire [31:0] _GEN_458 = _GEN_336 == 32'h4 ? _T_91[31:0] : 32'h1b; // @[ivncontrol4.scala 142:17 224:50 228:21]
  wire [31:0] _GEN_459 = _GEN_336 == 32'h5 ? _T_91[31:0] : _GEN_455; // @[ivncontrol4.scala 217:50 218:21]
  wire [31:0] _GEN_460 = _GEN_336 == 32'h5 ? _T_91[31:0] : _GEN_456; // @[ivncontrol4.scala 217:50 219:21]
  wire [31:0] _GEN_461 = _GEN_336 == 32'h5 ? _T_91[31:0] : _GEN_457; // @[ivncontrol4.scala 217:50 220:21]
  wire [31:0] _GEN_462 = _GEN_336 == 32'h5 ? _T_91[31:0] : _GEN_458; // @[ivncontrol4.scala 217:50 221:21]
  wire [31:0] _GEN_463 = _GEN_336 == 32'h5 ? _T_91[31:0] : 32'h1a; // @[ivncontrol4.scala 143:18 217:50 222:22]
  wire [31:0] _GEN_464 = _GEN_336 == 32'h6 ? _T_91[31:0] : _GEN_459; // @[ivncontrol4.scala 209:52 210:21]
  wire [31:0] _GEN_465 = _GEN_336 == 32'h6 ? _T_91[31:0] : _GEN_460; // @[ivncontrol4.scala 209:52 211:21]
  wire [31:0] _GEN_466 = _GEN_336 == 32'h6 ? _T_91[31:0] : _GEN_461; // @[ivncontrol4.scala 209:52 212:21]
  wire [31:0] _GEN_467 = _GEN_336 == 32'h6 ? _T_91[31:0] : _GEN_462; // @[ivncontrol4.scala 209:52 213:21]
  wire [31:0] _GEN_468 = _GEN_336 == 32'h6 ? _T_91[31:0] : _GEN_463; // @[ivncontrol4.scala 209:52 214:22]
  wire [31:0] _GEN_469 = _GEN_336 == 32'h6 ? _T_91[31:0] : 32'hb; // @[ivncontrol4.scala 143:18 209:52 215:22]
  wire [31:0] _GEN_470 = _GEN_336 == 32'h7 ? _T_91[31:0] : _GEN_464; // @[ivncontrol4.scala 201:52 202:21]
  wire [31:0] _GEN_471 = _GEN_336 == 32'h7 ? _T_91[31:0] : _GEN_465; // @[ivncontrol4.scala 201:52 203:21]
  wire [31:0] _GEN_472 = _GEN_336 == 32'h7 ? _T_91[31:0] : _GEN_466; // @[ivncontrol4.scala 201:52 204:21]
  wire [31:0] _GEN_473 = _GEN_336 == 32'h7 ? _T_91[31:0] : _GEN_467; // @[ivncontrol4.scala 201:52 205:21]
  wire [31:0] _GEN_474 = _GEN_336 == 32'h7 ? _T_91[31:0] : _GEN_468; // @[ivncontrol4.scala 201:52 206:22]
  wire [31:0] _GEN_475 = _GEN_336 == 32'h7 ? _T_91[31:0] : _GEN_469; // @[ivncontrol4.scala 201:52 207:22]
  wire [31:0] _GEN_476 = _GEN_336 == 32'h7 ? _T_91[31:0] : 32'he; // @[ivncontrol4.scala 143:18 201:52 208:22]
  wire [31:0] _GEN_477 = _GEN_336 >= 32'h8 ? _T_91[31:0] : _GEN_470; // @[ivncontrol4.scala 191:42 192:21]
  wire [31:0] _GEN_478 = _GEN_336 >= 32'h8 ? _T_91[31:0] : _GEN_471; // @[ivncontrol4.scala 191:42 193:21]
  wire [31:0] _GEN_479 = _GEN_336 >= 32'h8 ? _T_91[31:0] : _GEN_472; // @[ivncontrol4.scala 191:42 194:21]
  wire [31:0] _GEN_480 = _GEN_336 >= 32'h8 ? _T_91[31:0] : _GEN_473; // @[ivncontrol4.scala 191:42 195:21]
  wire [31:0] _GEN_481 = _GEN_336 >= 32'h8 ? _T_91[31:0] : _GEN_474; // @[ivncontrol4.scala 191:42 196:22]
  wire [31:0] _GEN_482 = _GEN_336 >= 32'h8 ? _T_91[31:0] : _GEN_475; // @[ivncontrol4.scala 191:42 197:22]
  wire [31:0] _GEN_483 = _GEN_336 >= 32'h8 ? _T_91[31:0] : _GEN_476; // @[ivncontrol4.scala 191:42 198:22]
  wire [31:0] _GEN_484 = _GEN_336 >= 32'h8 ? _T_91[31:0] : 32'h13; // @[ivncontrol4.scala 143:18 191:42 199:22]
  wire [31:0] _T_127 = 32'h8 - _GEN_336; // @[ivncontrol4.scala 245:18]
  wire [31:0] _i_vn_1_T_15 = 32'h1 + pin; // @[ivncontrol4.scala 246:29]
  wire [31:0] _GEN_597 = _T_127 == 32'h1 ? _i_vn_1_T_15 : _GEN_484; // @[ivncontrol4.scala 286:54 289:22]
  wire [31:0] _GEN_598 = _T_127 == 32'h2 ? _i_vn_1_T_15 : _GEN_483; // @[ivncontrol4.scala 281:54 284:22]
  wire [31:0] _GEN_599 = _T_127 == 32'h2 ? _i_vn_1_T_15 : _GEN_597; // @[ivncontrol4.scala 281:54 285:22]
  wire [31:0] _GEN_600 = _T_127 == 32'h3 ? _i_vn_1_T_15 : _GEN_482; // @[ivncontrol4.scala 274:54 276:22]
  wire [31:0] _GEN_601 = _T_127 == 32'h3 ? _i_vn_1_T_15 : _GEN_598; // @[ivncontrol4.scala 274:54 277:22]
  wire [31:0] _GEN_602 = _T_127 == 32'h3 ? _i_vn_1_T_15 : _GEN_599; // @[ivncontrol4.scala 274:54 278:22]
  wire [31:0] _GEN_603 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_481; // @[ivncontrol4.scala 268:54 270:22]
  wire [31:0] _GEN_604 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_600; // @[ivncontrol4.scala 268:54 271:22]
  wire [31:0] _GEN_605 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_601; // @[ivncontrol4.scala 268:54 272:22]
  wire [31:0] _GEN_606 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_602; // @[ivncontrol4.scala 268:54 273:22]
  wire [31:0] _GEN_607 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_480; // @[ivncontrol4.scala 261:54 263:21]
  wire [31:0] _GEN_608 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_603; // @[ivncontrol4.scala 261:54 264:22]
  wire [31:0] _GEN_609 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_604; // @[ivncontrol4.scala 261:54 265:22]
  wire [31:0] _GEN_610 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_605; // @[ivncontrol4.scala 261:54 266:22]
  wire [31:0] _GEN_611 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_606; // @[ivncontrol4.scala 261:54 267:22]
  wire [31:0] _GEN_612 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_479; // @[ivncontrol4.scala 254:54 255:22]
  wire [31:0] _GEN_613 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_607; // @[ivncontrol4.scala 254:54 256:21]
  wire [31:0] _GEN_614 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_608; // @[ivncontrol4.scala 254:54 257:22]
  wire [31:0] _GEN_615 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_609; // @[ivncontrol4.scala 254:54 258:22]
  wire [31:0] _GEN_616 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_610; // @[ivncontrol4.scala 254:54 259:22]
  wire [31:0] _GEN_617 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_611; // @[ivncontrol4.scala 254:54 260:22]
  wire [31:0] _GEN_618 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_478; // @[ivncontrol4.scala 245:49 246:22]
  wire [31:0] _GEN_619 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_612; // @[ivncontrol4.scala 245:49 247:21]
  wire [31:0] _GEN_620 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_613; // @[ivncontrol4.scala 245:49 248:21]
  wire [31:0] _GEN_621 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_614; // @[ivncontrol4.scala 245:49 249:22]
  wire [31:0] _GEN_622 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_615; // @[ivncontrol4.scala 245:49 250:22]
  wire [31:0] _GEN_623 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_616; // @[ivncontrol4.scala 245:49 251:22]
  wire [31:0] _GEN_624 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_617; // @[ivncontrol4.scala 245:49 252:22]
  wire [31:0] _GEN_642 = 4'h1 == _i_vn_1_T_15[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_643 = 4'h2 == _i_vn_1_T_15[3:0] ? rowcount_2 : _GEN_642; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_644 = 4'h3 == _i_vn_1_T_15[3:0] ? rowcount_3 : _GEN_643; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_645 = 4'h4 == _i_vn_1_T_15[3:0] ? rowcount_4 : _GEN_644; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_646 = 4'h5 == _i_vn_1_T_15[3:0] ? rowcount_5 : _GEN_645; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_647 = 4'h6 == _i_vn_1_T_15[3:0] ? rowcount_6 : _GEN_646; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_648 = 4'h7 == _i_vn_1_T_15[3:0] ? rowcount_7 : _GEN_647; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_649 = 4'h8 == _i_vn_1_T_15[3:0] ? rowcount_8 : _GEN_648; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_650 = 4'h9 == _i_vn_1_T_15[3:0] ? rowcount_9 : _GEN_649; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_651 = 4'ha == _i_vn_1_T_15[3:0] ? rowcount_10 : _GEN_650; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_652 = 4'hb == _i_vn_1_T_15[3:0] ? rowcount_11 : _GEN_651; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_653 = 4'hc == _i_vn_1_T_15[3:0] ? rowcount_12 : _GEN_652; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_654 = 4'hd == _i_vn_1_T_15[3:0] ? rowcount_13 : _GEN_653; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_655 = 4'he == _i_vn_1_T_15[3:0] ? rowcount_14 : _GEN_654; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_656 = 4'hf == _i_vn_1_T_15[3:0] ? rowcount_15 : _GEN_655; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _T_172 = _GEN_336 + _GEN_656; // @[ivncontrol4.scala 292:41]
  wire [31:0] _T_174 = 32'h8 - _T_172; // @[ivncontrol4.scala 292:18]
  wire [31:0] _i_vn_1_T_17 = 32'h2 + pin; // @[ivncontrol4.scala 293:29]
  wire [31:0] _GEN_849 = _T_174 == 32'h1 ? _i_vn_1_T_17 : _GEN_624; // @[ivncontrol4.scala 335:78 338:22]
  wire [31:0] _GEN_850 = _T_174 == 32'h2 ? _i_vn_1_T_17 : _GEN_623; // @[ivncontrol4.scala 329:76 332:22]
  wire [31:0] _GEN_851 = _T_174 == 32'h2 ? _i_vn_1_T_17 : _GEN_849; // @[ivncontrol4.scala 329:76 333:22]
  wire [31:0] _GEN_852 = _T_174 == 32'h3 ? _i_vn_1_T_17 : _GEN_622; // @[ivncontrol4.scala 322:78 324:23]
  wire [31:0] _GEN_853 = _T_174 == 32'h3 ? _i_vn_1_T_17 : _GEN_850; // @[ivncontrol4.scala 322:78 325:22]
  wire [31:0] _GEN_854 = _T_174 == 32'h3 ? _i_vn_1_T_17 : _GEN_851; // @[ivncontrol4.scala 322:78 326:22]
  wire [31:0] _GEN_855 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_621; // @[ivncontrol4.scala 316:78 318:22]
  wire [31:0] _GEN_856 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_852; // @[ivncontrol4.scala 316:78 319:22]
  wire [31:0] _GEN_857 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_853; // @[ivncontrol4.scala 316:78 320:22]
  wire [31:0] _GEN_858 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_854; // @[ivncontrol4.scala 316:78 321:22]
  wire [31:0] _GEN_859 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_620; // @[ivncontrol4.scala 309:76 311:23]
  wire [31:0] _GEN_860 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_855; // @[ivncontrol4.scala 309:76 312:22]
  wire [31:0] _GEN_861 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_856; // @[ivncontrol4.scala 309:76 313:22]
  wire [31:0] _GEN_862 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_857; // @[ivncontrol4.scala 309:76 314:22]
  wire [31:0] _GEN_863 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_858; // @[ivncontrol4.scala 309:76 315:22]
  wire [31:0] _GEN_864 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_619; // @[ivncontrol4.scala 301:77 303:22]
  wire [31:0] _GEN_865 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_859; // @[ivncontrol4.scala 301:77 304:21]
  wire [31:0] _GEN_866 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_860; // @[ivncontrol4.scala 301:77 305:22]
  wire [31:0] _GEN_867 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_861; // @[ivncontrol4.scala 301:77 306:22]
  wire [31:0] _GEN_868 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_862; // @[ivncontrol4.scala 301:77 307:22]
  wire [31:0] _GEN_869 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_863; // @[ivncontrol4.scala 301:77 308:22]
  wire [31:0] _GEN_870 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_618; // @[ivncontrol4.scala 292:73 293:22]
  wire [31:0] _GEN_871 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_864; // @[ivncontrol4.scala 292:73 294:21]
  wire [31:0] _GEN_872 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_865; // @[ivncontrol4.scala 292:73 295:21]
  wire [31:0] _GEN_873 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_866; // @[ivncontrol4.scala 292:73 296:22]
  wire [31:0] _GEN_874 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_867; // @[ivncontrol4.scala 292:73 297:22]
  wire [31:0] _GEN_875 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_868; // @[ivncontrol4.scala 292:73 298:22]
  wire [31:0] _GEN_876 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_869; // @[ivncontrol4.scala 292:73 299:22]
  wire [31:0] _GEN_910 = 4'h1 == _i_vn_1_T_17[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_911 = 4'h2 == _i_vn_1_T_17[3:0] ? rowcount_2 : _GEN_910; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_912 = 4'h3 == _i_vn_1_T_17[3:0] ? rowcount_3 : _GEN_911; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_913 = 4'h4 == _i_vn_1_T_17[3:0] ? rowcount_4 : _GEN_912; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_914 = 4'h5 == _i_vn_1_T_17[3:0] ? rowcount_5 : _GEN_913; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_915 = 4'h6 == _i_vn_1_T_17[3:0] ? rowcount_6 : _GEN_914; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_916 = 4'h7 == _i_vn_1_T_17[3:0] ? rowcount_7 : _GEN_915; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_917 = 4'h8 == _i_vn_1_T_17[3:0] ? rowcount_8 : _GEN_916; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_918 = 4'h9 == _i_vn_1_T_17[3:0] ? rowcount_9 : _GEN_917; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_919 = 4'ha == _i_vn_1_T_17[3:0] ? rowcount_10 : _GEN_918; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_920 = 4'hb == _i_vn_1_T_17[3:0] ? rowcount_11 : _GEN_919; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_921 = 4'hc == _i_vn_1_T_17[3:0] ? rowcount_12 : _GEN_920; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_922 = 4'hd == _i_vn_1_T_17[3:0] ? rowcount_13 : _GEN_921; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_923 = 4'he == _i_vn_1_T_17[3:0] ? rowcount_14 : _GEN_922; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_924 = 4'hf == _i_vn_1_T_17[3:0] ? rowcount_15 : _GEN_923; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _T_254 = _T_172 + _GEN_924; // @[ivncontrol4.scala 343:62]
  wire [31:0] _T_256 = 32'h8 - _T_254; // @[ivncontrol4.scala 343:17]
  wire [31:0] _i_vn_1_T_19 = 32'h3 + pin; // @[ivncontrol4.scala 344:29]
  wire [31:0] _GEN_1213 = _T_256 == 32'h1 ? _i_vn_1_T_19 : _GEN_876; // @[ivncontrol4.scala 386:100 389:22]
  wire [31:0] _GEN_1214 = _T_256 == 32'h2 ? _i_vn_1_T_19 : _GEN_875; // @[ivncontrol4.scala 380:98 383:22]
  wire [31:0] _GEN_1215 = _T_256 == 32'h2 ? _i_vn_1_T_19 : _GEN_1213; // @[ivncontrol4.scala 380:98 384:22]
  wire [31:0] _GEN_1216 = _T_256 == 32'h3 ? _i_vn_1_T_19 : _GEN_874; // @[ivncontrol4.scala 373:100 375:23]
  wire [31:0] _GEN_1217 = _T_256 == 32'h3 ? _i_vn_1_T_19 : _GEN_1214; // @[ivncontrol4.scala 373:100 376:22]
  wire [31:0] _GEN_1218 = _T_256 == 32'h3 ? _i_vn_1_T_19 : _GEN_1215; // @[ivncontrol4.scala 373:100 377:22]
  wire [31:0] _GEN_1219 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_873; // @[ivncontrol4.scala 367:100 369:22]
  wire [31:0] _GEN_1220 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_1216; // @[ivncontrol4.scala 367:100 370:22]
  wire [31:0] _GEN_1221 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_1217; // @[ivncontrol4.scala 367:100 371:22]
  wire [31:0] _GEN_1222 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_1218; // @[ivncontrol4.scala 367:100 372:22]
  wire [31:0] _GEN_1223 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_872; // @[ivncontrol4.scala 360:98 362:23]
  wire [31:0] _GEN_1224 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1219; // @[ivncontrol4.scala 360:98 363:22]
  wire [31:0] _GEN_1225 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1220; // @[ivncontrol4.scala 360:98 364:22]
  wire [31:0] _GEN_1226 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1221; // @[ivncontrol4.scala 360:98 365:22]
  wire [31:0] _GEN_1227 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1222; // @[ivncontrol4.scala 360:98 366:22]
  wire [31:0] _GEN_1228 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_871; // @[ivncontrol4.scala 352:99 354:22]
  wire [31:0] _GEN_1229 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1223; // @[ivncontrol4.scala 352:99 355:21]
  wire [31:0] _GEN_1230 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1224; // @[ivncontrol4.scala 352:99 356:22]
  wire [31:0] _GEN_1231 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1225; // @[ivncontrol4.scala 352:99 357:22]
  wire [31:0] _GEN_1232 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1226; // @[ivncontrol4.scala 352:99 358:22]
  wire [31:0] _GEN_1233 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1227; // @[ivncontrol4.scala 352:99 359:22]
  wire [31:0] _GEN_1234 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_870; // @[ivncontrol4.scala 343:94 344:22]
  wire [31:0] _GEN_1235 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1228; // @[ivncontrol4.scala 343:94 345:21]
  wire [31:0] _GEN_1236 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1229; // @[ivncontrol4.scala 343:94 346:21]
  wire [31:0] _GEN_1237 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1230; // @[ivncontrol4.scala 343:94 347:22]
  wire [31:0] _GEN_1238 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1231; // @[ivncontrol4.scala 343:94 348:22]
  wire [31:0] _GEN_1239 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1232; // @[ivncontrol4.scala 343:94 349:22]
  wire [31:0] _GEN_1240 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1233; // @[ivncontrol4.scala 343:94 350:22]
  wire [31:0] _GEN_1290 = 4'h1 == _i_vn_1_T_19[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1291 = 4'h2 == _i_vn_1_T_19[3:0] ? rowcount_2 : _GEN_1290; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1292 = 4'h3 == _i_vn_1_T_19[3:0] ? rowcount_3 : _GEN_1291; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1293 = 4'h4 == _i_vn_1_T_19[3:0] ? rowcount_4 : _GEN_1292; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1294 = 4'h5 == _i_vn_1_T_19[3:0] ? rowcount_5 : _GEN_1293; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1295 = 4'h6 == _i_vn_1_T_19[3:0] ? rowcount_6 : _GEN_1294; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1296 = 4'h7 == _i_vn_1_T_19[3:0] ? rowcount_7 : _GEN_1295; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1297 = 4'h8 == _i_vn_1_T_19[3:0] ? rowcount_8 : _GEN_1296; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1298 = 4'h9 == _i_vn_1_T_19[3:0] ? rowcount_9 : _GEN_1297; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1299 = 4'ha == _i_vn_1_T_19[3:0] ? rowcount_10 : _GEN_1298; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1300 = 4'hb == _i_vn_1_T_19[3:0] ? rowcount_11 : _GEN_1299; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1301 = 4'hc == _i_vn_1_T_19[3:0] ? rowcount_12 : _GEN_1300; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1302 = 4'hd == _i_vn_1_T_19[3:0] ? rowcount_13 : _GEN_1301; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1303 = 4'he == _i_vn_1_T_19[3:0] ? rowcount_14 : _GEN_1302; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1304 = 4'hf == _i_vn_1_T_19[3:0] ? rowcount_15 : _GEN_1303; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _T_371 = _T_254 + _GEN_1304; // @[ivncontrol4.scala 393:86]
  wire [31:0] _T_373 = 32'h8 - _T_371; // @[ivncontrol4.scala 393:19]
  wire [31:0] _i_vn_1_T_21 = 32'h4 + pin; // @[ivncontrol4.scala 394:29]
  wire [31:0] _GEN_1689 = _T_373 == 32'h1 ? _i_vn_1_T_21 : _GEN_1240; // @[ivncontrol4.scala 436:122 439:22]
  wire [31:0] _GEN_1690 = _T_373 == 32'h2 ? _i_vn_1_T_21 : _GEN_1239; // @[ivncontrol4.scala 430:121 433:22]
  wire [31:0] _GEN_1691 = _T_373 == 32'h2 ? _i_vn_1_T_21 : _GEN_1689; // @[ivncontrol4.scala 430:121 434:22]
  wire [31:0] _GEN_1692 = _T_373 == 32'h3 ? _i_vn_1_T_21 : _GEN_1238; // @[ivncontrol4.scala 423:123 425:23]
  wire [31:0] _GEN_1693 = _T_373 == 32'h3 ? _i_vn_1_T_21 : _GEN_1690; // @[ivncontrol4.scala 423:123 426:22]
  wire [31:0] _GEN_1694 = _T_373 == 32'h3 ? _i_vn_1_T_21 : _GEN_1691; // @[ivncontrol4.scala 423:123 427:22]
  wire [31:0] _GEN_1695 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1237; // @[ivncontrol4.scala 417:122 419:22]
  wire [31:0] _GEN_1696 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1692; // @[ivncontrol4.scala 417:122 420:22]
  wire [31:0] _GEN_1697 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1693; // @[ivncontrol4.scala 417:122 421:22]
  wire [31:0] _GEN_1698 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1694; // @[ivncontrol4.scala 417:122 422:22]
  wire [31:0] _GEN_1699 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1236; // @[ivncontrol4.scala 410:121 412:23]
  wire [31:0] _GEN_1700 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1695; // @[ivncontrol4.scala 410:121 413:22]
  wire [31:0] _GEN_1701 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1696; // @[ivncontrol4.scala 410:121 414:22]
  wire [31:0] _GEN_1702 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1697; // @[ivncontrol4.scala 410:121 415:22]
  wire [31:0] _GEN_1703 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1698; // @[ivncontrol4.scala 410:121 416:22]
  wire [31:0] _GEN_1704 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1235; // @[ivncontrol4.scala 402:121 404:22]
  wire [31:0] _GEN_1705 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1699; // @[ivncontrol4.scala 402:121 405:21]
  wire [31:0] _GEN_1706 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1700; // @[ivncontrol4.scala 402:121 406:22]
  wire [31:0] _GEN_1707 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1701; // @[ivncontrol4.scala 402:121 407:22]
  wire [31:0] _GEN_1708 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1702; // @[ivncontrol4.scala 402:121 408:22]
  wire [31:0] _GEN_1709 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1703; // @[ivncontrol4.scala 402:121 409:22]
  wire [31:0] _GEN_1710 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1234; // @[ivncontrol4.scala 393:118 394:22]
  wire [31:0] _GEN_1711 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1704; // @[ivncontrol4.scala 393:118 395:21]
  wire [31:0] _GEN_1712 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1705; // @[ivncontrol4.scala 393:118 396:21]
  wire [31:0] _GEN_1713 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1706; // @[ivncontrol4.scala 393:118 397:22]
  wire [31:0] _GEN_1714 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1707; // @[ivncontrol4.scala 393:118 398:22]
  wire [31:0] _GEN_1715 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1708; // @[ivncontrol4.scala 393:118 399:22]
  wire [31:0] _GEN_1716 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1709; // @[ivncontrol4.scala 393:118 400:22]
  wire [31:0] _GEN_1782 = 4'h1 == _i_vn_1_T_21[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1783 = 4'h2 == _i_vn_1_T_21[3:0] ? rowcount_2 : _GEN_1782; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1784 = 4'h3 == _i_vn_1_T_21[3:0] ? rowcount_3 : _GEN_1783; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1785 = 4'h4 == _i_vn_1_T_21[3:0] ? rowcount_4 : _GEN_1784; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1786 = 4'h5 == _i_vn_1_T_21[3:0] ? rowcount_5 : _GEN_1785; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1787 = 4'h6 == _i_vn_1_T_21[3:0] ? rowcount_6 : _GEN_1786; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1788 = 4'h7 == _i_vn_1_T_21[3:0] ? rowcount_7 : _GEN_1787; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1789 = 4'h8 == _i_vn_1_T_21[3:0] ? rowcount_8 : _GEN_1788; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1790 = 4'h9 == _i_vn_1_T_21[3:0] ? rowcount_9 : _GEN_1789; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1791 = 4'ha == _i_vn_1_T_21[3:0] ? rowcount_10 : _GEN_1790; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1792 = 4'hb == _i_vn_1_T_21[3:0] ? rowcount_11 : _GEN_1791; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1793 = 4'hc == _i_vn_1_T_21[3:0] ? rowcount_12 : _GEN_1792; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1794 = 4'hd == _i_vn_1_T_21[3:0] ? rowcount_13 : _GEN_1793; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1795 = 4'he == _i_vn_1_T_21[3:0] ? rowcount_14 : _GEN_1794; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1796 = 4'hf == _i_vn_1_T_21[3:0] ? rowcount_15 : _GEN_1795; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _T_523 = _T_371 + _GEN_1796; // @[ivncontrol4.scala 443:108]
  wire [31:0] _T_525 = 32'h8 - _T_523; // @[ivncontrol4.scala 443:19]
  wire [31:0] _i_vn_1_T_23 = 32'h5 + pin; // @[ivncontrol4.scala 444:29]
  wire [31:0] _GEN_2277 = _T_525 == 32'h1 ? _i_vn_1_T_23 : _GEN_1716; // @[ivncontrol4.scala 486:144 489:22]
  wire [31:0] _GEN_2278 = _T_525 == 32'h2 ? _i_vn_1_T_23 : _GEN_1715; // @[ivncontrol4.scala 480:143 483:22]
  wire [31:0] _GEN_2279 = _T_525 == 32'h2 ? _i_vn_1_T_23 : _GEN_2277; // @[ivncontrol4.scala 480:143 484:22]
  wire [31:0] _GEN_2280 = _T_525 == 32'h3 ? _i_vn_1_T_23 : _GEN_1714; // @[ivncontrol4.scala 473:145 475:23]
  wire [31:0] _GEN_2281 = _T_525 == 32'h3 ? _i_vn_1_T_23 : _GEN_2278; // @[ivncontrol4.scala 473:145 476:22]
  wire [31:0] _GEN_2282 = _T_525 == 32'h3 ? _i_vn_1_T_23 : _GEN_2279; // @[ivncontrol4.scala 473:145 477:22]
  wire [31:0] _GEN_2283 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_1713; // @[ivncontrol4.scala 467:143 469:22]
  wire [31:0] _GEN_2284 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_2280; // @[ivncontrol4.scala 467:143 470:22]
  wire [31:0] _GEN_2285 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_2281; // @[ivncontrol4.scala 467:143 471:22]
  wire [31:0] _GEN_2286 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_2282; // @[ivncontrol4.scala 467:143 472:22]
  wire [31:0] _GEN_2287 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_1712; // @[ivncontrol4.scala 460:143 462:23]
  wire [31:0] _GEN_2288 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2283; // @[ivncontrol4.scala 460:143 463:22]
  wire [31:0] _GEN_2289 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2284; // @[ivncontrol4.scala 460:143 464:22]
  wire [31:0] _GEN_2290 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2285; // @[ivncontrol4.scala 460:143 465:22]
  wire [31:0] _GEN_2291 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2286; // @[ivncontrol4.scala 460:143 466:22]
  wire [31:0] _GEN_2292 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_1711; // @[ivncontrol4.scala 452:143 454:22]
  wire [31:0] _GEN_2293 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2287; // @[ivncontrol4.scala 452:143 455:21]
  wire [31:0] _GEN_2294 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2288; // @[ivncontrol4.scala 452:143 456:22]
  wire [31:0] _GEN_2295 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2289; // @[ivncontrol4.scala 452:143 457:22]
  wire [31:0] _GEN_2296 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2290; // @[ivncontrol4.scala 452:143 458:22]
  wire [31:0] _GEN_2297 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2291; // @[ivncontrol4.scala 452:143 459:22]
  wire [31:0] _GEN_2298 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_1710; // @[ivncontrol4.scala 443:140 444:22]
  wire [31:0] _GEN_2299 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2292; // @[ivncontrol4.scala 443:140 445:21]
  wire [31:0] _GEN_2300 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2293; // @[ivncontrol4.scala 443:140 446:21]
  wire [31:0] _GEN_2301 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2294; // @[ivncontrol4.scala 443:140 447:22]
  wire [31:0] _GEN_2302 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2295; // @[ivncontrol4.scala 443:140 448:22]
  wire [31:0] _GEN_2303 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2296; // @[ivncontrol4.scala 443:140 449:22]
  wire [31:0] _GEN_2304 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2297; // @[ivncontrol4.scala 443:140 450:22]
  wire [31:0] _GEN_2386 = 4'h1 == _i_vn_1_T_23[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2387 = 4'h2 == _i_vn_1_T_23[3:0] ? rowcount_2 : _GEN_2386; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2388 = 4'h3 == _i_vn_1_T_23[3:0] ? rowcount_3 : _GEN_2387; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2389 = 4'h4 == _i_vn_1_T_23[3:0] ? rowcount_4 : _GEN_2388; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2390 = 4'h5 == _i_vn_1_T_23[3:0] ? rowcount_5 : _GEN_2389; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2391 = 4'h6 == _i_vn_1_T_23[3:0] ? rowcount_6 : _GEN_2390; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2392 = 4'h7 == _i_vn_1_T_23[3:0] ? rowcount_7 : _GEN_2391; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2393 = 4'h8 == _i_vn_1_T_23[3:0] ? rowcount_8 : _GEN_2392; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2394 = 4'h9 == _i_vn_1_T_23[3:0] ? rowcount_9 : _GEN_2393; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2395 = 4'ha == _i_vn_1_T_23[3:0] ? rowcount_10 : _GEN_2394; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2396 = 4'hb == _i_vn_1_T_23[3:0] ? rowcount_11 : _GEN_2395; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2397 = 4'hc == _i_vn_1_T_23[3:0] ? rowcount_12 : _GEN_2396; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2398 = 4'hd == _i_vn_1_T_23[3:0] ? rowcount_13 : _GEN_2397; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2399 = 4'he == _i_vn_1_T_23[3:0] ? rowcount_14 : _GEN_2398; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2400 = 4'hf == _i_vn_1_T_23[3:0] ? rowcount_15 : _GEN_2399; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _T_710 = _T_523 + _GEN_2400; // @[ivncontrol4.scala 494:130]
  wire [31:0] _T_712 = 32'h8 - _T_710; // @[ivncontrol4.scala 494:19]
  wire [31:0] _i_vn_1_T_25 = 32'h6 + pin; // @[ivncontrol4.scala 495:29]
  wire [31:0] _GEN_2977 = _T_712 == 32'h1 ? _i_vn_1_T_25 : _GEN_2304; // @[ivncontrol4.scala 537:166 540:22]
  wire [31:0] _GEN_2978 = _T_712 == 32'h2 ? _i_vn_1_T_25 : _GEN_2303; // @[ivncontrol4.scala 531:166 534:22]
  wire [31:0] _GEN_2979 = _T_712 == 32'h2 ? _i_vn_1_T_25 : _GEN_2977; // @[ivncontrol4.scala 531:166 535:22]
  wire [31:0] _GEN_2980 = _T_712 == 32'h3 ? _i_vn_1_T_25 : _GEN_2302; // @[ivncontrol4.scala 524:168 526:23]
  wire [31:0] _GEN_2981 = _T_712 == 32'h3 ? _i_vn_1_T_25 : _GEN_2978; // @[ivncontrol4.scala 524:168 527:22]
  wire [31:0] _GEN_2982 = _T_712 == 32'h3 ? _i_vn_1_T_25 : _GEN_2979; // @[ivncontrol4.scala 524:168 528:22]
  wire [31:0] _GEN_2983 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2301; // @[ivncontrol4.scala 518:166 520:22]
  wire [31:0] _GEN_2984 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2980; // @[ivncontrol4.scala 518:166 521:22]
  wire [31:0] _GEN_2985 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2981; // @[ivncontrol4.scala 518:166 522:22]
  wire [31:0] _GEN_2986 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2982; // @[ivncontrol4.scala 518:166 523:22]
  wire [31:0] _GEN_2987 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2300; // @[ivncontrol4.scala 511:166 513:23]
  wire [31:0] _GEN_2988 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2983; // @[ivncontrol4.scala 511:166 514:22]
  wire [31:0] _GEN_2989 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2984; // @[ivncontrol4.scala 511:166 515:22]
  wire [31:0] _GEN_2990 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2985; // @[ivncontrol4.scala 511:166 516:22]
  wire [31:0] _GEN_2991 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2986; // @[ivncontrol4.scala 511:166 517:22]
  wire [31:0] _GEN_2992 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2299; // @[ivncontrol4.scala 503:166 505:22]
  wire [31:0] _GEN_2993 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2987; // @[ivncontrol4.scala 503:166 506:21]
  wire [31:0] _GEN_2994 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2988; // @[ivncontrol4.scala 503:166 507:22]
  wire [31:0] _GEN_2995 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2989; // @[ivncontrol4.scala 503:166 508:22]
  wire [31:0] _GEN_2996 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2990; // @[ivncontrol4.scala 503:166 509:22]
  wire [31:0] _GEN_2997 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2991; // @[ivncontrol4.scala 503:166 510:22]
  wire [31:0] _GEN_2998 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2298; // @[ivncontrol4.scala 494:162 495:22]
  wire [31:0] _GEN_2999 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2992; // @[ivncontrol4.scala 494:162 496:21]
  wire [31:0] _GEN_3000 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2993; // @[ivncontrol4.scala 494:162 497:21]
  wire [31:0] _GEN_3001 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2994; // @[ivncontrol4.scala 494:162 498:22]
  wire [31:0] _GEN_3002 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2995; // @[ivncontrol4.scala 494:162 499:22]
  wire [31:0] _GEN_3003 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2996; // @[ivncontrol4.scala 494:162 500:22]
  wire [31:0] _GEN_3004 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2997; // @[ivncontrol4.scala 494:162 501:22]
  wire [31:0] _GEN_3102 = 4'h1 == _i_vn_1_T_25[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3103 = 4'h2 == _i_vn_1_T_25[3:0] ? rowcount_2 : _GEN_3102; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3104 = 4'h3 == _i_vn_1_T_25[3:0] ? rowcount_3 : _GEN_3103; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3105 = 4'h4 == _i_vn_1_T_25[3:0] ? rowcount_4 : _GEN_3104; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3106 = 4'h5 == _i_vn_1_T_25[3:0] ? rowcount_5 : _GEN_3105; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3107 = 4'h6 == _i_vn_1_T_25[3:0] ? rowcount_6 : _GEN_3106; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3108 = 4'h7 == _i_vn_1_T_25[3:0] ? rowcount_7 : _GEN_3107; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3109 = 4'h8 == _i_vn_1_T_25[3:0] ? rowcount_8 : _GEN_3108; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3110 = 4'h9 == _i_vn_1_T_25[3:0] ? rowcount_9 : _GEN_3109; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3111 = 4'ha == _i_vn_1_T_25[3:0] ? rowcount_10 : _GEN_3110; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3112 = 4'hb == _i_vn_1_T_25[3:0] ? rowcount_11 : _GEN_3111; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3113 = 4'hc == _i_vn_1_T_25[3:0] ? rowcount_12 : _GEN_3112; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3114 = 4'hd == _i_vn_1_T_25[3:0] ? rowcount_13 : _GEN_3113; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3115 = 4'he == _i_vn_1_T_25[3:0] ? rowcount_14 : _GEN_3114; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3116 = 4'hf == _i_vn_1_T_25[3:0] ? rowcount_15 : _GEN_3115; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _T_932 = _T_710 + _GEN_3116; // @[ivncontrol4.scala 545:152]
  wire [31:0] _T_934 = 32'h8 - _T_932; // @[ivncontrol4.scala 545:19]
  wire [31:0] _i_vn_1_T_27 = 32'h7 + pin; // @[ivncontrol4.scala 546:29]
  wire [31:0] _GEN_3789 = _T_934 == 32'h1 ? _i_vn_1_T_27 : _GEN_3004; // @[ivncontrol4.scala 588:188 591:22]
  wire [31:0] _GEN_3790 = _T_934 == 32'h2 ? _i_vn_1_T_27 : _GEN_3003; // @[ivncontrol4.scala 582:188 585:22]
  wire [31:0] _GEN_3791 = _T_934 == 32'h2 ? _i_vn_1_T_27 : _GEN_3789; // @[ivncontrol4.scala 582:188 586:22]
  wire [31:0] _GEN_3792 = _T_934 == 32'h3 ? _i_vn_1_T_27 : _GEN_3002; // @[ivncontrol4.scala 575:190 577:23]
  wire [31:0] _GEN_3793 = _T_934 == 32'h3 ? _i_vn_1_T_27 : _GEN_3790; // @[ivncontrol4.scala 575:190 578:22]
  wire [31:0] _GEN_3794 = _T_934 == 32'h3 ? _i_vn_1_T_27 : _GEN_3791; // @[ivncontrol4.scala 575:190 579:22]
  wire [31:0] _GEN_3795 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_3001; // @[ivncontrol4.scala 569:188 571:22]
  wire [31:0] _GEN_3796 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_3792; // @[ivncontrol4.scala 569:188 572:22]
  wire [31:0] _GEN_3797 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_3793; // @[ivncontrol4.scala 569:188 573:22]
  wire [31:0] _GEN_3798 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_3794; // @[ivncontrol4.scala 569:188 574:22]
  wire [31:0] _GEN_3799 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3000; // @[ivncontrol4.scala 562:188 564:23]
  wire [31:0] _GEN_3800 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3795; // @[ivncontrol4.scala 562:188 565:22]
  wire [31:0] _GEN_3801 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3796; // @[ivncontrol4.scala 562:188 566:22]
  wire [31:0] _GEN_3802 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3797; // @[ivncontrol4.scala 562:188 567:22]
  wire [31:0] _GEN_3803 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3798; // @[ivncontrol4.scala 562:188 568:22]
  wire [31:0] _GEN_3804 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_2999; // @[ivncontrol4.scala 554:188 556:22]
  wire [31:0] _GEN_3805 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3799; // @[ivncontrol4.scala 554:188 557:21]
  wire [31:0] _GEN_3806 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3800; // @[ivncontrol4.scala 554:188 558:22]
  wire [31:0] _GEN_3807 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3801; // @[ivncontrol4.scala 554:188 559:22]
  wire [31:0] _GEN_3808 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3802; // @[ivncontrol4.scala 554:188 560:22]
  wire [31:0] _GEN_3809 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3803; // @[ivncontrol4.scala 554:188 561:22]
  wire [31:0] _GEN_3810 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_2998; // @[ivncontrol4.scala 545:184 546:22]
  wire [31:0] _GEN_3811 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3804; // @[ivncontrol4.scala 545:184 547:21]
  wire [31:0] _GEN_3812 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3805; // @[ivncontrol4.scala 545:184 548:21]
  wire [31:0] _GEN_3813 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3806; // @[ivncontrol4.scala 545:184 549:22]
  wire [31:0] _GEN_3814 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3807; // @[ivncontrol4.scala 545:184 550:22]
  wire [31:0] _GEN_3815 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3808; // @[ivncontrol4.scala 545:184 551:22]
  wire [31:0] _GEN_3816 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3809; // @[ivncontrol4.scala 545:184 552:22]
  wire [31:0] _GEN_3817 = _GEN_312 ? _GEN_477 : 32'ha; // @[ivncontrol4.scala 142:17 189:28]
  wire [31:0] _GEN_3818 = _GEN_312 ? _GEN_3810 : 32'h12; // @[ivncontrol4.scala 142:17 189:28]
  wire [31:0] _GEN_3819 = _GEN_312 ? _GEN_3811 : 32'hd; // @[ivncontrol4.scala 142:17 189:28]
  wire [31:0] _GEN_3820 = _GEN_312 ? _GEN_3812 : 32'h1b; // @[ivncontrol4.scala 142:17 189:28]
  wire [31:0] _GEN_3821 = _GEN_312 ? _GEN_3813 : 32'h1a; // @[ivncontrol4.scala 143:18 189:28]
  wire [31:0] _GEN_3822 = _GEN_312 ? _GEN_3814 : 32'hb; // @[ivncontrol4.scala 143:18 189:28]
  wire [31:0] _GEN_3823 = _GEN_312 ? _GEN_3815 : 32'he; // @[ivncontrol4.scala 143:18 189:28]
  wire [31:0] _GEN_3824 = _GEN_312 ? _GEN_3816 : 32'h13; // @[ivncontrol4.scala 143:18 189:28]
  wire  valid1 = 1'h0;
  wire [31:0] _GEN_4221 = reset ? 32'h0 : _GEN_3817; // @[ivncontrol4.scala 17:{23,23}]
  wire [31:0] _GEN_4222 = reset ? 32'h0 : _GEN_3818; // @[ivncontrol4.scala 17:{23,23}]
  wire [31:0] _GEN_4223 = reset ? 32'h0 : _GEN_3819; // @[ivncontrol4.scala 17:{23,23}]
  wire [31:0] _GEN_4224 = reset ? 32'h0 : _GEN_3820; // @[ivncontrol4.scala 17:{23,23}]
  wire [31:0] _GEN_4225 = reset ? 32'h0 : _GEN_3821; // @[ivncontrol4.scala 18:{24,24}]
  wire [31:0] _GEN_4226 = reset ? 32'h0 : _GEN_3822; // @[ivncontrol4.scala 18:{24,24}]
  wire [31:0] _GEN_4227 = reset ? 32'h0 : _GEN_3823; // @[ivncontrol4.scala 18:{24,24}]
  wire [31:0] _GEN_4228 = reset ? 32'h0 : _GEN_3824; // @[ivncontrol4.scala 18:{24,24}]
  assign io_o_vn_0 = i_vn_0; // @[ivncontrol4.scala 138:13]
  assign io_o_vn_1 = i_vn_1; // @[ivncontrol4.scala 138:13]
  assign io_o_vn_2 = i_vn_2; // @[ivncontrol4.scala 138:13]
  assign io_o_vn_3 = i_vn_3; // @[ivncontrol4.scala 138:13]
  assign io_o_vn2_0 = i_vn2_0; // @[ivncontrol4.scala 139:14]
  assign io_o_vn2_1 = i_vn2_1; // @[ivncontrol4.scala 139:14]
  assign io_o_vn2_2 = i_vn2_2; // @[ivncontrol4.scala 139:14]
  assign io_o_vn2_3 = i_vn2_3; // @[ivncontrol4.scala 139:14]
  always @(posedge clock) begin
    i_vn_0 <= _GEN_4221[4:0]; // @[ivncontrol4.scala 17:{23,23}]
    i_vn_1 <= _GEN_4222[4:0]; // @[ivncontrol4.scala 17:{23,23}]
    i_vn_2 <= _GEN_4223[4:0]; // @[ivncontrol4.scala 17:{23,23}]
    i_vn_3 <= _GEN_4224[4:0]; // @[ivncontrol4.scala 17:{23,23}]
    i_vn2_0 <= _GEN_4225[4:0]; // @[ivncontrol4.scala 18:{24,24}]
    i_vn2_1 <= _GEN_4226[4:0]; // @[ivncontrol4.scala 18:{24,24}]
    i_vn2_2 <= _GEN_4227[4:0]; // @[ivncontrol4.scala 18:{24,24}]
    i_vn2_3 <= _GEN_4228[4:0]; // @[ivncontrol4.scala 18:{24,24}]
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_0 <= io_Stationary_matrix_0_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_1 <= io_Stationary_matrix_0_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_2 <= io_Stationary_matrix_0_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_3 <= io_Stationary_matrix_0_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_4 <= io_Stationary_matrix_0_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_5 <= io_Stationary_matrix_0_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_6 <= io_Stationary_matrix_0_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_7 <= io_Stationary_matrix_0_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_0 <= io_Stationary_matrix_1_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_1 <= io_Stationary_matrix_1_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_2 <= io_Stationary_matrix_1_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_3 <= io_Stationary_matrix_1_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_4 <= io_Stationary_matrix_1_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_5 <= io_Stationary_matrix_1_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_6 <= io_Stationary_matrix_1_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_7 <= io_Stationary_matrix_1_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_0 <= io_Stationary_matrix_2_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_1 <= io_Stationary_matrix_2_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_2 <= io_Stationary_matrix_2_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_3 <= io_Stationary_matrix_2_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_4 <= io_Stationary_matrix_2_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_5 <= io_Stationary_matrix_2_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_6 <= io_Stationary_matrix_2_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_7 <= io_Stationary_matrix_2_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_0 <= io_Stationary_matrix_3_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_1 <= io_Stationary_matrix_3_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_2 <= io_Stationary_matrix_3_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_3 <= io_Stationary_matrix_3_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_4 <= io_Stationary_matrix_3_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_5 <= io_Stationary_matrix_3_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_6 <= io_Stationary_matrix_3_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_7 <= io_Stationary_matrix_3_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_0 <= io_Stationary_matrix_4_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_1 <= io_Stationary_matrix_4_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_2 <= io_Stationary_matrix_4_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_3 <= io_Stationary_matrix_4_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_4 <= io_Stationary_matrix_4_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_5 <= io_Stationary_matrix_4_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_6 <= io_Stationary_matrix_4_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_7 <= io_Stationary_matrix_4_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_0 <= io_Stationary_matrix_5_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_1 <= io_Stationary_matrix_5_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_2 <= io_Stationary_matrix_5_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_3 <= io_Stationary_matrix_5_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_4 <= io_Stationary_matrix_5_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_5 <= io_Stationary_matrix_5_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_6 <= io_Stationary_matrix_5_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_7 <= io_Stationary_matrix_5_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_0 <= io_Stationary_matrix_6_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_1 <= io_Stationary_matrix_6_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_2 <= io_Stationary_matrix_6_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_3 <= io_Stationary_matrix_6_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_4 <= io_Stationary_matrix_6_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_5 <= io_Stationary_matrix_6_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_6 <= io_Stationary_matrix_6_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_7 <= io_Stationary_matrix_6_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_0 <= io_Stationary_matrix_7_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_1 <= io_Stationary_matrix_7_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_2 <= io_Stationary_matrix_7_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_3 <= io_Stationary_matrix_7_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_4 <= io_Stationary_matrix_7_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_5 <= io_Stationary_matrix_7_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_6 <= io_Stationary_matrix_7_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_7 <= io_Stationary_matrix_7_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_0 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_0 <= count_0; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_1 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_1 <= count_1; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_2 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_2 <= count_2; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_3 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_3 <= count_3; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_4 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_4 <= count_4; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_5 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_5 <= count_5; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_6 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_6 <= count_6; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_7 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_7 <= count_7; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_8 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_8 <= 32'h0; // @[ivncontrol4.scala 87:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_9 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_9 <= 32'h0; // @[ivncontrol4.scala 87:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_10 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_10 <= 32'h0; // @[ivncontrol4.scala 87:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_11 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_11 <= 32'h0; // @[ivncontrol4.scala 87:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_12 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_12 <= 32'h0; // @[ivncontrol4.scala 87:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_13 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_13 <= 32'h0; // @[ivncontrol4.scala 87:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_14 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_14 <= 32'h0; // @[ivncontrol4.scala 87:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_15 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end
    if (reset) begin // @[ivncontrol4.scala 37:22]
      pin <= 32'h0; // @[ivncontrol4.scala 37:22]
    end else if (_T_72 & rowcount_6 == 32'h0 & rowcount_7 != 32'h0) begin // @[ivncontrol4.scala 183:192]
      pin <= 32'h7; // @[ivncontrol4.scala 184:13]
    end else if (_T_59 & rowcount_5 == 32'h0 & rowcount_6 != 32'h0) begin // @[ivncontrol4.scala 180:169]
      pin <= 32'h6; // @[ivncontrol4.scala 181:13]
    end else if (_T_48 & rowcount_4 == 32'h0 & rowcount_5 != 32'h0) begin // @[ivncontrol4.scala 177:146]
      pin <= 32'h5; // @[ivncontrol4.scala 178:13]
    end else begin
      pin <= _GEN_317;
    end
    if (reset) begin // @[ivncontrol4.scala 41:20]
      i <= 32'h0; // @[ivncontrol4.scala 41:20]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
        i <= _GEN_247;
      end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
        i <= _GEN_247;
      end else begin
        i <= _GEN_265;
      end
    end
    if (reset) begin // @[ivncontrol4.scala 42:20]
      j <= 32'h0; // @[ivncontrol4.scala 42:20]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
        j <= 32'h8; // @[ivncontrol4.scala 116:11]
      end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
        j <= _j_T_1; // @[ivncontrol4.scala 118:11]
      end else begin
        j <= {{28'd0}, _GEN_264};
      end
    end
    if (3'h0 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h0 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h0 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h0 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h0 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h0 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h0 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h0 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_0 <= _GEN_224;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_0 <= _GEN_224;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h0 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_0 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_0 <= _GEN_224;
      end
    end else begin
      count_0 <= _GEN_224;
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_1 <= _GEN_225;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_1 <= _GEN_225;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h1 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_1 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_1 <= _GEN_225;
      end
    end else begin
      count_1 <= _GEN_225;
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_2 <= _GEN_226;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_2 <= _GEN_226;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h2 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_2 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_2 <= _GEN_226;
      end
    end else begin
      count_2 <= _GEN_226;
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_3 <= _GEN_227;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_3 <= _GEN_227;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h3 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_3 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_3 <= _GEN_227;
      end
    end else begin
      count_3 <= _GEN_227;
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_4 <= _GEN_228;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_4 <= _GEN_228;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h4 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_4 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_4 <= _GEN_228;
      end
    end else begin
      count_4 <= _GEN_228;
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_5 <= _GEN_229;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_5 <= _GEN_229;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h5 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_5 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_5 <= _GEN_229;
      end
    end else begin
      count_5 <= _GEN_229;
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_6 <= _GEN_230;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_6 <= _GEN_230;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h6 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_6 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_6 <= _GEN_230;
      end
    end else begin
      count_6 <= _GEN_230;
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_7 <= _GEN_231;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_7 <= _GEN_231;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h7 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_7 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_7 <= _GEN_231;
      end
    end else begin
      count_7 <= _GEN_231;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  i_vn_0 = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  i_vn_1 = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  i_vn_2 = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  i_vn_3 = _RAND_3[4:0];
  _RAND_4 = {1{`RANDOM}};
  i_vn2_0 = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  i_vn2_1 = _RAND_5[4:0];
  _RAND_6 = {1{`RANDOM}};
  i_vn2_2 = _RAND_6[4:0];
  _RAND_7 = {1{`RANDOM}};
  i_vn2_3 = _RAND_7[4:0];
  _RAND_8 = {1{`RANDOM}};
  solution_0_0 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  solution_0_1 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  solution_0_2 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  solution_0_3 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  solution_0_4 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  solution_0_5 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  solution_0_6 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  solution_0_7 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  solution_1_0 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  solution_1_1 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  solution_1_2 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  solution_1_3 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  solution_1_4 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  solution_1_5 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  solution_1_6 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  solution_1_7 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  solution_2_0 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  solution_2_1 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  solution_2_2 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  solution_2_3 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  solution_2_4 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  solution_2_5 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  solution_2_6 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  solution_2_7 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  solution_3_0 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  solution_3_1 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  solution_3_2 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  solution_3_3 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  solution_3_4 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  solution_3_5 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  solution_3_6 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  solution_3_7 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  solution_4_0 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  solution_4_1 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  solution_4_2 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  solution_4_3 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  solution_4_4 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  solution_4_5 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  solution_4_6 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  solution_4_7 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  solution_5_0 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  solution_5_1 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  solution_5_2 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  solution_5_3 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  solution_5_4 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  solution_5_5 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  solution_5_6 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  solution_5_7 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  solution_6_0 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  solution_6_1 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  solution_6_2 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  solution_6_3 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  solution_6_4 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  solution_6_5 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  solution_6_6 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  solution_6_7 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  solution_7_0 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  solution_7_1 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  solution_7_2 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  solution_7_3 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  solution_7_4 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  solution_7_5 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  solution_7_6 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  solution_7_7 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  rowcount_0 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  rowcount_1 = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  rowcount_2 = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  rowcount_3 = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  rowcount_4 = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  rowcount_5 = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  rowcount_6 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  rowcount_7 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  rowcount_8 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  rowcount_9 = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  rowcount_10 = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  rowcount_11 = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  rowcount_12 = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  rowcount_13 = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  rowcount_14 = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  rowcount_15 = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  pin = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  i = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  j = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  mat_0_0 = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  mat_0_1 = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  mat_0_2 = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  mat_0_3 = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  mat_0_4 = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  mat_0_5 = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  mat_0_6 = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  mat_0_7 = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  mat_1_0 = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  mat_1_1 = _RAND_100[31:0];
  _RAND_101 = {1{`RANDOM}};
  mat_1_2 = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  mat_1_3 = _RAND_102[31:0];
  _RAND_103 = {1{`RANDOM}};
  mat_1_4 = _RAND_103[31:0];
  _RAND_104 = {1{`RANDOM}};
  mat_1_5 = _RAND_104[31:0];
  _RAND_105 = {1{`RANDOM}};
  mat_1_6 = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  mat_1_7 = _RAND_106[31:0];
  _RAND_107 = {1{`RANDOM}};
  mat_2_0 = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  mat_2_1 = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  mat_2_2 = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  mat_2_3 = _RAND_110[31:0];
  _RAND_111 = {1{`RANDOM}};
  mat_2_4 = _RAND_111[31:0];
  _RAND_112 = {1{`RANDOM}};
  mat_2_5 = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  mat_2_6 = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  mat_2_7 = _RAND_114[31:0];
  _RAND_115 = {1{`RANDOM}};
  mat_3_0 = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  mat_3_1 = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  mat_3_2 = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  mat_3_3 = _RAND_118[31:0];
  _RAND_119 = {1{`RANDOM}};
  mat_3_4 = _RAND_119[31:0];
  _RAND_120 = {1{`RANDOM}};
  mat_3_5 = _RAND_120[31:0];
  _RAND_121 = {1{`RANDOM}};
  mat_3_6 = _RAND_121[31:0];
  _RAND_122 = {1{`RANDOM}};
  mat_3_7 = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  mat_4_0 = _RAND_123[31:0];
  _RAND_124 = {1{`RANDOM}};
  mat_4_1 = _RAND_124[31:0];
  _RAND_125 = {1{`RANDOM}};
  mat_4_2 = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  mat_4_3 = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  mat_4_4 = _RAND_127[31:0];
  _RAND_128 = {1{`RANDOM}};
  mat_4_5 = _RAND_128[31:0];
  _RAND_129 = {1{`RANDOM}};
  mat_4_6 = _RAND_129[31:0];
  _RAND_130 = {1{`RANDOM}};
  mat_4_7 = _RAND_130[31:0];
  _RAND_131 = {1{`RANDOM}};
  mat_5_0 = _RAND_131[31:0];
  _RAND_132 = {1{`RANDOM}};
  mat_5_1 = _RAND_132[31:0];
  _RAND_133 = {1{`RANDOM}};
  mat_5_2 = _RAND_133[31:0];
  _RAND_134 = {1{`RANDOM}};
  mat_5_3 = _RAND_134[31:0];
  _RAND_135 = {1{`RANDOM}};
  mat_5_4 = _RAND_135[31:0];
  _RAND_136 = {1{`RANDOM}};
  mat_5_5 = _RAND_136[31:0];
  _RAND_137 = {1{`RANDOM}};
  mat_5_6 = _RAND_137[31:0];
  _RAND_138 = {1{`RANDOM}};
  mat_5_7 = _RAND_138[31:0];
  _RAND_139 = {1{`RANDOM}};
  mat_6_0 = _RAND_139[31:0];
  _RAND_140 = {1{`RANDOM}};
  mat_6_1 = _RAND_140[31:0];
  _RAND_141 = {1{`RANDOM}};
  mat_6_2 = _RAND_141[31:0];
  _RAND_142 = {1{`RANDOM}};
  mat_6_3 = _RAND_142[31:0];
  _RAND_143 = {1{`RANDOM}};
  mat_6_4 = _RAND_143[31:0];
  _RAND_144 = {1{`RANDOM}};
  mat_6_5 = _RAND_144[31:0];
  _RAND_145 = {1{`RANDOM}};
  mat_6_6 = _RAND_145[31:0];
  _RAND_146 = {1{`RANDOM}};
  mat_6_7 = _RAND_146[31:0];
  _RAND_147 = {1{`RANDOM}};
  mat_7_0 = _RAND_147[31:0];
  _RAND_148 = {1{`RANDOM}};
  mat_7_1 = _RAND_148[31:0];
  _RAND_149 = {1{`RANDOM}};
  mat_7_2 = _RAND_149[31:0];
  _RAND_150 = {1{`RANDOM}};
  mat_7_3 = _RAND_150[31:0];
  _RAND_151 = {1{`RANDOM}};
  mat_7_4 = _RAND_151[31:0];
  _RAND_152 = {1{`RANDOM}};
  mat_7_5 = _RAND_152[31:0];
  _RAND_153 = {1{`RANDOM}};
  mat_7_6 = _RAND_153[31:0];
  _RAND_154 = {1{`RANDOM}};
  mat_7_7 = _RAND_154[31:0];
  _RAND_155 = {1{`RANDOM}};
  count_0 = _RAND_155[31:0];
  _RAND_156 = {1{`RANDOM}};
  count_1 = _RAND_156[31:0];
  _RAND_157 = {1{`RANDOM}};
  count_2 = _RAND_157[31:0];
  _RAND_158 = {1{`RANDOM}};
  count_3 = _RAND_158[31:0];
  _RAND_159 = {1{`RANDOM}};
  count_4 = _RAND_159[31:0];
  _RAND_160 = {1{`RANDOM}};
  count_5 = _RAND_160[31:0];
  _RAND_161 = {1{`RANDOM}};
  count_6 = _RAND_161[31:0];
  _RAND_162 = {1{`RANDOM}};
  count_7 = _RAND_162[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ivncontrol4_6(
  input         clock,
  input         reset,
  input  [15:0] io_Stationary_matrix_0_0,
  input  [15:0] io_Stationary_matrix_0_1,
  input  [15:0] io_Stationary_matrix_0_2,
  input  [15:0] io_Stationary_matrix_0_3,
  input  [15:0] io_Stationary_matrix_0_4,
  input  [15:0] io_Stationary_matrix_0_5,
  input  [15:0] io_Stationary_matrix_0_6,
  input  [15:0] io_Stationary_matrix_0_7,
  input  [15:0] io_Stationary_matrix_1_0,
  input  [15:0] io_Stationary_matrix_1_1,
  input  [15:0] io_Stationary_matrix_1_2,
  input  [15:0] io_Stationary_matrix_1_3,
  input  [15:0] io_Stationary_matrix_1_4,
  input  [15:0] io_Stationary_matrix_1_5,
  input  [15:0] io_Stationary_matrix_1_6,
  input  [15:0] io_Stationary_matrix_1_7,
  input  [15:0] io_Stationary_matrix_2_0,
  input  [15:0] io_Stationary_matrix_2_1,
  input  [15:0] io_Stationary_matrix_2_2,
  input  [15:0] io_Stationary_matrix_2_3,
  input  [15:0] io_Stationary_matrix_2_4,
  input  [15:0] io_Stationary_matrix_2_5,
  input  [15:0] io_Stationary_matrix_2_6,
  input  [15:0] io_Stationary_matrix_2_7,
  input  [15:0] io_Stationary_matrix_3_0,
  input  [15:0] io_Stationary_matrix_3_1,
  input  [15:0] io_Stationary_matrix_3_2,
  input  [15:0] io_Stationary_matrix_3_3,
  input  [15:0] io_Stationary_matrix_3_4,
  input  [15:0] io_Stationary_matrix_3_5,
  input  [15:0] io_Stationary_matrix_3_6,
  input  [15:0] io_Stationary_matrix_3_7,
  input  [15:0] io_Stationary_matrix_4_0,
  input  [15:0] io_Stationary_matrix_4_1,
  input  [15:0] io_Stationary_matrix_4_2,
  input  [15:0] io_Stationary_matrix_4_3,
  input  [15:0] io_Stationary_matrix_4_4,
  input  [15:0] io_Stationary_matrix_4_5,
  input  [15:0] io_Stationary_matrix_4_6,
  input  [15:0] io_Stationary_matrix_4_7,
  input  [15:0] io_Stationary_matrix_5_0,
  input  [15:0] io_Stationary_matrix_5_1,
  input  [15:0] io_Stationary_matrix_5_2,
  input  [15:0] io_Stationary_matrix_5_3,
  input  [15:0] io_Stationary_matrix_5_4,
  input  [15:0] io_Stationary_matrix_5_5,
  input  [15:0] io_Stationary_matrix_5_6,
  input  [15:0] io_Stationary_matrix_5_7,
  input  [15:0] io_Stationary_matrix_6_0,
  input  [15:0] io_Stationary_matrix_6_1,
  input  [15:0] io_Stationary_matrix_6_2,
  input  [15:0] io_Stationary_matrix_6_3,
  input  [15:0] io_Stationary_matrix_6_4,
  input  [15:0] io_Stationary_matrix_6_5,
  input  [15:0] io_Stationary_matrix_6_6,
  input  [15:0] io_Stationary_matrix_6_7,
  input  [15:0] io_Stationary_matrix_7_0,
  input  [15:0] io_Stationary_matrix_7_1,
  input  [15:0] io_Stationary_matrix_7_2,
  input  [15:0] io_Stationary_matrix_7_3,
  input  [15:0] io_Stationary_matrix_7_4,
  input  [15:0] io_Stationary_matrix_7_5,
  input  [15:0] io_Stationary_matrix_7_6,
  input  [15:0] io_Stationary_matrix_7_7,
  output [4:0]  io_o_vn_0,
  output [4:0]  io_o_vn_1,
  output [4:0]  io_o_vn_2,
  output [4:0]  io_o_vn_3,
  output [4:0]  io_o_vn2_0,
  output [4:0]  io_o_vn2_1,
  output [4:0]  io_o_vn2_2,
  output [4:0]  io_o_vn2_3,
  input         io_validpin
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
`endif // RANDOMIZE_REG_INIT
  reg [4:0] i_vn_0; // @[ivncontrol4.scala 17:23]
  reg [4:0] i_vn_1; // @[ivncontrol4.scala 17:23]
  reg [4:0] i_vn_2; // @[ivncontrol4.scala 17:23]
  reg [4:0] i_vn_3; // @[ivncontrol4.scala 17:23]
  reg [4:0] i_vn2_0; // @[ivncontrol4.scala 18:24]
  reg [4:0] i_vn2_1; // @[ivncontrol4.scala 18:24]
  reg [4:0] i_vn2_2; // @[ivncontrol4.scala 18:24]
  reg [4:0] i_vn2_3; // @[ivncontrol4.scala 18:24]
  reg [15:0] solution_0_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_0_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_0_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_0_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_0_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_0_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_0_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_0_7; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_7; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_7; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_7; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_7; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_7; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_7; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_7; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_0; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_1; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_2; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_3; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_4; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_5; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_6; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_7; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_8; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_9; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_10; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_11; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_12; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_13; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_14; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_15; // @[ivncontrol4.scala 27:27]
  reg [31:0] pin; // @[ivncontrol4.scala 37:22]
  reg [31:0] i; // @[ivncontrol4.scala 41:20]
  reg [31:0] j; // @[ivncontrol4.scala 42:20]
  wire  _io_ProcessValid_T = i == 32'h7; // @[ivncontrol4.scala 44:27]
  wire  _io_ProcessValid_T_1 = j == 32'h7; // @[ivncontrol4.scala 44:42]
  wire  _io_ProcessValid_T_2 = i == 32'h7 & j == 32'h7; // @[ivncontrol4.scala 44:36]
  reg [31:0] mat_0_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_0_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_0_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_0_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_0_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_0_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_0_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_0_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] count_0; // @[ivncontrol4.scala 58:20]
  reg [31:0] count_1; // @[ivncontrol4.scala 58:20]
  reg [31:0] count_2; // @[ivncontrol4.scala 58:20]
  reg [31:0] count_3; // @[ivncontrol4.scala 58:20]
  reg [31:0] count_4; // @[ivncontrol4.scala 58:20]
  reg [31:0] count_5; // @[ivncontrol4.scala 58:20]
  reg [31:0] count_6; // @[ivncontrol4.scala 58:20]
  reg [31:0] count_7; // @[ivncontrol4.scala 58:20]
  wire  _GEN_3825 = 3'h0 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_65 = 3'h0 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_0_1 : io_Stationary_matrix_0_0; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_66 = 3'h0 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_0_2 : _GEN_65; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_67 = 3'h0 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_0_3 : _GEN_66; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_68 = 3'h0 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_0_4 : _GEN_67; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_69 = 3'h0 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_0_5 : _GEN_68; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_70 = 3'h0 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_0_6 : _GEN_69; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_71 = 3'h0 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_0_7 : _GEN_70; // @[ivncontrol4.scala 63:{17,17}]
  wire  _GEN_3839 = 3'h1 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_72 = 3'h1 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_1_0 : _GEN_71; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_73 = 3'h1 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_1_1 : _GEN_72; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_74 = 3'h1 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_1_2 : _GEN_73; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_75 = 3'h1 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_1_3 : _GEN_74; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_76 = 3'h1 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_1_4 : _GEN_75; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_77 = 3'h1 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_1_5 : _GEN_76; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_78 = 3'h1 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_1_6 : _GEN_77; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_79 = 3'h1 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_1_7 : _GEN_78; // @[ivncontrol4.scala 63:{17,17}]
  wire  _GEN_3855 = 3'h2 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_80 = 3'h2 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_2_0 : _GEN_79; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_81 = 3'h2 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_2_1 : _GEN_80; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_82 = 3'h2 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_2_2 : _GEN_81; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_83 = 3'h2 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_2_3 : _GEN_82; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_84 = 3'h2 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_2_4 : _GEN_83; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_85 = 3'h2 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_2_5 : _GEN_84; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_86 = 3'h2 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_2_6 : _GEN_85; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_87 = 3'h2 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_2_7 : _GEN_86; // @[ivncontrol4.scala 63:{17,17}]
  wire  _GEN_3871 = 3'h3 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_88 = 3'h3 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_3_0 : _GEN_87; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_89 = 3'h3 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_3_1 : _GEN_88; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_90 = 3'h3 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_3_2 : _GEN_89; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_91 = 3'h3 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_3_3 : _GEN_90; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_92 = 3'h3 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_3_4 : _GEN_91; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_93 = 3'h3 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_3_5 : _GEN_92; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_94 = 3'h3 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_3_6 : _GEN_93; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_95 = 3'h3 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_3_7 : _GEN_94; // @[ivncontrol4.scala 63:{17,17}]
  wire  _GEN_3887 = 3'h4 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_96 = 3'h4 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_4_0 : _GEN_95; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_97 = 3'h4 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_4_1 : _GEN_96; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_98 = 3'h4 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_4_2 : _GEN_97; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_99 = 3'h4 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_4_3 : _GEN_98; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_100 = 3'h4 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_4_4 : _GEN_99; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_101 = 3'h4 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_4_5 : _GEN_100; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_102 = 3'h4 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_4_6 : _GEN_101; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_103 = 3'h4 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_4_7 : _GEN_102; // @[ivncontrol4.scala 63:{17,17}]
  wire  _GEN_3903 = 3'h5 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_104 = 3'h5 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_5_0 : _GEN_103; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_105 = 3'h5 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_5_1 : _GEN_104; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_106 = 3'h5 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_5_2 : _GEN_105; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_107 = 3'h5 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_5_3 : _GEN_106; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_108 = 3'h5 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_5_4 : _GEN_107; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_109 = 3'h5 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_5_5 : _GEN_108; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_110 = 3'h5 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_5_6 : _GEN_109; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_111 = 3'h5 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_5_7 : _GEN_110; // @[ivncontrol4.scala 63:{17,17}]
  wire  _GEN_3919 = 3'h6 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_112 = 3'h6 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_6_0 : _GEN_111; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_113 = 3'h6 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_6_1 : _GEN_112; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_114 = 3'h6 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_6_2 : _GEN_113; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_115 = 3'h6 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_6_3 : _GEN_114; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_116 = 3'h6 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_6_4 : _GEN_115; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_117 = 3'h6 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_6_5 : _GEN_116; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_118 = 3'h6 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_6_6 : _GEN_117; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_119 = 3'h6 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_6_7 : _GEN_118; // @[ivncontrol4.scala 63:{17,17}]
  wire  _GEN_3935 = 3'h7 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_120 = 3'h7 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_7_0 : _GEN_119; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_121 = 3'h7 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_7_1 : _GEN_120; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_122 = 3'h7 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_7_2 : _GEN_121; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_123 = 3'h7 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_7_3 : _GEN_122; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_124 = 3'h7 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_7_4 : _GEN_123; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_125 = 3'h7 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_7_5 : _GEN_124; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_126 = 3'h7 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_7_6 : _GEN_125; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_127 = 3'h7 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_7_7 : _GEN_126; // @[ivncontrol4.scala 63:{17,17}]
  wire [31:0] _mat_T_1_T_2 = {{16'd0}, _GEN_127}; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_129 = _GEN_3825 & 4'h1 == j[3:0] ? solution_0_1 : solution_0_0; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_130 = _GEN_3825 & 4'h2 == j[3:0] ? solution_0_2 : _GEN_129; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_131 = _GEN_3825 & 4'h3 == j[3:0] ? solution_0_3 : _GEN_130; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_132 = _GEN_3825 & 4'h4 == j[3:0] ? solution_0_4 : _GEN_131; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_133 = _GEN_3825 & 4'h5 == j[3:0] ? solution_0_5 : _GEN_132; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_134 = _GEN_3825 & 4'h6 == j[3:0] ? solution_0_6 : _GEN_133; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_135 = _GEN_3825 & 4'h7 == j[3:0] ? solution_0_7 : _GEN_134; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_136 = _GEN_3825 & 4'h8 == j[3:0] ? 16'h0 : _GEN_135; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_137 = _GEN_3839 & 4'h0 == j[3:0] ? solution_1_0 : _GEN_136; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_138 = _GEN_3839 & 4'h1 == j[3:0] ? solution_1_1 : _GEN_137; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_139 = _GEN_3839 & 4'h2 == j[3:0] ? solution_1_2 : _GEN_138; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_140 = _GEN_3839 & 4'h3 == j[3:0] ? solution_1_3 : _GEN_139; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_141 = _GEN_3839 & 4'h4 == j[3:0] ? solution_1_4 : _GEN_140; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_142 = _GEN_3839 & 4'h5 == j[3:0] ? solution_1_5 : _GEN_141; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_143 = _GEN_3839 & 4'h6 == j[3:0] ? solution_1_6 : _GEN_142; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_144 = _GEN_3839 & 4'h7 == j[3:0] ? solution_1_7 : _GEN_143; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_145 = _GEN_3839 & 4'h8 == j[3:0] ? 16'h0 : _GEN_144; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_146 = _GEN_3855 & 4'h0 == j[3:0] ? solution_2_0 : _GEN_145; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_147 = _GEN_3855 & 4'h1 == j[3:0] ? solution_2_1 : _GEN_146; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_148 = _GEN_3855 & 4'h2 == j[3:0] ? solution_2_2 : _GEN_147; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_149 = _GEN_3855 & 4'h3 == j[3:0] ? solution_2_3 : _GEN_148; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_150 = _GEN_3855 & 4'h4 == j[3:0] ? solution_2_4 : _GEN_149; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_151 = _GEN_3855 & 4'h5 == j[3:0] ? solution_2_5 : _GEN_150; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_152 = _GEN_3855 & 4'h6 == j[3:0] ? solution_2_6 : _GEN_151; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_153 = _GEN_3855 & 4'h7 == j[3:0] ? solution_2_7 : _GEN_152; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_154 = _GEN_3855 & 4'h8 == j[3:0] ? 16'h0 : _GEN_153; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_155 = _GEN_3871 & 4'h0 == j[3:0] ? solution_3_0 : _GEN_154; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_156 = _GEN_3871 & 4'h1 == j[3:0] ? solution_3_1 : _GEN_155; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_157 = _GEN_3871 & 4'h2 == j[3:0] ? solution_3_2 : _GEN_156; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_158 = _GEN_3871 & 4'h3 == j[3:0] ? solution_3_3 : _GEN_157; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_159 = _GEN_3871 & 4'h4 == j[3:0] ? solution_3_4 : _GEN_158; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_160 = _GEN_3871 & 4'h5 == j[3:0] ? solution_3_5 : _GEN_159; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_161 = _GEN_3871 & 4'h6 == j[3:0] ? solution_3_6 : _GEN_160; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_162 = _GEN_3871 & 4'h7 == j[3:0] ? solution_3_7 : _GEN_161; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_163 = _GEN_3871 & 4'h8 == j[3:0] ? 16'h0 : _GEN_162; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_164 = _GEN_3887 & 4'h0 == j[3:0] ? solution_4_0 : _GEN_163; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_165 = _GEN_3887 & 4'h1 == j[3:0] ? solution_4_1 : _GEN_164; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_166 = _GEN_3887 & 4'h2 == j[3:0] ? solution_4_2 : _GEN_165; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_167 = _GEN_3887 & 4'h3 == j[3:0] ? solution_4_3 : _GEN_166; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_168 = _GEN_3887 & 4'h4 == j[3:0] ? solution_4_4 : _GEN_167; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_169 = _GEN_3887 & 4'h5 == j[3:0] ? solution_4_5 : _GEN_168; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_170 = _GEN_3887 & 4'h6 == j[3:0] ? solution_4_6 : _GEN_169; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_171 = _GEN_3887 & 4'h7 == j[3:0] ? solution_4_7 : _GEN_170; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_172 = _GEN_3887 & 4'h8 == j[3:0] ? 16'h0 : _GEN_171; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_173 = _GEN_3903 & 4'h0 == j[3:0] ? solution_5_0 : _GEN_172; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_174 = _GEN_3903 & 4'h1 == j[3:0] ? solution_5_1 : _GEN_173; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_175 = _GEN_3903 & 4'h2 == j[3:0] ? solution_5_2 : _GEN_174; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_176 = _GEN_3903 & 4'h3 == j[3:0] ? solution_5_3 : _GEN_175; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_177 = _GEN_3903 & 4'h4 == j[3:0] ? solution_5_4 : _GEN_176; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_178 = _GEN_3903 & 4'h5 == j[3:0] ? solution_5_5 : _GEN_177; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_179 = _GEN_3903 & 4'h6 == j[3:0] ? solution_5_6 : _GEN_178; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_180 = _GEN_3903 & 4'h7 == j[3:0] ? solution_5_7 : _GEN_179; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_181 = _GEN_3903 & 4'h8 == j[3:0] ? 16'h0 : _GEN_180; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_182 = _GEN_3919 & 4'h0 == j[3:0] ? solution_6_0 : _GEN_181; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_183 = _GEN_3919 & 4'h1 == j[3:0] ? solution_6_1 : _GEN_182; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_184 = _GEN_3919 & 4'h2 == j[3:0] ? solution_6_2 : _GEN_183; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_185 = _GEN_3919 & 4'h3 == j[3:0] ? solution_6_3 : _GEN_184; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_186 = _GEN_3919 & 4'h4 == j[3:0] ? solution_6_4 : _GEN_185; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_187 = _GEN_3919 & 4'h5 == j[3:0] ? solution_6_5 : _GEN_186; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_188 = _GEN_3919 & 4'h6 == j[3:0] ? solution_6_6 : _GEN_187; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_189 = _GEN_3919 & 4'h7 == j[3:0] ? solution_6_7 : _GEN_188; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_190 = _GEN_3919 & 4'h8 == j[3:0] ? 16'h0 : _GEN_189; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_191 = _GEN_3935 & 4'h0 == j[3:0] ? solution_7_0 : _GEN_190; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_192 = _GEN_3935 & 4'h1 == j[3:0] ? solution_7_1 : _GEN_191; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_193 = _GEN_3935 & 4'h2 == j[3:0] ? solution_7_2 : _GEN_192; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_194 = _GEN_3935 & 4'h3 == j[3:0] ? solution_7_3 : _GEN_193; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_195 = _GEN_3935 & 4'h4 == j[3:0] ? solution_7_4 : _GEN_194; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_196 = _GEN_3935 & 4'h5 == j[3:0] ? solution_7_5 : _GEN_195; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_197 = _GEN_3935 & 4'h6 == j[3:0] ? solution_7_6 : _GEN_196; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_198 = _GEN_3935 & 4'h7 == j[3:0] ? solution_7_7 : _GEN_197; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_199 = _GEN_3935 & 4'h8 == j[3:0] ? 16'h0 : _GEN_198; // @[ivncontrol4.scala 65:{31,31}]
  wire [31:0] _GEN_201 = 3'h1 == i[2:0] ? count_1 : count_0; // @[ivncontrol4.scala 66:{33,33}]
  wire [31:0] _GEN_202 = 3'h2 == i[2:0] ? count_2 : _GEN_201; // @[ivncontrol4.scala 66:{33,33}]
  wire [31:0] _GEN_203 = 3'h3 == i[2:0] ? count_3 : _GEN_202; // @[ivncontrol4.scala 66:{33,33}]
  wire [31:0] _GEN_204 = 3'h4 == i[2:0] ? count_4 : _GEN_203; // @[ivncontrol4.scala 66:{33,33}]
  wire [31:0] _GEN_205 = 3'h5 == i[2:0] ? count_5 : _GEN_204; // @[ivncontrol4.scala 66:{33,33}]
  wire [31:0] _GEN_206 = 3'h6 == i[2:0] ? count_6 : _GEN_205; // @[ivncontrol4.scala 66:{33,33}]
  wire [31:0] _GEN_207 = 3'h7 == i[2:0] ? count_7 : _GEN_206; // @[ivncontrol4.scala 66:{33,33}]
  wire [31:0] _count_T_2 = _GEN_207 + 32'h1; // @[ivncontrol4.scala 66:33]
  wire [31:0] _GEN_208 = 3'h0 == i[2:0] ? _count_T_2 : count_0; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_209 = 3'h1 == i[2:0] ? _count_T_2 : count_1; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_210 = 3'h2 == i[2:0] ? _count_T_2 : count_2; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_211 = 3'h3 == i[2:0] ? _count_T_2 : count_3; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_212 = 3'h4 == i[2:0] ? _count_T_2 : count_4; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_213 = 3'h5 == i[2:0] ? _count_T_2 : count_5; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_214 = 3'h6 == i[2:0] ? _count_T_2 : count_6; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_215 = 3'h7 == i[2:0] ? _count_T_2 : count_7; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_216 = _GEN_199 != 16'h0 ? _GEN_208 : count_0; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_217 = _GEN_199 != 16'h0 ? _GEN_209 : count_1; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_218 = _GEN_199 != 16'h0 ? _GEN_210 : count_2; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_219 = _GEN_199 != 16'h0 ? _GEN_211 : count_3; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_220 = _GEN_199 != 16'h0 ? _GEN_212 : count_4; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_221 = _GEN_199 != 16'h0 ? _GEN_213 : count_5; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_222 = _GEN_199 != 16'h0 ? _GEN_214 : count_6; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_223 = _GEN_199 != 16'h0 ? _GEN_215 : count_7; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_224 = io_validpin ? _GEN_216 : count_0; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _GEN_225 = io_validpin ? _GEN_217 : count_1; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _GEN_226 = io_validpin ? _GEN_218 : count_2; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _GEN_227 = io_validpin ? _GEN_219 : count_3; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _GEN_228 = io_validpin ? _GEN_220 : count_4; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _GEN_229 = io_validpin ? _GEN_221 : count_5; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _GEN_230 = io_validpin ? _GEN_222 : count_6; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _GEN_231 = io_validpin ? _GEN_223 : count_7; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _i_T_1 = i + 32'h1; // @[ivncontrol4.scala 113:16]
  wire [31:0] _GEN_247 = i < 32'h7 & _io_ProcessValid_T_1 ? _i_T_1 : i; // @[ivncontrol4.scala 112:74 113:11 41:20]
  wire [31:0] _j_T_1 = j + 32'h1; // @[ivncontrol4.scala 118:16]
  wire [3:0] _GEN_264 = _io_ProcessValid_T & j == 32'h8 ? 4'h8 : 4'h0; // @[ivncontrol4.scala 120:77 121:11 129:11]
  wire [31:0] _GEN_265 = _io_ProcessValid_T & j == 32'h8 ? 32'h7 : _GEN_247; // @[ivncontrol4.scala 120:77 122:11]
  wire  _GEN_312 = _io_ProcessValid_T_2; // @[ivncontrol4.scala 153:41]
  wire [31:0] _GEN_313 = rowcount_0 != 32'h0 ? 32'h0 : pin; // @[ivncontrol4.scala 162:30 163:13 37:22]
  wire  _T_27 = rowcount_0 == 32'h0; // @[ivncontrol4.scala 165:23]
  wire [31:0] _GEN_314 = rowcount_0 == 32'h0 & rowcount_1 != 32'h0 ? 32'h1 : _GEN_313; // @[ivncontrol4.scala 165:54 166:13]
  wire  _T_32 = _T_27 & rowcount_1 == 32'h0; // @[ivncontrol4.scala 168:31]
  wire [31:0] _GEN_315 = _T_27 & rowcount_1 == 32'h0 & rowcount_2 != 32'h0 ? 32'h2 : _GEN_314; // @[ivncontrol4.scala 168:77 169:13]
  wire  _T_39 = _T_32 & rowcount_2 == 32'h0; // @[ivncontrol4.scala 171:54]
  wire [31:0] _GEN_316 = _T_32 & rowcount_2 == 32'h0 & rowcount_3 != 32'h0 ? 32'h3 : _GEN_315; // @[ivncontrol4.scala 171:100 172:13]
  wire  _T_48 = _T_39 & rowcount_3 == 32'h0; // @[ivncontrol4.scala 174:77]
  wire [31:0] _GEN_317 = _T_39 & rowcount_3 == 32'h0 & rowcount_4 != 32'h0 ? 32'h4 : _GEN_316; // @[ivncontrol4.scala 174:123 175:13]
  wire  _T_59 = _T_48 & rowcount_4 == 32'h0; // @[ivncontrol4.scala 177:100]
  wire  _T_72 = _T_59 & rowcount_5 == 32'h0; // @[ivncontrol4.scala 180:123]
  wire  valid = _io_ProcessValid_T_2; // @[ivncontrol4.scala 153:41]
  wire [32:0] _T_91 = {{1'd0}, pin}; // @[ivncontrol4.scala 191:27]
  wire [31:0] _GEN_322 = 4'h1 == _T_91[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_323 = 4'h2 == _T_91[3:0] ? rowcount_2 : _GEN_322; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_324 = 4'h3 == _T_91[3:0] ? rowcount_3 : _GEN_323; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_325 = 4'h4 == _T_91[3:0] ? rowcount_4 : _GEN_324; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_326 = 4'h5 == _T_91[3:0] ? rowcount_5 : _GEN_325; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_327 = 4'h6 == _T_91[3:0] ? rowcount_6 : _GEN_326; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_328 = 4'h7 == _T_91[3:0] ? rowcount_7 : _GEN_327; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_329 = 4'h8 == _T_91[3:0] ? rowcount_8 : _GEN_328; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_330 = 4'h9 == _T_91[3:0] ? rowcount_9 : _GEN_329; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_331 = 4'ha == _T_91[3:0] ? rowcount_10 : _GEN_330; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_332 = 4'hb == _T_91[3:0] ? rowcount_11 : _GEN_331; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_333 = 4'hc == _T_91[3:0] ? rowcount_12 : _GEN_332; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_334 = 4'hd == _T_91[3:0] ? rowcount_13 : _GEN_333; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_335 = 4'he == _T_91[3:0] ? rowcount_14 : _GEN_334; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_336 = 4'hf == _T_91[3:0] ? rowcount_15 : _GEN_335; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_449 = _GEN_336 == 32'h1 ? _T_91[31:0] : 32'hc; // @[ivncontrol4.scala 142:17 241:50 242:21]
  wire [31:0] _GEN_450 = _GEN_336 == 32'h2 ? _T_91[31:0] : _GEN_449; // @[ivncontrol4.scala 237:51 238:21]
  wire [31:0] _GEN_451 = _GEN_336 == 32'h2 ? _T_91[31:0] : 32'h1; // @[ivncontrol4.scala 142:17 237:51 239:21]
  wire [31:0] _GEN_452 = _GEN_336 == 32'h3 ? _T_91[31:0] : _GEN_450; // @[ivncontrol4.scala 232:50 233:21]
  wire [31:0] _GEN_453 = _GEN_336 == 32'h3 ? _T_91[31:0] : _GEN_451; // @[ivncontrol4.scala 232:50 234:21]
  wire [31:0] _GEN_454 = _GEN_336 == 32'h3 ? _T_91[31:0] : 32'h1a; // @[ivncontrol4.scala 142:17 232:50 235:21]
  wire [31:0] _GEN_455 = _GEN_336 == 32'h4 ? _T_91[31:0] : _GEN_452; // @[ivncontrol4.scala 224:50 225:21]
  wire [31:0] _GEN_456 = _GEN_336 == 32'h4 ? _T_91[31:0] : _GEN_453; // @[ivncontrol4.scala 224:50 226:21]
  wire [31:0] _GEN_457 = _GEN_336 == 32'h4 ? _T_91[31:0] : _GEN_454; // @[ivncontrol4.scala 224:50 227:21]
  wire [31:0] _GEN_458 = _GEN_336 == 32'h4 ? _T_91[31:0] : 32'h1b; // @[ivncontrol4.scala 142:17 224:50 228:21]
  wire [31:0] _GEN_459 = _GEN_336 == 32'h5 ? _T_91[31:0] : _GEN_455; // @[ivncontrol4.scala 217:50 218:21]
  wire [31:0] _GEN_460 = _GEN_336 == 32'h5 ? _T_91[31:0] : _GEN_456; // @[ivncontrol4.scala 217:50 219:21]
  wire [31:0] _GEN_461 = _GEN_336 == 32'h5 ? _T_91[31:0] : _GEN_457; // @[ivncontrol4.scala 217:50 220:21]
  wire [31:0] _GEN_462 = _GEN_336 == 32'h5 ? _T_91[31:0] : _GEN_458; // @[ivncontrol4.scala 217:50 221:21]
  wire [31:0] _GEN_463 = _GEN_336 == 32'h5 ? _T_91[31:0] : 32'h13; // @[ivncontrol4.scala 143:18 217:50 222:22]
  wire [31:0] _GEN_464 = _GEN_336 == 32'h6 ? _T_91[31:0] : _GEN_459; // @[ivncontrol4.scala 209:52 210:21]
  wire [31:0] _GEN_465 = _GEN_336 == 32'h6 ? _T_91[31:0] : _GEN_460; // @[ivncontrol4.scala 209:52 211:21]
  wire [31:0] _GEN_466 = _GEN_336 == 32'h6 ? _T_91[31:0] : _GEN_461; // @[ivncontrol4.scala 209:52 212:21]
  wire [31:0] _GEN_467 = _GEN_336 == 32'h6 ? _T_91[31:0] : _GEN_462; // @[ivncontrol4.scala 209:52 213:21]
  wire [31:0] _GEN_468 = _GEN_336 == 32'h6 ? _T_91[31:0] : _GEN_463; // @[ivncontrol4.scala 209:52 214:22]
  wire [31:0] _GEN_469 = _GEN_336 == 32'h6 ? _T_91[31:0] : 32'ha; // @[ivncontrol4.scala 143:18 209:52 215:22]
  wire [31:0] _GEN_470 = _GEN_336 == 32'h7 ? _T_91[31:0] : _GEN_464; // @[ivncontrol4.scala 201:52 202:21]
  wire [31:0] _GEN_471 = _GEN_336 == 32'h7 ? _T_91[31:0] : _GEN_465; // @[ivncontrol4.scala 201:52 203:21]
  wire [31:0] _GEN_472 = _GEN_336 == 32'h7 ? _T_91[31:0] : _GEN_466; // @[ivncontrol4.scala 201:52 204:21]
  wire [31:0] _GEN_473 = _GEN_336 == 32'h7 ? _T_91[31:0] : _GEN_467; // @[ivncontrol4.scala 201:52 205:21]
  wire [31:0] _GEN_474 = _GEN_336 == 32'h7 ? _T_91[31:0] : _GEN_468; // @[ivncontrol4.scala 201:52 206:22]
  wire [31:0] _GEN_475 = _GEN_336 == 32'h7 ? _T_91[31:0] : _GEN_469; // @[ivncontrol4.scala 201:52 207:22]
  wire [31:0] _GEN_476 = _GEN_336 == 32'h7 ? _T_91[31:0] : 32'h6; // @[ivncontrol4.scala 143:18 201:52 208:22]
  wire [31:0] _GEN_477 = _GEN_336 >= 32'h8 ? _T_91[31:0] : _GEN_470; // @[ivncontrol4.scala 191:42 192:21]
  wire [31:0] _GEN_478 = _GEN_336 >= 32'h8 ? _T_91[31:0] : _GEN_471; // @[ivncontrol4.scala 191:42 193:21]
  wire [31:0] _GEN_479 = _GEN_336 >= 32'h8 ? _T_91[31:0] : _GEN_472; // @[ivncontrol4.scala 191:42 194:21]
  wire [31:0] _GEN_480 = _GEN_336 >= 32'h8 ? _T_91[31:0] : _GEN_473; // @[ivncontrol4.scala 191:42 195:21]
  wire [31:0] _GEN_481 = _GEN_336 >= 32'h8 ? _T_91[31:0] : _GEN_474; // @[ivncontrol4.scala 191:42 196:22]
  wire [31:0] _GEN_482 = _GEN_336 >= 32'h8 ? _T_91[31:0] : _GEN_475; // @[ivncontrol4.scala 191:42 197:22]
  wire [31:0] _GEN_483 = _GEN_336 >= 32'h8 ? _T_91[31:0] : _GEN_476; // @[ivncontrol4.scala 191:42 198:22]
  wire [31:0] _GEN_484 = _GEN_336 >= 32'h8 ? _T_91[31:0] : 32'h1b; // @[ivncontrol4.scala 143:18 191:42 199:22]
  wire [31:0] _T_127 = 32'h8 - _GEN_336; // @[ivncontrol4.scala 245:18]
  wire [31:0] _i_vn_1_T_15 = 32'h1 + pin; // @[ivncontrol4.scala 246:29]
  wire [31:0] _GEN_597 = _T_127 == 32'h1 ? _i_vn_1_T_15 : _GEN_484; // @[ivncontrol4.scala 286:54 289:22]
  wire [31:0] _GEN_598 = _T_127 == 32'h2 ? _i_vn_1_T_15 : _GEN_483; // @[ivncontrol4.scala 281:54 284:22]
  wire [31:0] _GEN_599 = _T_127 == 32'h2 ? _i_vn_1_T_15 : _GEN_597; // @[ivncontrol4.scala 281:54 285:22]
  wire [31:0] _GEN_600 = _T_127 == 32'h3 ? _i_vn_1_T_15 : _GEN_482; // @[ivncontrol4.scala 274:54 276:22]
  wire [31:0] _GEN_601 = _T_127 == 32'h3 ? _i_vn_1_T_15 : _GEN_598; // @[ivncontrol4.scala 274:54 277:22]
  wire [31:0] _GEN_602 = _T_127 == 32'h3 ? _i_vn_1_T_15 : _GEN_599; // @[ivncontrol4.scala 274:54 278:22]
  wire [31:0] _GEN_603 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_481; // @[ivncontrol4.scala 268:54 270:22]
  wire [31:0] _GEN_604 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_600; // @[ivncontrol4.scala 268:54 271:22]
  wire [31:0] _GEN_605 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_601; // @[ivncontrol4.scala 268:54 272:22]
  wire [31:0] _GEN_606 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_602; // @[ivncontrol4.scala 268:54 273:22]
  wire [31:0] _GEN_607 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_480; // @[ivncontrol4.scala 261:54 263:21]
  wire [31:0] _GEN_608 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_603; // @[ivncontrol4.scala 261:54 264:22]
  wire [31:0] _GEN_609 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_604; // @[ivncontrol4.scala 261:54 265:22]
  wire [31:0] _GEN_610 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_605; // @[ivncontrol4.scala 261:54 266:22]
  wire [31:0] _GEN_611 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_606; // @[ivncontrol4.scala 261:54 267:22]
  wire [31:0] _GEN_612 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_479; // @[ivncontrol4.scala 254:54 255:22]
  wire [31:0] _GEN_613 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_607; // @[ivncontrol4.scala 254:54 256:21]
  wire [31:0] _GEN_614 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_608; // @[ivncontrol4.scala 254:54 257:22]
  wire [31:0] _GEN_615 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_609; // @[ivncontrol4.scala 254:54 258:22]
  wire [31:0] _GEN_616 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_610; // @[ivncontrol4.scala 254:54 259:22]
  wire [31:0] _GEN_617 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_611; // @[ivncontrol4.scala 254:54 260:22]
  wire [31:0] _GEN_618 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_478; // @[ivncontrol4.scala 245:49 246:22]
  wire [31:0] _GEN_619 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_612; // @[ivncontrol4.scala 245:49 247:21]
  wire [31:0] _GEN_620 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_613; // @[ivncontrol4.scala 245:49 248:21]
  wire [31:0] _GEN_621 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_614; // @[ivncontrol4.scala 245:49 249:22]
  wire [31:0] _GEN_622 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_615; // @[ivncontrol4.scala 245:49 250:22]
  wire [31:0] _GEN_623 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_616; // @[ivncontrol4.scala 245:49 251:22]
  wire [31:0] _GEN_624 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_617; // @[ivncontrol4.scala 245:49 252:22]
  wire [31:0] _GEN_642 = 4'h1 == _i_vn_1_T_15[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_643 = 4'h2 == _i_vn_1_T_15[3:0] ? rowcount_2 : _GEN_642; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_644 = 4'h3 == _i_vn_1_T_15[3:0] ? rowcount_3 : _GEN_643; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_645 = 4'h4 == _i_vn_1_T_15[3:0] ? rowcount_4 : _GEN_644; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_646 = 4'h5 == _i_vn_1_T_15[3:0] ? rowcount_5 : _GEN_645; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_647 = 4'h6 == _i_vn_1_T_15[3:0] ? rowcount_6 : _GEN_646; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_648 = 4'h7 == _i_vn_1_T_15[3:0] ? rowcount_7 : _GEN_647; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_649 = 4'h8 == _i_vn_1_T_15[3:0] ? rowcount_8 : _GEN_648; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_650 = 4'h9 == _i_vn_1_T_15[3:0] ? rowcount_9 : _GEN_649; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_651 = 4'ha == _i_vn_1_T_15[3:0] ? rowcount_10 : _GEN_650; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_652 = 4'hb == _i_vn_1_T_15[3:0] ? rowcount_11 : _GEN_651; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_653 = 4'hc == _i_vn_1_T_15[3:0] ? rowcount_12 : _GEN_652; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_654 = 4'hd == _i_vn_1_T_15[3:0] ? rowcount_13 : _GEN_653; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_655 = 4'he == _i_vn_1_T_15[3:0] ? rowcount_14 : _GEN_654; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_656 = 4'hf == _i_vn_1_T_15[3:0] ? rowcount_15 : _GEN_655; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _T_172 = _GEN_336 + _GEN_656; // @[ivncontrol4.scala 292:41]
  wire [31:0] _T_174 = 32'h8 - _T_172; // @[ivncontrol4.scala 292:18]
  wire [31:0] _i_vn_1_T_17 = 32'h2 + pin; // @[ivncontrol4.scala 293:29]
  wire [31:0] _GEN_849 = _T_174 == 32'h1 ? _i_vn_1_T_17 : _GEN_624; // @[ivncontrol4.scala 335:78 338:22]
  wire [31:0] _GEN_850 = _T_174 == 32'h2 ? _i_vn_1_T_17 : _GEN_623; // @[ivncontrol4.scala 329:76 332:22]
  wire [31:0] _GEN_851 = _T_174 == 32'h2 ? _i_vn_1_T_17 : _GEN_849; // @[ivncontrol4.scala 329:76 333:22]
  wire [31:0] _GEN_852 = _T_174 == 32'h3 ? _i_vn_1_T_17 : _GEN_622; // @[ivncontrol4.scala 322:78 324:23]
  wire [31:0] _GEN_853 = _T_174 == 32'h3 ? _i_vn_1_T_17 : _GEN_850; // @[ivncontrol4.scala 322:78 325:22]
  wire [31:0] _GEN_854 = _T_174 == 32'h3 ? _i_vn_1_T_17 : _GEN_851; // @[ivncontrol4.scala 322:78 326:22]
  wire [31:0] _GEN_855 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_621; // @[ivncontrol4.scala 316:78 318:22]
  wire [31:0] _GEN_856 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_852; // @[ivncontrol4.scala 316:78 319:22]
  wire [31:0] _GEN_857 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_853; // @[ivncontrol4.scala 316:78 320:22]
  wire [31:0] _GEN_858 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_854; // @[ivncontrol4.scala 316:78 321:22]
  wire [31:0] _GEN_859 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_620; // @[ivncontrol4.scala 309:76 311:23]
  wire [31:0] _GEN_860 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_855; // @[ivncontrol4.scala 309:76 312:22]
  wire [31:0] _GEN_861 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_856; // @[ivncontrol4.scala 309:76 313:22]
  wire [31:0] _GEN_862 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_857; // @[ivncontrol4.scala 309:76 314:22]
  wire [31:0] _GEN_863 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_858; // @[ivncontrol4.scala 309:76 315:22]
  wire [31:0] _GEN_864 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_619; // @[ivncontrol4.scala 301:77 303:22]
  wire [31:0] _GEN_865 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_859; // @[ivncontrol4.scala 301:77 304:21]
  wire [31:0] _GEN_866 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_860; // @[ivncontrol4.scala 301:77 305:22]
  wire [31:0] _GEN_867 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_861; // @[ivncontrol4.scala 301:77 306:22]
  wire [31:0] _GEN_868 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_862; // @[ivncontrol4.scala 301:77 307:22]
  wire [31:0] _GEN_869 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_863; // @[ivncontrol4.scala 301:77 308:22]
  wire [31:0] _GEN_870 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_618; // @[ivncontrol4.scala 292:73 293:22]
  wire [31:0] _GEN_871 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_864; // @[ivncontrol4.scala 292:73 294:21]
  wire [31:0] _GEN_872 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_865; // @[ivncontrol4.scala 292:73 295:21]
  wire [31:0] _GEN_873 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_866; // @[ivncontrol4.scala 292:73 296:22]
  wire [31:0] _GEN_874 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_867; // @[ivncontrol4.scala 292:73 297:22]
  wire [31:0] _GEN_875 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_868; // @[ivncontrol4.scala 292:73 298:22]
  wire [31:0] _GEN_876 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_869; // @[ivncontrol4.scala 292:73 299:22]
  wire [31:0] _GEN_910 = 4'h1 == _i_vn_1_T_17[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_911 = 4'h2 == _i_vn_1_T_17[3:0] ? rowcount_2 : _GEN_910; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_912 = 4'h3 == _i_vn_1_T_17[3:0] ? rowcount_3 : _GEN_911; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_913 = 4'h4 == _i_vn_1_T_17[3:0] ? rowcount_4 : _GEN_912; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_914 = 4'h5 == _i_vn_1_T_17[3:0] ? rowcount_5 : _GEN_913; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_915 = 4'h6 == _i_vn_1_T_17[3:0] ? rowcount_6 : _GEN_914; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_916 = 4'h7 == _i_vn_1_T_17[3:0] ? rowcount_7 : _GEN_915; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_917 = 4'h8 == _i_vn_1_T_17[3:0] ? rowcount_8 : _GEN_916; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_918 = 4'h9 == _i_vn_1_T_17[3:0] ? rowcount_9 : _GEN_917; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_919 = 4'ha == _i_vn_1_T_17[3:0] ? rowcount_10 : _GEN_918; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_920 = 4'hb == _i_vn_1_T_17[3:0] ? rowcount_11 : _GEN_919; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_921 = 4'hc == _i_vn_1_T_17[3:0] ? rowcount_12 : _GEN_920; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_922 = 4'hd == _i_vn_1_T_17[3:0] ? rowcount_13 : _GEN_921; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_923 = 4'he == _i_vn_1_T_17[3:0] ? rowcount_14 : _GEN_922; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_924 = 4'hf == _i_vn_1_T_17[3:0] ? rowcount_15 : _GEN_923; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _T_254 = _T_172 + _GEN_924; // @[ivncontrol4.scala 343:62]
  wire [31:0] _T_256 = 32'h8 - _T_254; // @[ivncontrol4.scala 343:17]
  wire [31:0] _i_vn_1_T_19 = 32'h3 + pin; // @[ivncontrol4.scala 344:29]
  wire [31:0] _GEN_1213 = _T_256 == 32'h1 ? _i_vn_1_T_19 : _GEN_876; // @[ivncontrol4.scala 386:100 389:22]
  wire [31:0] _GEN_1214 = _T_256 == 32'h2 ? _i_vn_1_T_19 : _GEN_875; // @[ivncontrol4.scala 380:98 383:22]
  wire [31:0] _GEN_1215 = _T_256 == 32'h2 ? _i_vn_1_T_19 : _GEN_1213; // @[ivncontrol4.scala 380:98 384:22]
  wire [31:0] _GEN_1216 = _T_256 == 32'h3 ? _i_vn_1_T_19 : _GEN_874; // @[ivncontrol4.scala 373:100 375:23]
  wire [31:0] _GEN_1217 = _T_256 == 32'h3 ? _i_vn_1_T_19 : _GEN_1214; // @[ivncontrol4.scala 373:100 376:22]
  wire [31:0] _GEN_1218 = _T_256 == 32'h3 ? _i_vn_1_T_19 : _GEN_1215; // @[ivncontrol4.scala 373:100 377:22]
  wire [31:0] _GEN_1219 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_873; // @[ivncontrol4.scala 367:100 369:22]
  wire [31:0] _GEN_1220 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_1216; // @[ivncontrol4.scala 367:100 370:22]
  wire [31:0] _GEN_1221 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_1217; // @[ivncontrol4.scala 367:100 371:22]
  wire [31:0] _GEN_1222 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_1218; // @[ivncontrol4.scala 367:100 372:22]
  wire [31:0] _GEN_1223 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_872; // @[ivncontrol4.scala 360:98 362:23]
  wire [31:0] _GEN_1224 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1219; // @[ivncontrol4.scala 360:98 363:22]
  wire [31:0] _GEN_1225 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1220; // @[ivncontrol4.scala 360:98 364:22]
  wire [31:0] _GEN_1226 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1221; // @[ivncontrol4.scala 360:98 365:22]
  wire [31:0] _GEN_1227 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1222; // @[ivncontrol4.scala 360:98 366:22]
  wire [31:0] _GEN_1228 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_871; // @[ivncontrol4.scala 352:99 354:22]
  wire [31:0] _GEN_1229 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1223; // @[ivncontrol4.scala 352:99 355:21]
  wire [31:0] _GEN_1230 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1224; // @[ivncontrol4.scala 352:99 356:22]
  wire [31:0] _GEN_1231 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1225; // @[ivncontrol4.scala 352:99 357:22]
  wire [31:0] _GEN_1232 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1226; // @[ivncontrol4.scala 352:99 358:22]
  wire [31:0] _GEN_1233 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1227; // @[ivncontrol4.scala 352:99 359:22]
  wire [31:0] _GEN_1234 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_870; // @[ivncontrol4.scala 343:94 344:22]
  wire [31:0] _GEN_1235 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1228; // @[ivncontrol4.scala 343:94 345:21]
  wire [31:0] _GEN_1236 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1229; // @[ivncontrol4.scala 343:94 346:21]
  wire [31:0] _GEN_1237 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1230; // @[ivncontrol4.scala 343:94 347:22]
  wire [31:0] _GEN_1238 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1231; // @[ivncontrol4.scala 343:94 348:22]
  wire [31:0] _GEN_1239 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1232; // @[ivncontrol4.scala 343:94 349:22]
  wire [31:0] _GEN_1240 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1233; // @[ivncontrol4.scala 343:94 350:22]
  wire [31:0] _GEN_1290 = 4'h1 == _i_vn_1_T_19[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1291 = 4'h2 == _i_vn_1_T_19[3:0] ? rowcount_2 : _GEN_1290; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1292 = 4'h3 == _i_vn_1_T_19[3:0] ? rowcount_3 : _GEN_1291; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1293 = 4'h4 == _i_vn_1_T_19[3:0] ? rowcount_4 : _GEN_1292; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1294 = 4'h5 == _i_vn_1_T_19[3:0] ? rowcount_5 : _GEN_1293; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1295 = 4'h6 == _i_vn_1_T_19[3:0] ? rowcount_6 : _GEN_1294; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1296 = 4'h7 == _i_vn_1_T_19[3:0] ? rowcount_7 : _GEN_1295; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1297 = 4'h8 == _i_vn_1_T_19[3:0] ? rowcount_8 : _GEN_1296; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1298 = 4'h9 == _i_vn_1_T_19[3:0] ? rowcount_9 : _GEN_1297; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1299 = 4'ha == _i_vn_1_T_19[3:0] ? rowcount_10 : _GEN_1298; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1300 = 4'hb == _i_vn_1_T_19[3:0] ? rowcount_11 : _GEN_1299; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1301 = 4'hc == _i_vn_1_T_19[3:0] ? rowcount_12 : _GEN_1300; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1302 = 4'hd == _i_vn_1_T_19[3:0] ? rowcount_13 : _GEN_1301; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1303 = 4'he == _i_vn_1_T_19[3:0] ? rowcount_14 : _GEN_1302; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1304 = 4'hf == _i_vn_1_T_19[3:0] ? rowcount_15 : _GEN_1303; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _T_371 = _T_254 + _GEN_1304; // @[ivncontrol4.scala 393:86]
  wire [31:0] _T_373 = 32'h8 - _T_371; // @[ivncontrol4.scala 393:19]
  wire [31:0] _i_vn_1_T_21 = 32'h4 + pin; // @[ivncontrol4.scala 394:29]
  wire [31:0] _GEN_1689 = _T_373 == 32'h1 ? _i_vn_1_T_21 : _GEN_1240; // @[ivncontrol4.scala 436:122 439:22]
  wire [31:0] _GEN_1690 = _T_373 == 32'h2 ? _i_vn_1_T_21 : _GEN_1239; // @[ivncontrol4.scala 430:121 433:22]
  wire [31:0] _GEN_1691 = _T_373 == 32'h2 ? _i_vn_1_T_21 : _GEN_1689; // @[ivncontrol4.scala 430:121 434:22]
  wire [31:0] _GEN_1692 = _T_373 == 32'h3 ? _i_vn_1_T_21 : _GEN_1238; // @[ivncontrol4.scala 423:123 425:23]
  wire [31:0] _GEN_1693 = _T_373 == 32'h3 ? _i_vn_1_T_21 : _GEN_1690; // @[ivncontrol4.scala 423:123 426:22]
  wire [31:0] _GEN_1694 = _T_373 == 32'h3 ? _i_vn_1_T_21 : _GEN_1691; // @[ivncontrol4.scala 423:123 427:22]
  wire [31:0] _GEN_1695 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1237; // @[ivncontrol4.scala 417:122 419:22]
  wire [31:0] _GEN_1696 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1692; // @[ivncontrol4.scala 417:122 420:22]
  wire [31:0] _GEN_1697 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1693; // @[ivncontrol4.scala 417:122 421:22]
  wire [31:0] _GEN_1698 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1694; // @[ivncontrol4.scala 417:122 422:22]
  wire [31:0] _GEN_1699 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1236; // @[ivncontrol4.scala 410:121 412:23]
  wire [31:0] _GEN_1700 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1695; // @[ivncontrol4.scala 410:121 413:22]
  wire [31:0] _GEN_1701 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1696; // @[ivncontrol4.scala 410:121 414:22]
  wire [31:0] _GEN_1702 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1697; // @[ivncontrol4.scala 410:121 415:22]
  wire [31:0] _GEN_1703 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1698; // @[ivncontrol4.scala 410:121 416:22]
  wire [31:0] _GEN_1704 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1235; // @[ivncontrol4.scala 402:121 404:22]
  wire [31:0] _GEN_1705 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1699; // @[ivncontrol4.scala 402:121 405:21]
  wire [31:0] _GEN_1706 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1700; // @[ivncontrol4.scala 402:121 406:22]
  wire [31:0] _GEN_1707 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1701; // @[ivncontrol4.scala 402:121 407:22]
  wire [31:0] _GEN_1708 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1702; // @[ivncontrol4.scala 402:121 408:22]
  wire [31:0] _GEN_1709 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1703; // @[ivncontrol4.scala 402:121 409:22]
  wire [31:0] _GEN_1710 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1234; // @[ivncontrol4.scala 393:118 394:22]
  wire [31:0] _GEN_1711 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1704; // @[ivncontrol4.scala 393:118 395:21]
  wire [31:0] _GEN_1712 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1705; // @[ivncontrol4.scala 393:118 396:21]
  wire [31:0] _GEN_1713 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1706; // @[ivncontrol4.scala 393:118 397:22]
  wire [31:0] _GEN_1714 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1707; // @[ivncontrol4.scala 393:118 398:22]
  wire [31:0] _GEN_1715 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1708; // @[ivncontrol4.scala 393:118 399:22]
  wire [31:0] _GEN_1716 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1709; // @[ivncontrol4.scala 393:118 400:22]
  wire [31:0] _GEN_1782 = 4'h1 == _i_vn_1_T_21[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1783 = 4'h2 == _i_vn_1_T_21[3:0] ? rowcount_2 : _GEN_1782; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1784 = 4'h3 == _i_vn_1_T_21[3:0] ? rowcount_3 : _GEN_1783; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1785 = 4'h4 == _i_vn_1_T_21[3:0] ? rowcount_4 : _GEN_1784; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1786 = 4'h5 == _i_vn_1_T_21[3:0] ? rowcount_5 : _GEN_1785; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1787 = 4'h6 == _i_vn_1_T_21[3:0] ? rowcount_6 : _GEN_1786; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1788 = 4'h7 == _i_vn_1_T_21[3:0] ? rowcount_7 : _GEN_1787; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1789 = 4'h8 == _i_vn_1_T_21[3:0] ? rowcount_8 : _GEN_1788; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1790 = 4'h9 == _i_vn_1_T_21[3:0] ? rowcount_9 : _GEN_1789; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1791 = 4'ha == _i_vn_1_T_21[3:0] ? rowcount_10 : _GEN_1790; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1792 = 4'hb == _i_vn_1_T_21[3:0] ? rowcount_11 : _GEN_1791; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1793 = 4'hc == _i_vn_1_T_21[3:0] ? rowcount_12 : _GEN_1792; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1794 = 4'hd == _i_vn_1_T_21[3:0] ? rowcount_13 : _GEN_1793; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1795 = 4'he == _i_vn_1_T_21[3:0] ? rowcount_14 : _GEN_1794; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1796 = 4'hf == _i_vn_1_T_21[3:0] ? rowcount_15 : _GEN_1795; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _T_523 = _T_371 + _GEN_1796; // @[ivncontrol4.scala 443:108]
  wire [31:0] _T_525 = 32'h8 - _T_523; // @[ivncontrol4.scala 443:19]
  wire [31:0] _i_vn_1_T_23 = 32'h5 + pin; // @[ivncontrol4.scala 444:29]
  wire [31:0] _GEN_2277 = _T_525 == 32'h1 ? _i_vn_1_T_23 : _GEN_1716; // @[ivncontrol4.scala 486:144 489:22]
  wire [31:0] _GEN_2278 = _T_525 == 32'h2 ? _i_vn_1_T_23 : _GEN_1715; // @[ivncontrol4.scala 480:143 483:22]
  wire [31:0] _GEN_2279 = _T_525 == 32'h2 ? _i_vn_1_T_23 : _GEN_2277; // @[ivncontrol4.scala 480:143 484:22]
  wire [31:0] _GEN_2280 = _T_525 == 32'h3 ? _i_vn_1_T_23 : _GEN_1714; // @[ivncontrol4.scala 473:145 475:23]
  wire [31:0] _GEN_2281 = _T_525 == 32'h3 ? _i_vn_1_T_23 : _GEN_2278; // @[ivncontrol4.scala 473:145 476:22]
  wire [31:0] _GEN_2282 = _T_525 == 32'h3 ? _i_vn_1_T_23 : _GEN_2279; // @[ivncontrol4.scala 473:145 477:22]
  wire [31:0] _GEN_2283 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_1713; // @[ivncontrol4.scala 467:143 469:22]
  wire [31:0] _GEN_2284 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_2280; // @[ivncontrol4.scala 467:143 470:22]
  wire [31:0] _GEN_2285 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_2281; // @[ivncontrol4.scala 467:143 471:22]
  wire [31:0] _GEN_2286 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_2282; // @[ivncontrol4.scala 467:143 472:22]
  wire [31:0] _GEN_2287 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_1712; // @[ivncontrol4.scala 460:143 462:23]
  wire [31:0] _GEN_2288 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2283; // @[ivncontrol4.scala 460:143 463:22]
  wire [31:0] _GEN_2289 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2284; // @[ivncontrol4.scala 460:143 464:22]
  wire [31:0] _GEN_2290 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2285; // @[ivncontrol4.scala 460:143 465:22]
  wire [31:0] _GEN_2291 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2286; // @[ivncontrol4.scala 460:143 466:22]
  wire [31:0] _GEN_2292 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_1711; // @[ivncontrol4.scala 452:143 454:22]
  wire [31:0] _GEN_2293 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2287; // @[ivncontrol4.scala 452:143 455:21]
  wire [31:0] _GEN_2294 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2288; // @[ivncontrol4.scala 452:143 456:22]
  wire [31:0] _GEN_2295 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2289; // @[ivncontrol4.scala 452:143 457:22]
  wire [31:0] _GEN_2296 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2290; // @[ivncontrol4.scala 452:143 458:22]
  wire [31:0] _GEN_2297 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2291; // @[ivncontrol4.scala 452:143 459:22]
  wire [31:0] _GEN_2298 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_1710; // @[ivncontrol4.scala 443:140 444:22]
  wire [31:0] _GEN_2299 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2292; // @[ivncontrol4.scala 443:140 445:21]
  wire [31:0] _GEN_2300 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2293; // @[ivncontrol4.scala 443:140 446:21]
  wire [31:0] _GEN_2301 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2294; // @[ivncontrol4.scala 443:140 447:22]
  wire [31:0] _GEN_2302 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2295; // @[ivncontrol4.scala 443:140 448:22]
  wire [31:0] _GEN_2303 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2296; // @[ivncontrol4.scala 443:140 449:22]
  wire [31:0] _GEN_2304 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2297; // @[ivncontrol4.scala 443:140 450:22]
  wire [31:0] _GEN_2386 = 4'h1 == _i_vn_1_T_23[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2387 = 4'h2 == _i_vn_1_T_23[3:0] ? rowcount_2 : _GEN_2386; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2388 = 4'h3 == _i_vn_1_T_23[3:0] ? rowcount_3 : _GEN_2387; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2389 = 4'h4 == _i_vn_1_T_23[3:0] ? rowcount_4 : _GEN_2388; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2390 = 4'h5 == _i_vn_1_T_23[3:0] ? rowcount_5 : _GEN_2389; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2391 = 4'h6 == _i_vn_1_T_23[3:0] ? rowcount_6 : _GEN_2390; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2392 = 4'h7 == _i_vn_1_T_23[3:0] ? rowcount_7 : _GEN_2391; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2393 = 4'h8 == _i_vn_1_T_23[3:0] ? rowcount_8 : _GEN_2392; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2394 = 4'h9 == _i_vn_1_T_23[3:0] ? rowcount_9 : _GEN_2393; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2395 = 4'ha == _i_vn_1_T_23[3:0] ? rowcount_10 : _GEN_2394; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2396 = 4'hb == _i_vn_1_T_23[3:0] ? rowcount_11 : _GEN_2395; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2397 = 4'hc == _i_vn_1_T_23[3:0] ? rowcount_12 : _GEN_2396; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2398 = 4'hd == _i_vn_1_T_23[3:0] ? rowcount_13 : _GEN_2397; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2399 = 4'he == _i_vn_1_T_23[3:0] ? rowcount_14 : _GEN_2398; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2400 = 4'hf == _i_vn_1_T_23[3:0] ? rowcount_15 : _GEN_2399; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _T_710 = _T_523 + _GEN_2400; // @[ivncontrol4.scala 494:130]
  wire [31:0] _T_712 = 32'h8 - _T_710; // @[ivncontrol4.scala 494:19]
  wire [31:0] _i_vn_1_T_25 = 32'h6 + pin; // @[ivncontrol4.scala 495:29]
  wire [31:0] _GEN_2977 = _T_712 == 32'h1 ? _i_vn_1_T_25 : _GEN_2304; // @[ivncontrol4.scala 537:166 540:22]
  wire [31:0] _GEN_2978 = _T_712 == 32'h2 ? _i_vn_1_T_25 : _GEN_2303; // @[ivncontrol4.scala 531:166 534:22]
  wire [31:0] _GEN_2979 = _T_712 == 32'h2 ? _i_vn_1_T_25 : _GEN_2977; // @[ivncontrol4.scala 531:166 535:22]
  wire [31:0] _GEN_2980 = _T_712 == 32'h3 ? _i_vn_1_T_25 : _GEN_2302; // @[ivncontrol4.scala 524:168 526:23]
  wire [31:0] _GEN_2981 = _T_712 == 32'h3 ? _i_vn_1_T_25 : _GEN_2978; // @[ivncontrol4.scala 524:168 527:22]
  wire [31:0] _GEN_2982 = _T_712 == 32'h3 ? _i_vn_1_T_25 : _GEN_2979; // @[ivncontrol4.scala 524:168 528:22]
  wire [31:0] _GEN_2983 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2301; // @[ivncontrol4.scala 518:166 520:22]
  wire [31:0] _GEN_2984 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2980; // @[ivncontrol4.scala 518:166 521:22]
  wire [31:0] _GEN_2985 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2981; // @[ivncontrol4.scala 518:166 522:22]
  wire [31:0] _GEN_2986 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2982; // @[ivncontrol4.scala 518:166 523:22]
  wire [31:0] _GEN_2987 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2300; // @[ivncontrol4.scala 511:166 513:23]
  wire [31:0] _GEN_2988 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2983; // @[ivncontrol4.scala 511:166 514:22]
  wire [31:0] _GEN_2989 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2984; // @[ivncontrol4.scala 511:166 515:22]
  wire [31:0] _GEN_2990 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2985; // @[ivncontrol4.scala 511:166 516:22]
  wire [31:0] _GEN_2991 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2986; // @[ivncontrol4.scala 511:166 517:22]
  wire [31:0] _GEN_2992 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2299; // @[ivncontrol4.scala 503:166 505:22]
  wire [31:0] _GEN_2993 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2987; // @[ivncontrol4.scala 503:166 506:21]
  wire [31:0] _GEN_2994 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2988; // @[ivncontrol4.scala 503:166 507:22]
  wire [31:0] _GEN_2995 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2989; // @[ivncontrol4.scala 503:166 508:22]
  wire [31:0] _GEN_2996 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2990; // @[ivncontrol4.scala 503:166 509:22]
  wire [31:0] _GEN_2997 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2991; // @[ivncontrol4.scala 503:166 510:22]
  wire [31:0] _GEN_2998 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2298; // @[ivncontrol4.scala 494:162 495:22]
  wire [31:0] _GEN_2999 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2992; // @[ivncontrol4.scala 494:162 496:21]
  wire [31:0] _GEN_3000 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2993; // @[ivncontrol4.scala 494:162 497:21]
  wire [31:0] _GEN_3001 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2994; // @[ivncontrol4.scala 494:162 498:22]
  wire [31:0] _GEN_3002 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2995; // @[ivncontrol4.scala 494:162 499:22]
  wire [31:0] _GEN_3003 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2996; // @[ivncontrol4.scala 494:162 500:22]
  wire [31:0] _GEN_3004 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2997; // @[ivncontrol4.scala 494:162 501:22]
  wire [31:0] _GEN_3102 = 4'h1 == _i_vn_1_T_25[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3103 = 4'h2 == _i_vn_1_T_25[3:0] ? rowcount_2 : _GEN_3102; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3104 = 4'h3 == _i_vn_1_T_25[3:0] ? rowcount_3 : _GEN_3103; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3105 = 4'h4 == _i_vn_1_T_25[3:0] ? rowcount_4 : _GEN_3104; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3106 = 4'h5 == _i_vn_1_T_25[3:0] ? rowcount_5 : _GEN_3105; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3107 = 4'h6 == _i_vn_1_T_25[3:0] ? rowcount_6 : _GEN_3106; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3108 = 4'h7 == _i_vn_1_T_25[3:0] ? rowcount_7 : _GEN_3107; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3109 = 4'h8 == _i_vn_1_T_25[3:0] ? rowcount_8 : _GEN_3108; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3110 = 4'h9 == _i_vn_1_T_25[3:0] ? rowcount_9 : _GEN_3109; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3111 = 4'ha == _i_vn_1_T_25[3:0] ? rowcount_10 : _GEN_3110; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3112 = 4'hb == _i_vn_1_T_25[3:0] ? rowcount_11 : _GEN_3111; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3113 = 4'hc == _i_vn_1_T_25[3:0] ? rowcount_12 : _GEN_3112; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3114 = 4'hd == _i_vn_1_T_25[3:0] ? rowcount_13 : _GEN_3113; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3115 = 4'he == _i_vn_1_T_25[3:0] ? rowcount_14 : _GEN_3114; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3116 = 4'hf == _i_vn_1_T_25[3:0] ? rowcount_15 : _GEN_3115; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _T_932 = _T_710 + _GEN_3116; // @[ivncontrol4.scala 545:152]
  wire [31:0] _T_934 = 32'h8 - _T_932; // @[ivncontrol4.scala 545:19]
  wire [31:0] _i_vn_1_T_27 = 32'h7 + pin; // @[ivncontrol4.scala 546:29]
  wire [31:0] _GEN_3789 = _T_934 == 32'h1 ? _i_vn_1_T_27 : _GEN_3004; // @[ivncontrol4.scala 588:188 591:22]
  wire [31:0] _GEN_3790 = _T_934 == 32'h2 ? _i_vn_1_T_27 : _GEN_3003; // @[ivncontrol4.scala 582:188 585:22]
  wire [31:0] _GEN_3791 = _T_934 == 32'h2 ? _i_vn_1_T_27 : _GEN_3789; // @[ivncontrol4.scala 582:188 586:22]
  wire [31:0] _GEN_3792 = _T_934 == 32'h3 ? _i_vn_1_T_27 : _GEN_3002; // @[ivncontrol4.scala 575:190 577:23]
  wire [31:0] _GEN_3793 = _T_934 == 32'h3 ? _i_vn_1_T_27 : _GEN_3790; // @[ivncontrol4.scala 575:190 578:22]
  wire [31:0] _GEN_3794 = _T_934 == 32'h3 ? _i_vn_1_T_27 : _GEN_3791; // @[ivncontrol4.scala 575:190 579:22]
  wire [31:0] _GEN_3795 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_3001; // @[ivncontrol4.scala 569:188 571:22]
  wire [31:0] _GEN_3796 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_3792; // @[ivncontrol4.scala 569:188 572:22]
  wire [31:0] _GEN_3797 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_3793; // @[ivncontrol4.scala 569:188 573:22]
  wire [31:0] _GEN_3798 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_3794; // @[ivncontrol4.scala 569:188 574:22]
  wire [31:0] _GEN_3799 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3000; // @[ivncontrol4.scala 562:188 564:23]
  wire [31:0] _GEN_3800 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3795; // @[ivncontrol4.scala 562:188 565:22]
  wire [31:0] _GEN_3801 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3796; // @[ivncontrol4.scala 562:188 566:22]
  wire [31:0] _GEN_3802 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3797; // @[ivncontrol4.scala 562:188 567:22]
  wire [31:0] _GEN_3803 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3798; // @[ivncontrol4.scala 562:188 568:22]
  wire [31:0] _GEN_3804 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_2999; // @[ivncontrol4.scala 554:188 556:22]
  wire [31:0] _GEN_3805 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3799; // @[ivncontrol4.scala 554:188 557:21]
  wire [31:0] _GEN_3806 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3800; // @[ivncontrol4.scala 554:188 558:22]
  wire [31:0] _GEN_3807 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3801; // @[ivncontrol4.scala 554:188 559:22]
  wire [31:0] _GEN_3808 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3802; // @[ivncontrol4.scala 554:188 560:22]
  wire [31:0] _GEN_3809 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3803; // @[ivncontrol4.scala 554:188 561:22]
  wire [31:0] _GEN_3810 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_2998; // @[ivncontrol4.scala 545:184 546:22]
  wire [31:0] _GEN_3811 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3804; // @[ivncontrol4.scala 545:184 547:21]
  wire [31:0] _GEN_3812 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3805; // @[ivncontrol4.scala 545:184 548:21]
  wire [31:0] _GEN_3813 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3806; // @[ivncontrol4.scala 545:184 549:22]
  wire [31:0] _GEN_3814 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3807; // @[ivncontrol4.scala 545:184 550:22]
  wire [31:0] _GEN_3815 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3808; // @[ivncontrol4.scala 545:184 551:22]
  wire [31:0] _GEN_3816 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3809; // @[ivncontrol4.scala 545:184 552:22]
  wire [31:0] _GEN_3817 = _GEN_312 ? _GEN_477 : 32'hc; // @[ivncontrol4.scala 142:17 189:28]
  wire [31:0] _GEN_3818 = _GEN_312 ? _GEN_3810 : 32'h1; // @[ivncontrol4.scala 142:17 189:28]
  wire [31:0] _GEN_3819 = _GEN_312 ? _GEN_3811 : 32'h1a; // @[ivncontrol4.scala 142:17 189:28]
  wire [31:0] _GEN_3820 = _GEN_312 ? _GEN_3812 : 32'h1b; // @[ivncontrol4.scala 142:17 189:28]
  wire [31:0] _GEN_3821 = _GEN_312 ? _GEN_3813 : 32'h13; // @[ivncontrol4.scala 143:18 189:28]
  wire [31:0] _GEN_3822 = _GEN_312 ? _GEN_3814 : 32'ha; // @[ivncontrol4.scala 143:18 189:28]
  wire [31:0] _GEN_3823 = _GEN_312 ? _GEN_3815 : 32'h6; // @[ivncontrol4.scala 143:18 189:28]
  wire [31:0] _GEN_3824 = _GEN_312 ? _GEN_3816 : 32'h1b; // @[ivncontrol4.scala 143:18 189:28]
  wire  valid1 = 1'h0;
  wire [31:0] _GEN_4221 = reset ? 32'h0 : _GEN_3817; // @[ivncontrol4.scala 17:{23,23}]
  wire [31:0] _GEN_4222 = reset ? 32'h0 : _GEN_3818; // @[ivncontrol4.scala 17:{23,23}]
  wire [31:0] _GEN_4223 = reset ? 32'h0 : _GEN_3819; // @[ivncontrol4.scala 17:{23,23}]
  wire [31:0] _GEN_4224 = reset ? 32'h0 : _GEN_3820; // @[ivncontrol4.scala 17:{23,23}]
  wire [31:0] _GEN_4225 = reset ? 32'h0 : _GEN_3821; // @[ivncontrol4.scala 18:{24,24}]
  wire [31:0] _GEN_4226 = reset ? 32'h0 : _GEN_3822; // @[ivncontrol4.scala 18:{24,24}]
  wire [31:0] _GEN_4227 = reset ? 32'h0 : _GEN_3823; // @[ivncontrol4.scala 18:{24,24}]
  wire [31:0] _GEN_4228 = reset ? 32'h0 : _GEN_3824; // @[ivncontrol4.scala 18:{24,24}]
  assign io_o_vn_0 = i_vn_0; // @[ivncontrol4.scala 138:13]
  assign io_o_vn_1 = i_vn_1; // @[ivncontrol4.scala 138:13]
  assign io_o_vn_2 = i_vn_2; // @[ivncontrol4.scala 138:13]
  assign io_o_vn_3 = i_vn_3; // @[ivncontrol4.scala 138:13]
  assign io_o_vn2_0 = i_vn2_0; // @[ivncontrol4.scala 139:14]
  assign io_o_vn2_1 = i_vn2_1; // @[ivncontrol4.scala 139:14]
  assign io_o_vn2_2 = i_vn2_2; // @[ivncontrol4.scala 139:14]
  assign io_o_vn2_3 = i_vn2_3; // @[ivncontrol4.scala 139:14]
  always @(posedge clock) begin
    i_vn_0 <= _GEN_4221[4:0]; // @[ivncontrol4.scala 17:{23,23}]
    i_vn_1 <= _GEN_4222[4:0]; // @[ivncontrol4.scala 17:{23,23}]
    i_vn_2 <= _GEN_4223[4:0]; // @[ivncontrol4.scala 17:{23,23}]
    i_vn_3 <= _GEN_4224[4:0]; // @[ivncontrol4.scala 17:{23,23}]
    i_vn2_0 <= _GEN_4225[4:0]; // @[ivncontrol4.scala 18:{24,24}]
    i_vn2_1 <= _GEN_4226[4:0]; // @[ivncontrol4.scala 18:{24,24}]
    i_vn2_2 <= _GEN_4227[4:0]; // @[ivncontrol4.scala 18:{24,24}]
    i_vn2_3 <= _GEN_4228[4:0]; // @[ivncontrol4.scala 18:{24,24}]
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_0 <= io_Stationary_matrix_0_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_1 <= io_Stationary_matrix_0_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_2 <= io_Stationary_matrix_0_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_3 <= io_Stationary_matrix_0_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_4 <= io_Stationary_matrix_0_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_5 <= io_Stationary_matrix_0_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_6 <= io_Stationary_matrix_0_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_7 <= io_Stationary_matrix_0_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_0 <= io_Stationary_matrix_1_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_1 <= io_Stationary_matrix_1_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_2 <= io_Stationary_matrix_1_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_3 <= io_Stationary_matrix_1_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_4 <= io_Stationary_matrix_1_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_5 <= io_Stationary_matrix_1_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_6 <= io_Stationary_matrix_1_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_7 <= io_Stationary_matrix_1_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_0 <= io_Stationary_matrix_2_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_1 <= io_Stationary_matrix_2_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_2 <= io_Stationary_matrix_2_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_3 <= io_Stationary_matrix_2_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_4 <= io_Stationary_matrix_2_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_5 <= io_Stationary_matrix_2_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_6 <= io_Stationary_matrix_2_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_7 <= io_Stationary_matrix_2_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_0 <= io_Stationary_matrix_3_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_1 <= io_Stationary_matrix_3_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_2 <= io_Stationary_matrix_3_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_3 <= io_Stationary_matrix_3_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_4 <= io_Stationary_matrix_3_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_5 <= io_Stationary_matrix_3_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_6 <= io_Stationary_matrix_3_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_7 <= io_Stationary_matrix_3_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_0 <= io_Stationary_matrix_4_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_1 <= io_Stationary_matrix_4_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_2 <= io_Stationary_matrix_4_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_3 <= io_Stationary_matrix_4_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_4 <= io_Stationary_matrix_4_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_5 <= io_Stationary_matrix_4_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_6 <= io_Stationary_matrix_4_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_7 <= io_Stationary_matrix_4_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_0 <= io_Stationary_matrix_5_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_1 <= io_Stationary_matrix_5_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_2 <= io_Stationary_matrix_5_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_3 <= io_Stationary_matrix_5_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_4 <= io_Stationary_matrix_5_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_5 <= io_Stationary_matrix_5_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_6 <= io_Stationary_matrix_5_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_7 <= io_Stationary_matrix_5_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_0 <= io_Stationary_matrix_6_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_1 <= io_Stationary_matrix_6_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_2 <= io_Stationary_matrix_6_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_3 <= io_Stationary_matrix_6_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_4 <= io_Stationary_matrix_6_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_5 <= io_Stationary_matrix_6_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_6 <= io_Stationary_matrix_6_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_7 <= io_Stationary_matrix_6_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_0 <= io_Stationary_matrix_7_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_1 <= io_Stationary_matrix_7_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_2 <= io_Stationary_matrix_7_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_3 <= io_Stationary_matrix_7_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_4 <= io_Stationary_matrix_7_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_5 <= io_Stationary_matrix_7_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_6 <= io_Stationary_matrix_7_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_7 <= io_Stationary_matrix_7_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_0 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_0 <= count_0; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_1 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_1 <= count_1; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_2 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_2 <= count_2; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_3 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_3 <= count_3; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_4 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_4 <= count_4; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_5 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_5 <= count_5; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_6 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_6 <= count_6; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_7 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_7 <= count_7; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_8 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_8 <= 32'h0; // @[ivncontrol4.scala 87:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_9 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_9 <= 32'h0; // @[ivncontrol4.scala 87:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_10 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_10 <= 32'h0; // @[ivncontrol4.scala 87:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_11 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_11 <= 32'h0; // @[ivncontrol4.scala 87:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_12 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_12 <= 32'h0; // @[ivncontrol4.scala 87:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_13 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_13 <= 32'h0; // @[ivncontrol4.scala 87:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_14 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_14 <= 32'h0; // @[ivncontrol4.scala 87:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_15 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end
    if (reset) begin // @[ivncontrol4.scala 37:22]
      pin <= 32'h0; // @[ivncontrol4.scala 37:22]
    end else if (_T_72 & rowcount_6 == 32'h0 & rowcount_7 != 32'h0) begin // @[ivncontrol4.scala 183:192]
      pin <= 32'h7; // @[ivncontrol4.scala 184:13]
    end else if (_T_59 & rowcount_5 == 32'h0 & rowcount_6 != 32'h0) begin // @[ivncontrol4.scala 180:169]
      pin <= 32'h6; // @[ivncontrol4.scala 181:13]
    end else if (_T_48 & rowcount_4 == 32'h0 & rowcount_5 != 32'h0) begin // @[ivncontrol4.scala 177:146]
      pin <= 32'h5; // @[ivncontrol4.scala 178:13]
    end else begin
      pin <= _GEN_317;
    end
    if (reset) begin // @[ivncontrol4.scala 41:20]
      i <= 32'h0; // @[ivncontrol4.scala 41:20]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
        i <= _GEN_247;
      end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
        i <= _GEN_247;
      end else begin
        i <= _GEN_265;
      end
    end
    if (reset) begin // @[ivncontrol4.scala 42:20]
      j <= 32'h0; // @[ivncontrol4.scala 42:20]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
        j <= 32'h8; // @[ivncontrol4.scala 116:11]
      end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
        j <= _j_T_1; // @[ivncontrol4.scala 118:11]
      end else begin
        j <= {{28'd0}, _GEN_264};
      end
    end
    if (3'h0 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h0 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h0 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h0 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h0 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h0 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h0 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h0 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_0 <= _GEN_224;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_0 <= _GEN_224;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h0 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_0 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_0 <= _GEN_224;
      end
    end else begin
      count_0 <= _GEN_224;
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_1 <= _GEN_225;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_1 <= _GEN_225;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h1 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_1 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_1 <= _GEN_225;
      end
    end else begin
      count_1 <= _GEN_225;
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_2 <= _GEN_226;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_2 <= _GEN_226;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h2 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_2 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_2 <= _GEN_226;
      end
    end else begin
      count_2 <= _GEN_226;
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_3 <= _GEN_227;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_3 <= _GEN_227;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h3 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_3 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_3 <= _GEN_227;
      end
    end else begin
      count_3 <= _GEN_227;
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_4 <= _GEN_228;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_4 <= _GEN_228;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h4 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_4 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_4 <= _GEN_228;
      end
    end else begin
      count_4 <= _GEN_228;
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_5 <= _GEN_229;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_5 <= _GEN_229;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h5 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_5 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_5 <= _GEN_229;
      end
    end else begin
      count_5 <= _GEN_229;
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_6 <= _GEN_230;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_6 <= _GEN_230;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h6 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_6 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_6 <= _GEN_230;
      end
    end else begin
      count_6 <= _GEN_230;
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_7 <= _GEN_231;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_7 <= _GEN_231;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h7 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_7 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_7 <= _GEN_231;
      end
    end else begin
      count_7 <= _GEN_231;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  i_vn_0 = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  i_vn_1 = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  i_vn_2 = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  i_vn_3 = _RAND_3[4:0];
  _RAND_4 = {1{`RANDOM}};
  i_vn2_0 = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  i_vn2_1 = _RAND_5[4:0];
  _RAND_6 = {1{`RANDOM}};
  i_vn2_2 = _RAND_6[4:0];
  _RAND_7 = {1{`RANDOM}};
  i_vn2_3 = _RAND_7[4:0];
  _RAND_8 = {1{`RANDOM}};
  solution_0_0 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  solution_0_1 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  solution_0_2 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  solution_0_3 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  solution_0_4 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  solution_0_5 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  solution_0_6 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  solution_0_7 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  solution_1_0 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  solution_1_1 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  solution_1_2 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  solution_1_3 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  solution_1_4 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  solution_1_5 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  solution_1_6 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  solution_1_7 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  solution_2_0 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  solution_2_1 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  solution_2_2 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  solution_2_3 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  solution_2_4 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  solution_2_5 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  solution_2_6 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  solution_2_7 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  solution_3_0 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  solution_3_1 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  solution_3_2 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  solution_3_3 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  solution_3_4 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  solution_3_5 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  solution_3_6 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  solution_3_7 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  solution_4_0 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  solution_4_1 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  solution_4_2 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  solution_4_3 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  solution_4_4 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  solution_4_5 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  solution_4_6 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  solution_4_7 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  solution_5_0 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  solution_5_1 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  solution_5_2 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  solution_5_3 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  solution_5_4 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  solution_5_5 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  solution_5_6 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  solution_5_7 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  solution_6_0 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  solution_6_1 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  solution_6_2 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  solution_6_3 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  solution_6_4 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  solution_6_5 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  solution_6_6 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  solution_6_7 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  solution_7_0 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  solution_7_1 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  solution_7_2 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  solution_7_3 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  solution_7_4 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  solution_7_5 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  solution_7_6 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  solution_7_7 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  rowcount_0 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  rowcount_1 = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  rowcount_2 = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  rowcount_3 = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  rowcount_4 = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  rowcount_5 = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  rowcount_6 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  rowcount_7 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  rowcount_8 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  rowcount_9 = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  rowcount_10 = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  rowcount_11 = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  rowcount_12 = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  rowcount_13 = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  rowcount_14 = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  rowcount_15 = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  pin = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  i = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  j = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  mat_0_0 = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  mat_0_1 = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  mat_0_2 = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  mat_0_3 = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  mat_0_4 = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  mat_0_5 = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  mat_0_6 = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  mat_0_7 = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  mat_1_0 = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  mat_1_1 = _RAND_100[31:0];
  _RAND_101 = {1{`RANDOM}};
  mat_1_2 = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  mat_1_3 = _RAND_102[31:0];
  _RAND_103 = {1{`RANDOM}};
  mat_1_4 = _RAND_103[31:0];
  _RAND_104 = {1{`RANDOM}};
  mat_1_5 = _RAND_104[31:0];
  _RAND_105 = {1{`RANDOM}};
  mat_1_6 = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  mat_1_7 = _RAND_106[31:0];
  _RAND_107 = {1{`RANDOM}};
  mat_2_0 = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  mat_2_1 = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  mat_2_2 = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  mat_2_3 = _RAND_110[31:0];
  _RAND_111 = {1{`RANDOM}};
  mat_2_4 = _RAND_111[31:0];
  _RAND_112 = {1{`RANDOM}};
  mat_2_5 = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  mat_2_6 = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  mat_2_7 = _RAND_114[31:0];
  _RAND_115 = {1{`RANDOM}};
  mat_3_0 = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  mat_3_1 = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  mat_3_2 = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  mat_3_3 = _RAND_118[31:0];
  _RAND_119 = {1{`RANDOM}};
  mat_3_4 = _RAND_119[31:0];
  _RAND_120 = {1{`RANDOM}};
  mat_3_5 = _RAND_120[31:0];
  _RAND_121 = {1{`RANDOM}};
  mat_3_6 = _RAND_121[31:0];
  _RAND_122 = {1{`RANDOM}};
  mat_3_7 = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  mat_4_0 = _RAND_123[31:0];
  _RAND_124 = {1{`RANDOM}};
  mat_4_1 = _RAND_124[31:0];
  _RAND_125 = {1{`RANDOM}};
  mat_4_2 = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  mat_4_3 = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  mat_4_4 = _RAND_127[31:0];
  _RAND_128 = {1{`RANDOM}};
  mat_4_5 = _RAND_128[31:0];
  _RAND_129 = {1{`RANDOM}};
  mat_4_6 = _RAND_129[31:0];
  _RAND_130 = {1{`RANDOM}};
  mat_4_7 = _RAND_130[31:0];
  _RAND_131 = {1{`RANDOM}};
  mat_5_0 = _RAND_131[31:0];
  _RAND_132 = {1{`RANDOM}};
  mat_5_1 = _RAND_132[31:0];
  _RAND_133 = {1{`RANDOM}};
  mat_5_2 = _RAND_133[31:0];
  _RAND_134 = {1{`RANDOM}};
  mat_5_3 = _RAND_134[31:0];
  _RAND_135 = {1{`RANDOM}};
  mat_5_4 = _RAND_135[31:0];
  _RAND_136 = {1{`RANDOM}};
  mat_5_5 = _RAND_136[31:0];
  _RAND_137 = {1{`RANDOM}};
  mat_5_6 = _RAND_137[31:0];
  _RAND_138 = {1{`RANDOM}};
  mat_5_7 = _RAND_138[31:0];
  _RAND_139 = {1{`RANDOM}};
  mat_6_0 = _RAND_139[31:0];
  _RAND_140 = {1{`RANDOM}};
  mat_6_1 = _RAND_140[31:0];
  _RAND_141 = {1{`RANDOM}};
  mat_6_2 = _RAND_141[31:0];
  _RAND_142 = {1{`RANDOM}};
  mat_6_3 = _RAND_142[31:0];
  _RAND_143 = {1{`RANDOM}};
  mat_6_4 = _RAND_143[31:0];
  _RAND_144 = {1{`RANDOM}};
  mat_6_5 = _RAND_144[31:0];
  _RAND_145 = {1{`RANDOM}};
  mat_6_6 = _RAND_145[31:0];
  _RAND_146 = {1{`RANDOM}};
  mat_6_7 = _RAND_146[31:0];
  _RAND_147 = {1{`RANDOM}};
  mat_7_0 = _RAND_147[31:0];
  _RAND_148 = {1{`RANDOM}};
  mat_7_1 = _RAND_148[31:0];
  _RAND_149 = {1{`RANDOM}};
  mat_7_2 = _RAND_149[31:0];
  _RAND_150 = {1{`RANDOM}};
  mat_7_3 = _RAND_150[31:0];
  _RAND_151 = {1{`RANDOM}};
  mat_7_4 = _RAND_151[31:0];
  _RAND_152 = {1{`RANDOM}};
  mat_7_5 = _RAND_152[31:0];
  _RAND_153 = {1{`RANDOM}};
  mat_7_6 = _RAND_153[31:0];
  _RAND_154 = {1{`RANDOM}};
  mat_7_7 = _RAND_154[31:0];
  _RAND_155 = {1{`RANDOM}};
  count_0 = _RAND_155[31:0];
  _RAND_156 = {1{`RANDOM}};
  count_1 = _RAND_156[31:0];
  _RAND_157 = {1{`RANDOM}};
  count_2 = _RAND_157[31:0];
  _RAND_158 = {1{`RANDOM}};
  count_3 = _RAND_158[31:0];
  _RAND_159 = {1{`RANDOM}};
  count_4 = _RAND_159[31:0];
  _RAND_160 = {1{`RANDOM}};
  count_5 = _RAND_160[31:0];
  _RAND_161 = {1{`RANDOM}};
  count_6 = _RAND_161[31:0];
  _RAND_162 = {1{`RANDOM}};
  count_7 = _RAND_162[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ivncontrol4_7(
  input         clock,
  input         reset,
  input  [15:0] io_Stationary_matrix_0_0,
  input  [15:0] io_Stationary_matrix_0_1,
  input  [15:0] io_Stationary_matrix_0_2,
  input  [15:0] io_Stationary_matrix_0_3,
  input  [15:0] io_Stationary_matrix_0_4,
  input  [15:0] io_Stationary_matrix_0_5,
  input  [15:0] io_Stationary_matrix_0_6,
  input  [15:0] io_Stationary_matrix_0_7,
  input  [15:0] io_Stationary_matrix_1_0,
  input  [15:0] io_Stationary_matrix_1_1,
  input  [15:0] io_Stationary_matrix_1_2,
  input  [15:0] io_Stationary_matrix_1_3,
  input  [15:0] io_Stationary_matrix_1_4,
  input  [15:0] io_Stationary_matrix_1_5,
  input  [15:0] io_Stationary_matrix_1_6,
  input  [15:0] io_Stationary_matrix_1_7,
  input  [15:0] io_Stationary_matrix_2_0,
  input  [15:0] io_Stationary_matrix_2_1,
  input  [15:0] io_Stationary_matrix_2_2,
  input  [15:0] io_Stationary_matrix_2_3,
  input  [15:0] io_Stationary_matrix_2_4,
  input  [15:0] io_Stationary_matrix_2_5,
  input  [15:0] io_Stationary_matrix_2_6,
  input  [15:0] io_Stationary_matrix_2_7,
  input  [15:0] io_Stationary_matrix_3_0,
  input  [15:0] io_Stationary_matrix_3_1,
  input  [15:0] io_Stationary_matrix_3_2,
  input  [15:0] io_Stationary_matrix_3_3,
  input  [15:0] io_Stationary_matrix_3_4,
  input  [15:0] io_Stationary_matrix_3_5,
  input  [15:0] io_Stationary_matrix_3_6,
  input  [15:0] io_Stationary_matrix_3_7,
  input  [15:0] io_Stationary_matrix_4_0,
  input  [15:0] io_Stationary_matrix_4_1,
  input  [15:0] io_Stationary_matrix_4_2,
  input  [15:0] io_Stationary_matrix_4_3,
  input  [15:0] io_Stationary_matrix_4_4,
  input  [15:0] io_Stationary_matrix_4_5,
  input  [15:0] io_Stationary_matrix_4_6,
  input  [15:0] io_Stationary_matrix_4_7,
  input  [15:0] io_Stationary_matrix_5_0,
  input  [15:0] io_Stationary_matrix_5_1,
  input  [15:0] io_Stationary_matrix_5_2,
  input  [15:0] io_Stationary_matrix_5_3,
  input  [15:0] io_Stationary_matrix_5_4,
  input  [15:0] io_Stationary_matrix_5_5,
  input  [15:0] io_Stationary_matrix_5_6,
  input  [15:0] io_Stationary_matrix_5_7,
  input  [15:0] io_Stationary_matrix_6_0,
  input  [15:0] io_Stationary_matrix_6_1,
  input  [15:0] io_Stationary_matrix_6_2,
  input  [15:0] io_Stationary_matrix_6_3,
  input  [15:0] io_Stationary_matrix_6_4,
  input  [15:0] io_Stationary_matrix_6_5,
  input  [15:0] io_Stationary_matrix_6_6,
  input  [15:0] io_Stationary_matrix_6_7,
  input  [15:0] io_Stationary_matrix_7_0,
  input  [15:0] io_Stationary_matrix_7_1,
  input  [15:0] io_Stationary_matrix_7_2,
  input  [15:0] io_Stationary_matrix_7_3,
  input  [15:0] io_Stationary_matrix_7_4,
  input  [15:0] io_Stationary_matrix_7_5,
  input  [15:0] io_Stationary_matrix_7_6,
  input  [15:0] io_Stationary_matrix_7_7,
  output [4:0]  io_o_vn_0,
  output [4:0]  io_o_vn_1,
  output [4:0]  io_o_vn_2,
  output [4:0]  io_o_vn_3,
  output [4:0]  io_o_vn2_0,
  output [4:0]  io_o_vn2_1,
  output [4:0]  io_o_vn2_2,
  output [4:0]  io_o_vn2_3,
  input         io_validpin
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
`endif // RANDOMIZE_REG_INIT
  reg [4:0] i_vn_0; // @[ivncontrol4.scala 17:23]
  reg [4:0] i_vn_1; // @[ivncontrol4.scala 17:23]
  reg [4:0] i_vn_2; // @[ivncontrol4.scala 17:23]
  reg [4:0] i_vn_3; // @[ivncontrol4.scala 17:23]
  reg [4:0] i_vn2_0; // @[ivncontrol4.scala 18:24]
  reg [4:0] i_vn2_1; // @[ivncontrol4.scala 18:24]
  reg [4:0] i_vn2_2; // @[ivncontrol4.scala 18:24]
  reg [4:0] i_vn2_3; // @[ivncontrol4.scala 18:24]
  reg [15:0] solution_0_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_0_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_0_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_0_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_0_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_0_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_0_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_0_7; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_1_7; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_2_7; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_3_7; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_4_7; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_5_7; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_6_7; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_0; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_1; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_2; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_3; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_4; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_5; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_6; // @[ivncontrol4.scala 21:27]
  reg [15:0] solution_7_7; // @[ivncontrol4.scala 21:27]
  reg [31:0] rowcount_0; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_1; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_2; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_3; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_4; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_5; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_6; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_7; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_8; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_9; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_10; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_11; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_12; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_13; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_14; // @[ivncontrol4.scala 27:27]
  reg [31:0] rowcount_15; // @[ivncontrol4.scala 27:27]
  reg [31:0] pin; // @[ivncontrol4.scala 37:22]
  reg [31:0] i; // @[ivncontrol4.scala 41:20]
  reg [31:0] j; // @[ivncontrol4.scala 42:20]
  wire  _io_ProcessValid_T = i == 32'h7; // @[ivncontrol4.scala 44:27]
  wire  _io_ProcessValid_T_1 = j == 32'h7; // @[ivncontrol4.scala 44:42]
  wire  _io_ProcessValid_T_2 = i == 32'h7 & j == 32'h7; // @[ivncontrol4.scala 44:36]
  reg [31:0] mat_0_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_0_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_0_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_0_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_0_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_0_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_0_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_0_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_1_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_2_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_3_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_4_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_5_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_6_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_0; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_1; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_2; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_3; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_4; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_5; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_6; // @[ivncontrol4.scala 54:18]
  reg [31:0] mat_7_7; // @[ivncontrol4.scala 54:18]
  reg [31:0] count_0; // @[ivncontrol4.scala 58:20]
  reg [31:0] count_1; // @[ivncontrol4.scala 58:20]
  reg [31:0] count_2; // @[ivncontrol4.scala 58:20]
  reg [31:0] count_3; // @[ivncontrol4.scala 58:20]
  reg [31:0] count_4; // @[ivncontrol4.scala 58:20]
  reg [31:0] count_5; // @[ivncontrol4.scala 58:20]
  reg [31:0] count_6; // @[ivncontrol4.scala 58:20]
  reg [31:0] count_7; // @[ivncontrol4.scala 58:20]
  wire  _GEN_3825 = 3'h0 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_65 = 3'h0 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_0_1 : io_Stationary_matrix_0_0; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_66 = 3'h0 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_0_2 : _GEN_65; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_67 = 3'h0 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_0_3 : _GEN_66; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_68 = 3'h0 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_0_4 : _GEN_67; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_69 = 3'h0 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_0_5 : _GEN_68; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_70 = 3'h0 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_0_6 : _GEN_69; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_71 = 3'h0 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_0_7 : _GEN_70; // @[ivncontrol4.scala 63:{17,17}]
  wire  _GEN_3839 = 3'h1 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_72 = 3'h1 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_1_0 : _GEN_71; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_73 = 3'h1 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_1_1 : _GEN_72; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_74 = 3'h1 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_1_2 : _GEN_73; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_75 = 3'h1 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_1_3 : _GEN_74; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_76 = 3'h1 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_1_4 : _GEN_75; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_77 = 3'h1 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_1_5 : _GEN_76; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_78 = 3'h1 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_1_6 : _GEN_77; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_79 = 3'h1 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_1_7 : _GEN_78; // @[ivncontrol4.scala 63:{17,17}]
  wire  _GEN_3855 = 3'h2 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_80 = 3'h2 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_2_0 : _GEN_79; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_81 = 3'h2 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_2_1 : _GEN_80; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_82 = 3'h2 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_2_2 : _GEN_81; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_83 = 3'h2 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_2_3 : _GEN_82; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_84 = 3'h2 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_2_4 : _GEN_83; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_85 = 3'h2 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_2_5 : _GEN_84; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_86 = 3'h2 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_2_6 : _GEN_85; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_87 = 3'h2 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_2_7 : _GEN_86; // @[ivncontrol4.scala 63:{17,17}]
  wire  _GEN_3871 = 3'h3 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_88 = 3'h3 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_3_0 : _GEN_87; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_89 = 3'h3 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_3_1 : _GEN_88; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_90 = 3'h3 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_3_2 : _GEN_89; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_91 = 3'h3 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_3_3 : _GEN_90; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_92 = 3'h3 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_3_4 : _GEN_91; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_93 = 3'h3 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_3_5 : _GEN_92; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_94 = 3'h3 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_3_6 : _GEN_93; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_95 = 3'h3 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_3_7 : _GEN_94; // @[ivncontrol4.scala 63:{17,17}]
  wire  _GEN_3887 = 3'h4 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_96 = 3'h4 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_4_0 : _GEN_95; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_97 = 3'h4 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_4_1 : _GEN_96; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_98 = 3'h4 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_4_2 : _GEN_97; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_99 = 3'h4 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_4_3 : _GEN_98; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_100 = 3'h4 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_4_4 : _GEN_99; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_101 = 3'h4 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_4_5 : _GEN_100; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_102 = 3'h4 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_4_6 : _GEN_101; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_103 = 3'h4 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_4_7 : _GEN_102; // @[ivncontrol4.scala 63:{17,17}]
  wire  _GEN_3903 = 3'h5 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_104 = 3'h5 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_5_0 : _GEN_103; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_105 = 3'h5 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_5_1 : _GEN_104; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_106 = 3'h5 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_5_2 : _GEN_105; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_107 = 3'h5 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_5_3 : _GEN_106; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_108 = 3'h5 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_5_4 : _GEN_107; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_109 = 3'h5 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_5_5 : _GEN_108; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_110 = 3'h5 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_5_6 : _GEN_109; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_111 = 3'h5 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_5_7 : _GEN_110; // @[ivncontrol4.scala 63:{17,17}]
  wire  _GEN_3919 = 3'h6 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_112 = 3'h6 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_6_0 : _GEN_111; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_113 = 3'h6 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_6_1 : _GEN_112; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_114 = 3'h6 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_6_2 : _GEN_113; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_115 = 3'h6 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_6_3 : _GEN_114; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_116 = 3'h6 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_6_4 : _GEN_115; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_117 = 3'h6 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_6_5 : _GEN_116; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_118 = 3'h6 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_6_6 : _GEN_117; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_119 = 3'h6 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_6_7 : _GEN_118; // @[ivncontrol4.scala 63:{17,17}]
  wire  _GEN_3935 = 3'h7 == i[2:0]; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_120 = 3'h7 == i[2:0] & 3'h0 == j[2:0] ? io_Stationary_matrix_7_0 : _GEN_119; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_121 = 3'h7 == i[2:0] & 3'h1 == j[2:0] ? io_Stationary_matrix_7_1 : _GEN_120; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_122 = 3'h7 == i[2:0] & 3'h2 == j[2:0] ? io_Stationary_matrix_7_2 : _GEN_121; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_123 = 3'h7 == i[2:0] & 3'h3 == j[2:0] ? io_Stationary_matrix_7_3 : _GEN_122; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_124 = 3'h7 == i[2:0] & 3'h4 == j[2:0] ? io_Stationary_matrix_7_4 : _GEN_123; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_125 = 3'h7 == i[2:0] & 3'h5 == j[2:0] ? io_Stationary_matrix_7_5 : _GEN_124; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_126 = 3'h7 == i[2:0] & 3'h6 == j[2:0] ? io_Stationary_matrix_7_6 : _GEN_125; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_127 = 3'h7 == i[2:0] & 3'h7 == j[2:0] ? io_Stationary_matrix_7_7 : _GEN_126; // @[ivncontrol4.scala 63:{17,17}]
  wire [31:0] _mat_T_1_T_2 = {{16'd0}, _GEN_127}; // @[ivncontrol4.scala 63:{17,17}]
  wire [15:0] _GEN_129 = _GEN_3825 & 4'h1 == j[3:0] ? solution_0_1 : solution_0_0; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_130 = _GEN_3825 & 4'h2 == j[3:0] ? solution_0_2 : _GEN_129; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_131 = _GEN_3825 & 4'h3 == j[3:0] ? solution_0_3 : _GEN_130; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_132 = _GEN_3825 & 4'h4 == j[3:0] ? solution_0_4 : _GEN_131; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_133 = _GEN_3825 & 4'h5 == j[3:0] ? solution_0_5 : _GEN_132; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_134 = _GEN_3825 & 4'h6 == j[3:0] ? solution_0_6 : _GEN_133; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_135 = _GEN_3825 & 4'h7 == j[3:0] ? solution_0_7 : _GEN_134; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_136 = _GEN_3825 & 4'h8 == j[3:0] ? 16'h0 : _GEN_135; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_137 = _GEN_3839 & 4'h0 == j[3:0] ? solution_1_0 : _GEN_136; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_138 = _GEN_3839 & 4'h1 == j[3:0] ? solution_1_1 : _GEN_137; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_139 = _GEN_3839 & 4'h2 == j[3:0] ? solution_1_2 : _GEN_138; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_140 = _GEN_3839 & 4'h3 == j[3:0] ? solution_1_3 : _GEN_139; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_141 = _GEN_3839 & 4'h4 == j[3:0] ? solution_1_4 : _GEN_140; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_142 = _GEN_3839 & 4'h5 == j[3:0] ? solution_1_5 : _GEN_141; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_143 = _GEN_3839 & 4'h6 == j[3:0] ? solution_1_6 : _GEN_142; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_144 = _GEN_3839 & 4'h7 == j[3:0] ? solution_1_7 : _GEN_143; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_145 = _GEN_3839 & 4'h8 == j[3:0] ? 16'h0 : _GEN_144; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_146 = _GEN_3855 & 4'h0 == j[3:0] ? solution_2_0 : _GEN_145; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_147 = _GEN_3855 & 4'h1 == j[3:0] ? solution_2_1 : _GEN_146; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_148 = _GEN_3855 & 4'h2 == j[3:0] ? solution_2_2 : _GEN_147; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_149 = _GEN_3855 & 4'h3 == j[3:0] ? solution_2_3 : _GEN_148; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_150 = _GEN_3855 & 4'h4 == j[3:0] ? solution_2_4 : _GEN_149; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_151 = _GEN_3855 & 4'h5 == j[3:0] ? solution_2_5 : _GEN_150; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_152 = _GEN_3855 & 4'h6 == j[3:0] ? solution_2_6 : _GEN_151; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_153 = _GEN_3855 & 4'h7 == j[3:0] ? solution_2_7 : _GEN_152; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_154 = _GEN_3855 & 4'h8 == j[3:0] ? 16'h0 : _GEN_153; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_155 = _GEN_3871 & 4'h0 == j[3:0] ? solution_3_0 : _GEN_154; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_156 = _GEN_3871 & 4'h1 == j[3:0] ? solution_3_1 : _GEN_155; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_157 = _GEN_3871 & 4'h2 == j[3:0] ? solution_3_2 : _GEN_156; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_158 = _GEN_3871 & 4'h3 == j[3:0] ? solution_3_3 : _GEN_157; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_159 = _GEN_3871 & 4'h4 == j[3:0] ? solution_3_4 : _GEN_158; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_160 = _GEN_3871 & 4'h5 == j[3:0] ? solution_3_5 : _GEN_159; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_161 = _GEN_3871 & 4'h6 == j[3:0] ? solution_3_6 : _GEN_160; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_162 = _GEN_3871 & 4'h7 == j[3:0] ? solution_3_7 : _GEN_161; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_163 = _GEN_3871 & 4'h8 == j[3:0] ? 16'h0 : _GEN_162; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_164 = _GEN_3887 & 4'h0 == j[3:0] ? solution_4_0 : _GEN_163; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_165 = _GEN_3887 & 4'h1 == j[3:0] ? solution_4_1 : _GEN_164; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_166 = _GEN_3887 & 4'h2 == j[3:0] ? solution_4_2 : _GEN_165; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_167 = _GEN_3887 & 4'h3 == j[3:0] ? solution_4_3 : _GEN_166; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_168 = _GEN_3887 & 4'h4 == j[3:0] ? solution_4_4 : _GEN_167; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_169 = _GEN_3887 & 4'h5 == j[3:0] ? solution_4_5 : _GEN_168; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_170 = _GEN_3887 & 4'h6 == j[3:0] ? solution_4_6 : _GEN_169; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_171 = _GEN_3887 & 4'h7 == j[3:0] ? solution_4_7 : _GEN_170; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_172 = _GEN_3887 & 4'h8 == j[3:0] ? 16'h0 : _GEN_171; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_173 = _GEN_3903 & 4'h0 == j[3:0] ? solution_5_0 : _GEN_172; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_174 = _GEN_3903 & 4'h1 == j[3:0] ? solution_5_1 : _GEN_173; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_175 = _GEN_3903 & 4'h2 == j[3:0] ? solution_5_2 : _GEN_174; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_176 = _GEN_3903 & 4'h3 == j[3:0] ? solution_5_3 : _GEN_175; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_177 = _GEN_3903 & 4'h4 == j[3:0] ? solution_5_4 : _GEN_176; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_178 = _GEN_3903 & 4'h5 == j[3:0] ? solution_5_5 : _GEN_177; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_179 = _GEN_3903 & 4'h6 == j[3:0] ? solution_5_6 : _GEN_178; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_180 = _GEN_3903 & 4'h7 == j[3:0] ? solution_5_7 : _GEN_179; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_181 = _GEN_3903 & 4'h8 == j[3:0] ? 16'h0 : _GEN_180; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_182 = _GEN_3919 & 4'h0 == j[3:0] ? solution_6_0 : _GEN_181; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_183 = _GEN_3919 & 4'h1 == j[3:0] ? solution_6_1 : _GEN_182; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_184 = _GEN_3919 & 4'h2 == j[3:0] ? solution_6_2 : _GEN_183; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_185 = _GEN_3919 & 4'h3 == j[3:0] ? solution_6_3 : _GEN_184; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_186 = _GEN_3919 & 4'h4 == j[3:0] ? solution_6_4 : _GEN_185; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_187 = _GEN_3919 & 4'h5 == j[3:0] ? solution_6_5 : _GEN_186; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_188 = _GEN_3919 & 4'h6 == j[3:0] ? solution_6_6 : _GEN_187; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_189 = _GEN_3919 & 4'h7 == j[3:0] ? solution_6_7 : _GEN_188; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_190 = _GEN_3919 & 4'h8 == j[3:0] ? 16'h0 : _GEN_189; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_191 = _GEN_3935 & 4'h0 == j[3:0] ? solution_7_0 : _GEN_190; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_192 = _GEN_3935 & 4'h1 == j[3:0] ? solution_7_1 : _GEN_191; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_193 = _GEN_3935 & 4'h2 == j[3:0] ? solution_7_2 : _GEN_192; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_194 = _GEN_3935 & 4'h3 == j[3:0] ? solution_7_3 : _GEN_193; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_195 = _GEN_3935 & 4'h4 == j[3:0] ? solution_7_4 : _GEN_194; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_196 = _GEN_3935 & 4'h5 == j[3:0] ? solution_7_5 : _GEN_195; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_197 = _GEN_3935 & 4'h6 == j[3:0] ? solution_7_6 : _GEN_196; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_198 = _GEN_3935 & 4'h7 == j[3:0] ? solution_7_7 : _GEN_197; // @[ivncontrol4.scala 65:{31,31}]
  wire [15:0] _GEN_199 = _GEN_3935 & 4'h8 == j[3:0] ? 16'h0 : _GEN_198; // @[ivncontrol4.scala 65:{31,31}]
  wire [31:0] _GEN_201 = 3'h1 == i[2:0] ? count_1 : count_0; // @[ivncontrol4.scala 66:{33,33}]
  wire [31:0] _GEN_202 = 3'h2 == i[2:0] ? count_2 : _GEN_201; // @[ivncontrol4.scala 66:{33,33}]
  wire [31:0] _GEN_203 = 3'h3 == i[2:0] ? count_3 : _GEN_202; // @[ivncontrol4.scala 66:{33,33}]
  wire [31:0] _GEN_204 = 3'h4 == i[2:0] ? count_4 : _GEN_203; // @[ivncontrol4.scala 66:{33,33}]
  wire [31:0] _GEN_205 = 3'h5 == i[2:0] ? count_5 : _GEN_204; // @[ivncontrol4.scala 66:{33,33}]
  wire [31:0] _GEN_206 = 3'h6 == i[2:0] ? count_6 : _GEN_205; // @[ivncontrol4.scala 66:{33,33}]
  wire [31:0] _GEN_207 = 3'h7 == i[2:0] ? count_7 : _GEN_206; // @[ivncontrol4.scala 66:{33,33}]
  wire [31:0] _count_T_2 = _GEN_207 + 32'h1; // @[ivncontrol4.scala 66:33]
  wire [31:0] _GEN_208 = 3'h0 == i[2:0] ? _count_T_2 : count_0; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_209 = 3'h1 == i[2:0] ? _count_T_2 : count_1; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_210 = 3'h2 == i[2:0] ? _count_T_2 : count_2; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_211 = 3'h3 == i[2:0] ? _count_T_2 : count_3; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_212 = 3'h4 == i[2:0] ? _count_T_2 : count_4; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_213 = 3'h5 == i[2:0] ? _count_T_2 : count_5; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_214 = 3'h6 == i[2:0] ? _count_T_2 : count_6; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_215 = 3'h7 == i[2:0] ? _count_T_2 : count_7; // @[ivncontrol4.scala 58:20 66:{22,22}]
  wire [31:0] _GEN_216 = _GEN_199 != 16'h0 ? _GEN_208 : count_0; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_217 = _GEN_199 != 16'h0 ? _GEN_209 : count_1; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_218 = _GEN_199 != 16'h0 ? _GEN_210 : count_2; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_219 = _GEN_199 != 16'h0 ? _GEN_211 : count_3; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_220 = _GEN_199 != 16'h0 ? _GEN_212 : count_4; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_221 = _GEN_199 != 16'h0 ? _GEN_213 : count_5; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_222 = _GEN_199 != 16'h0 ? _GEN_214 : count_6; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_223 = _GEN_199 != 16'h0 ? _GEN_215 : count_7; // @[ivncontrol4.scala 58:20 65:39]
  wire [31:0] _GEN_224 = io_validpin ? _GEN_216 : count_0; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _GEN_225 = io_validpin ? _GEN_217 : count_1; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _GEN_226 = io_validpin ? _GEN_218 : count_2; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _GEN_227 = io_validpin ? _GEN_219 : count_3; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _GEN_228 = io_validpin ? _GEN_220 : count_4; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _GEN_229 = io_validpin ? _GEN_221 : count_5; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _GEN_230 = io_validpin ? _GEN_222 : count_6; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _GEN_231 = io_validpin ? _GEN_223 : count_7; // @[ivncontrol4.scala 58:20 64:22]
  wire [31:0] _i_T_1 = i + 32'h1; // @[ivncontrol4.scala 113:16]
  wire [31:0] _GEN_247 = i < 32'h7 & _io_ProcessValid_T_1 ? _i_T_1 : i; // @[ivncontrol4.scala 112:74 113:11 41:20]
  wire [31:0] _j_T_1 = j + 32'h1; // @[ivncontrol4.scala 118:16]
  wire [3:0] _GEN_264 = _io_ProcessValid_T & j == 32'h8 ? 4'h8 : 4'h0; // @[ivncontrol4.scala 120:77 121:11 129:11]
  wire [31:0] _GEN_265 = _io_ProcessValid_T & j == 32'h8 ? 32'h7 : _GEN_247; // @[ivncontrol4.scala 120:77 122:11]
  wire  _GEN_312 = _io_ProcessValid_T_2; // @[ivncontrol4.scala 153:41]
  wire [31:0] _GEN_313 = rowcount_0 != 32'h0 ? 32'h0 : pin; // @[ivncontrol4.scala 162:30 163:13 37:22]
  wire  _T_27 = rowcount_0 == 32'h0; // @[ivncontrol4.scala 165:23]
  wire [31:0] _GEN_314 = rowcount_0 == 32'h0 & rowcount_1 != 32'h0 ? 32'h1 : _GEN_313; // @[ivncontrol4.scala 165:54 166:13]
  wire  _T_32 = _T_27 & rowcount_1 == 32'h0; // @[ivncontrol4.scala 168:31]
  wire [31:0] _GEN_315 = _T_27 & rowcount_1 == 32'h0 & rowcount_2 != 32'h0 ? 32'h2 : _GEN_314; // @[ivncontrol4.scala 168:77 169:13]
  wire  _T_39 = _T_32 & rowcount_2 == 32'h0; // @[ivncontrol4.scala 171:54]
  wire [31:0] _GEN_316 = _T_32 & rowcount_2 == 32'h0 & rowcount_3 != 32'h0 ? 32'h3 : _GEN_315; // @[ivncontrol4.scala 171:100 172:13]
  wire  _T_48 = _T_39 & rowcount_3 == 32'h0; // @[ivncontrol4.scala 174:77]
  wire [31:0] _GEN_317 = _T_39 & rowcount_3 == 32'h0 & rowcount_4 != 32'h0 ? 32'h4 : _GEN_316; // @[ivncontrol4.scala 174:123 175:13]
  wire  _T_59 = _T_48 & rowcount_4 == 32'h0; // @[ivncontrol4.scala 177:100]
  wire  _T_72 = _T_59 & rowcount_5 == 32'h0; // @[ivncontrol4.scala 180:123]
  wire  valid = _io_ProcessValid_T_2; // @[ivncontrol4.scala 153:41]
  wire [32:0] _T_91 = {{1'd0}, pin}; // @[ivncontrol4.scala 191:27]
  wire [31:0] _GEN_322 = 4'h1 == _T_91[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_323 = 4'h2 == _T_91[3:0] ? rowcount_2 : _GEN_322; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_324 = 4'h3 == _T_91[3:0] ? rowcount_3 : _GEN_323; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_325 = 4'h4 == _T_91[3:0] ? rowcount_4 : _GEN_324; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_326 = 4'h5 == _T_91[3:0] ? rowcount_5 : _GEN_325; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_327 = 4'h6 == _T_91[3:0] ? rowcount_6 : _GEN_326; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_328 = 4'h7 == _T_91[3:0] ? rowcount_7 : _GEN_327; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_329 = 4'h8 == _T_91[3:0] ? rowcount_8 : _GEN_328; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_330 = 4'h9 == _T_91[3:0] ? rowcount_9 : _GEN_329; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_331 = 4'ha == _T_91[3:0] ? rowcount_10 : _GEN_330; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_332 = 4'hb == _T_91[3:0] ? rowcount_11 : _GEN_331; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_333 = 4'hc == _T_91[3:0] ? rowcount_12 : _GEN_332; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_334 = 4'hd == _T_91[3:0] ? rowcount_13 : _GEN_333; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_335 = 4'he == _T_91[3:0] ? rowcount_14 : _GEN_334; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_336 = 4'hf == _T_91[3:0] ? rowcount_15 : _GEN_335; // @[ivncontrol4.scala 191:{35,35}]
  wire [31:0] _GEN_449 = _GEN_336 == 32'h1 ? _T_91[31:0] : 32'h1c; // @[ivncontrol4.scala 142:17 241:50 242:21]
  wire [31:0] _GEN_450 = _GEN_336 == 32'h2 ? _T_91[31:0] : _GEN_449; // @[ivncontrol4.scala 237:51 238:21]
  wire [31:0] _GEN_451 = _GEN_336 == 32'h2 ? _T_91[31:0] : 32'h11; // @[ivncontrol4.scala 142:17 237:51 239:21]
  wire [31:0] _GEN_452 = _GEN_336 == 32'h3 ? _T_91[31:0] : _GEN_450; // @[ivncontrol4.scala 232:50 233:21]
  wire [31:0] _GEN_453 = _GEN_336 == 32'h3 ? _T_91[31:0] : _GEN_451; // @[ivncontrol4.scala 232:50 234:21]
  wire [31:0] _GEN_454 = _GEN_336 == 32'h3 ? _T_91[31:0] : 32'hc; // @[ivncontrol4.scala 142:17 232:50 235:21]
  wire [31:0] _GEN_455 = _GEN_336 == 32'h4 ? _T_91[31:0] : _GEN_452; // @[ivncontrol4.scala 224:50 225:21]
  wire [31:0] _GEN_456 = _GEN_336 == 32'h4 ? _T_91[31:0] : _GEN_453; // @[ivncontrol4.scala 224:50 226:21]
  wire [31:0] _GEN_457 = _GEN_336 == 32'h4 ? _T_91[31:0] : _GEN_454; // @[ivncontrol4.scala 224:50 227:21]
  wire [31:0] _GEN_458 = _GEN_336 == 32'h4 ? _T_91[31:0] : 32'h7; // @[ivncontrol4.scala 142:17 224:50 228:21]
  wire [31:0] _GEN_459 = _GEN_336 == 32'h5 ? _T_91[31:0] : _GEN_455; // @[ivncontrol4.scala 217:50 218:21]
  wire [31:0] _GEN_460 = _GEN_336 == 32'h5 ? _T_91[31:0] : _GEN_456; // @[ivncontrol4.scala 217:50 219:21]
  wire [31:0] _GEN_461 = _GEN_336 == 32'h5 ? _T_91[31:0] : _GEN_457; // @[ivncontrol4.scala 217:50 220:21]
  wire [31:0] _GEN_462 = _GEN_336 == 32'h5 ? _T_91[31:0] : _GEN_458; // @[ivncontrol4.scala 217:50 221:21]
  wire [31:0] _GEN_463 = _GEN_336 == 32'h5 ? _T_91[31:0] : 32'ha; // @[ivncontrol4.scala 143:18 217:50 222:22]
  wire [31:0] _GEN_464 = _GEN_336 == 32'h6 ? _T_91[31:0] : _GEN_459; // @[ivncontrol4.scala 209:52 210:21]
  wire [31:0] _GEN_465 = _GEN_336 == 32'h6 ? _T_91[31:0] : _GEN_460; // @[ivncontrol4.scala 209:52 211:21]
  wire [31:0] _GEN_466 = _GEN_336 == 32'h6 ? _T_91[31:0] : _GEN_461; // @[ivncontrol4.scala 209:52 212:21]
  wire [31:0] _GEN_467 = _GEN_336 == 32'h6 ? _T_91[31:0] : _GEN_462; // @[ivncontrol4.scala 209:52 213:21]
  wire [31:0] _GEN_468 = _GEN_336 == 32'h6 ? _T_91[31:0] : _GEN_463; // @[ivncontrol4.scala 209:52 214:22]
  wire [31:0] _GEN_469 = _GEN_336 == 32'h6 ? _T_91[31:0] : 32'h3; // @[ivncontrol4.scala 143:18 209:52 215:22]
  wire [31:0] _GEN_470 = _GEN_336 == 32'h7 ? _T_91[31:0] : _GEN_464; // @[ivncontrol4.scala 201:52 202:21]
  wire [31:0] _GEN_471 = _GEN_336 == 32'h7 ? _T_91[31:0] : _GEN_465; // @[ivncontrol4.scala 201:52 203:21]
  wire [31:0] _GEN_472 = _GEN_336 == 32'h7 ? _T_91[31:0] : _GEN_466; // @[ivncontrol4.scala 201:52 204:21]
  wire [31:0] _GEN_473 = _GEN_336 == 32'h7 ? _T_91[31:0] : _GEN_467; // @[ivncontrol4.scala 201:52 205:21]
  wire [31:0] _GEN_474 = _GEN_336 == 32'h7 ? _T_91[31:0] : _GEN_468; // @[ivncontrol4.scala 201:52 206:22]
  wire [31:0] _GEN_475 = _GEN_336 == 32'h7 ? _T_91[31:0] : _GEN_469; // @[ivncontrol4.scala 201:52 207:22]
  wire [31:0] _GEN_476 = _GEN_336 == 32'h7 ? _T_91[31:0] : 32'h1b; // @[ivncontrol4.scala 143:18 201:52 208:22]
  wire [31:0] _GEN_477 = _GEN_336 >= 32'h8 ? _T_91[31:0] : _GEN_470; // @[ivncontrol4.scala 191:42 192:21]
  wire [31:0] _GEN_478 = _GEN_336 >= 32'h8 ? _T_91[31:0] : _GEN_471; // @[ivncontrol4.scala 191:42 193:21]
  wire [31:0] _GEN_479 = _GEN_336 >= 32'h8 ? _T_91[31:0] : _GEN_472; // @[ivncontrol4.scala 191:42 194:21]
  wire [31:0] _GEN_480 = _GEN_336 >= 32'h8 ? _T_91[31:0] : _GEN_473; // @[ivncontrol4.scala 191:42 195:21]
  wire [31:0] _GEN_481 = _GEN_336 >= 32'h8 ? _T_91[31:0] : _GEN_474; // @[ivncontrol4.scala 191:42 196:22]
  wire [31:0] _GEN_482 = _GEN_336 >= 32'h8 ? _T_91[31:0] : _GEN_475; // @[ivncontrol4.scala 191:42 197:22]
  wire [31:0] _GEN_483 = _GEN_336 >= 32'h8 ? _T_91[31:0] : _GEN_476; // @[ivncontrol4.scala 191:42 198:22]
  wire [31:0] _GEN_484 = _GEN_336 >= 32'h8 ? _T_91[31:0] : 32'h15; // @[ivncontrol4.scala 143:18 191:42 199:22]
  wire [31:0] _T_127 = 32'h8 - _GEN_336; // @[ivncontrol4.scala 245:18]
  wire [31:0] _i_vn_1_T_15 = 32'h1 + pin; // @[ivncontrol4.scala 246:29]
  wire [31:0] _GEN_597 = _T_127 == 32'h1 ? _i_vn_1_T_15 : _GEN_484; // @[ivncontrol4.scala 286:54 289:22]
  wire [31:0] _GEN_598 = _T_127 == 32'h2 ? _i_vn_1_T_15 : _GEN_483; // @[ivncontrol4.scala 281:54 284:22]
  wire [31:0] _GEN_599 = _T_127 == 32'h2 ? _i_vn_1_T_15 : _GEN_597; // @[ivncontrol4.scala 281:54 285:22]
  wire [31:0] _GEN_600 = _T_127 == 32'h3 ? _i_vn_1_T_15 : _GEN_482; // @[ivncontrol4.scala 274:54 276:22]
  wire [31:0] _GEN_601 = _T_127 == 32'h3 ? _i_vn_1_T_15 : _GEN_598; // @[ivncontrol4.scala 274:54 277:22]
  wire [31:0] _GEN_602 = _T_127 == 32'h3 ? _i_vn_1_T_15 : _GEN_599; // @[ivncontrol4.scala 274:54 278:22]
  wire [31:0] _GEN_603 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_481; // @[ivncontrol4.scala 268:54 270:22]
  wire [31:0] _GEN_604 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_600; // @[ivncontrol4.scala 268:54 271:22]
  wire [31:0] _GEN_605 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_601; // @[ivncontrol4.scala 268:54 272:22]
  wire [31:0] _GEN_606 = _T_127 == 32'h4 ? _i_vn_1_T_15 : _GEN_602; // @[ivncontrol4.scala 268:54 273:22]
  wire [31:0] _GEN_607 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_480; // @[ivncontrol4.scala 261:54 263:21]
  wire [31:0] _GEN_608 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_603; // @[ivncontrol4.scala 261:54 264:22]
  wire [31:0] _GEN_609 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_604; // @[ivncontrol4.scala 261:54 265:22]
  wire [31:0] _GEN_610 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_605; // @[ivncontrol4.scala 261:54 266:22]
  wire [31:0] _GEN_611 = _T_127 == 32'h5 ? _i_vn_1_T_15 : _GEN_606; // @[ivncontrol4.scala 261:54 267:22]
  wire [31:0] _GEN_612 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_479; // @[ivncontrol4.scala 254:54 255:22]
  wire [31:0] _GEN_613 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_607; // @[ivncontrol4.scala 254:54 256:21]
  wire [31:0] _GEN_614 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_608; // @[ivncontrol4.scala 254:54 257:22]
  wire [31:0] _GEN_615 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_609; // @[ivncontrol4.scala 254:54 258:22]
  wire [31:0] _GEN_616 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_610; // @[ivncontrol4.scala 254:54 259:22]
  wire [31:0] _GEN_617 = _T_127 == 32'h6 ? _i_vn_1_T_15 : _GEN_611; // @[ivncontrol4.scala 254:54 260:22]
  wire [31:0] _GEN_618 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_478; // @[ivncontrol4.scala 245:49 246:22]
  wire [31:0] _GEN_619 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_612; // @[ivncontrol4.scala 245:49 247:21]
  wire [31:0] _GEN_620 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_613; // @[ivncontrol4.scala 245:49 248:21]
  wire [31:0] _GEN_621 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_614; // @[ivncontrol4.scala 245:49 249:22]
  wire [31:0] _GEN_622 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_615; // @[ivncontrol4.scala 245:49 250:22]
  wire [31:0] _GEN_623 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_616; // @[ivncontrol4.scala 245:49 251:22]
  wire [31:0] _GEN_624 = _T_127 == 32'h7 ? _i_vn_1_T_15 : _GEN_617; // @[ivncontrol4.scala 245:49 252:22]
  wire [31:0] _GEN_642 = 4'h1 == _i_vn_1_T_15[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_643 = 4'h2 == _i_vn_1_T_15[3:0] ? rowcount_2 : _GEN_642; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_644 = 4'h3 == _i_vn_1_T_15[3:0] ? rowcount_3 : _GEN_643; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_645 = 4'h4 == _i_vn_1_T_15[3:0] ? rowcount_4 : _GEN_644; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_646 = 4'h5 == _i_vn_1_T_15[3:0] ? rowcount_5 : _GEN_645; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_647 = 4'h6 == _i_vn_1_T_15[3:0] ? rowcount_6 : _GEN_646; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_648 = 4'h7 == _i_vn_1_T_15[3:0] ? rowcount_7 : _GEN_647; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_649 = 4'h8 == _i_vn_1_T_15[3:0] ? rowcount_8 : _GEN_648; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_650 = 4'h9 == _i_vn_1_T_15[3:0] ? rowcount_9 : _GEN_649; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_651 = 4'ha == _i_vn_1_T_15[3:0] ? rowcount_10 : _GEN_650; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_652 = 4'hb == _i_vn_1_T_15[3:0] ? rowcount_11 : _GEN_651; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_653 = 4'hc == _i_vn_1_T_15[3:0] ? rowcount_12 : _GEN_652; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_654 = 4'hd == _i_vn_1_T_15[3:0] ? rowcount_13 : _GEN_653; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_655 = 4'he == _i_vn_1_T_15[3:0] ? rowcount_14 : _GEN_654; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _GEN_656 = 4'hf == _i_vn_1_T_15[3:0] ? rowcount_15 : _GEN_655; // @[ivncontrol4.scala 292:{41,41}]
  wire [31:0] _T_172 = _GEN_336 + _GEN_656; // @[ivncontrol4.scala 292:41]
  wire [31:0] _T_174 = 32'h8 - _T_172; // @[ivncontrol4.scala 292:18]
  wire [31:0] _i_vn_1_T_17 = 32'h2 + pin; // @[ivncontrol4.scala 293:29]
  wire [31:0] _GEN_849 = _T_174 == 32'h1 ? _i_vn_1_T_17 : _GEN_624; // @[ivncontrol4.scala 335:78 338:22]
  wire [31:0] _GEN_850 = _T_174 == 32'h2 ? _i_vn_1_T_17 : _GEN_623; // @[ivncontrol4.scala 329:76 332:22]
  wire [31:0] _GEN_851 = _T_174 == 32'h2 ? _i_vn_1_T_17 : _GEN_849; // @[ivncontrol4.scala 329:76 333:22]
  wire [31:0] _GEN_852 = _T_174 == 32'h3 ? _i_vn_1_T_17 : _GEN_622; // @[ivncontrol4.scala 322:78 324:23]
  wire [31:0] _GEN_853 = _T_174 == 32'h3 ? _i_vn_1_T_17 : _GEN_850; // @[ivncontrol4.scala 322:78 325:22]
  wire [31:0] _GEN_854 = _T_174 == 32'h3 ? _i_vn_1_T_17 : _GEN_851; // @[ivncontrol4.scala 322:78 326:22]
  wire [31:0] _GEN_855 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_621; // @[ivncontrol4.scala 316:78 318:22]
  wire [31:0] _GEN_856 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_852; // @[ivncontrol4.scala 316:78 319:22]
  wire [31:0] _GEN_857 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_853; // @[ivncontrol4.scala 316:78 320:22]
  wire [31:0] _GEN_858 = _T_174 == 32'h4 ? _i_vn_1_T_17 : _GEN_854; // @[ivncontrol4.scala 316:78 321:22]
  wire [31:0] _GEN_859 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_620; // @[ivncontrol4.scala 309:76 311:23]
  wire [31:0] _GEN_860 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_855; // @[ivncontrol4.scala 309:76 312:22]
  wire [31:0] _GEN_861 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_856; // @[ivncontrol4.scala 309:76 313:22]
  wire [31:0] _GEN_862 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_857; // @[ivncontrol4.scala 309:76 314:22]
  wire [31:0] _GEN_863 = _T_174 == 32'h5 ? _i_vn_1_T_17 : _GEN_858; // @[ivncontrol4.scala 309:76 315:22]
  wire [31:0] _GEN_864 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_619; // @[ivncontrol4.scala 301:77 303:22]
  wire [31:0] _GEN_865 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_859; // @[ivncontrol4.scala 301:77 304:21]
  wire [31:0] _GEN_866 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_860; // @[ivncontrol4.scala 301:77 305:22]
  wire [31:0] _GEN_867 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_861; // @[ivncontrol4.scala 301:77 306:22]
  wire [31:0] _GEN_868 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_862; // @[ivncontrol4.scala 301:77 307:22]
  wire [31:0] _GEN_869 = _T_174 == 32'h6 ? _i_vn_1_T_17 : _GEN_863; // @[ivncontrol4.scala 301:77 308:22]
  wire [31:0] _GEN_870 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_618; // @[ivncontrol4.scala 292:73 293:22]
  wire [31:0] _GEN_871 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_864; // @[ivncontrol4.scala 292:73 294:21]
  wire [31:0] _GEN_872 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_865; // @[ivncontrol4.scala 292:73 295:21]
  wire [31:0] _GEN_873 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_866; // @[ivncontrol4.scala 292:73 296:22]
  wire [31:0] _GEN_874 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_867; // @[ivncontrol4.scala 292:73 297:22]
  wire [31:0] _GEN_875 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_868; // @[ivncontrol4.scala 292:73 298:22]
  wire [31:0] _GEN_876 = _T_174 == 32'h7 ? _i_vn_1_T_17 : _GEN_869; // @[ivncontrol4.scala 292:73 299:22]
  wire [31:0] _GEN_910 = 4'h1 == _i_vn_1_T_17[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_911 = 4'h2 == _i_vn_1_T_17[3:0] ? rowcount_2 : _GEN_910; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_912 = 4'h3 == _i_vn_1_T_17[3:0] ? rowcount_3 : _GEN_911; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_913 = 4'h4 == _i_vn_1_T_17[3:0] ? rowcount_4 : _GEN_912; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_914 = 4'h5 == _i_vn_1_T_17[3:0] ? rowcount_5 : _GEN_913; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_915 = 4'h6 == _i_vn_1_T_17[3:0] ? rowcount_6 : _GEN_914; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_916 = 4'h7 == _i_vn_1_T_17[3:0] ? rowcount_7 : _GEN_915; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_917 = 4'h8 == _i_vn_1_T_17[3:0] ? rowcount_8 : _GEN_916; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_918 = 4'h9 == _i_vn_1_T_17[3:0] ? rowcount_9 : _GEN_917; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_919 = 4'ha == _i_vn_1_T_17[3:0] ? rowcount_10 : _GEN_918; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_920 = 4'hb == _i_vn_1_T_17[3:0] ? rowcount_11 : _GEN_919; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_921 = 4'hc == _i_vn_1_T_17[3:0] ? rowcount_12 : _GEN_920; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_922 = 4'hd == _i_vn_1_T_17[3:0] ? rowcount_13 : _GEN_921; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_923 = 4'he == _i_vn_1_T_17[3:0] ? rowcount_14 : _GEN_922; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _GEN_924 = 4'hf == _i_vn_1_T_17[3:0] ? rowcount_15 : _GEN_923; // @[ivncontrol4.scala 343:{62,62}]
  wire [31:0] _T_254 = _T_172 + _GEN_924; // @[ivncontrol4.scala 343:62]
  wire [31:0] _T_256 = 32'h8 - _T_254; // @[ivncontrol4.scala 343:17]
  wire [31:0] _i_vn_1_T_19 = 32'h3 + pin; // @[ivncontrol4.scala 344:29]
  wire [31:0] _GEN_1213 = _T_256 == 32'h1 ? _i_vn_1_T_19 : _GEN_876; // @[ivncontrol4.scala 386:100 389:22]
  wire [31:0] _GEN_1214 = _T_256 == 32'h2 ? _i_vn_1_T_19 : _GEN_875; // @[ivncontrol4.scala 380:98 383:22]
  wire [31:0] _GEN_1215 = _T_256 == 32'h2 ? _i_vn_1_T_19 : _GEN_1213; // @[ivncontrol4.scala 380:98 384:22]
  wire [31:0] _GEN_1216 = _T_256 == 32'h3 ? _i_vn_1_T_19 : _GEN_874; // @[ivncontrol4.scala 373:100 375:23]
  wire [31:0] _GEN_1217 = _T_256 == 32'h3 ? _i_vn_1_T_19 : _GEN_1214; // @[ivncontrol4.scala 373:100 376:22]
  wire [31:0] _GEN_1218 = _T_256 == 32'h3 ? _i_vn_1_T_19 : _GEN_1215; // @[ivncontrol4.scala 373:100 377:22]
  wire [31:0] _GEN_1219 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_873; // @[ivncontrol4.scala 367:100 369:22]
  wire [31:0] _GEN_1220 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_1216; // @[ivncontrol4.scala 367:100 370:22]
  wire [31:0] _GEN_1221 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_1217; // @[ivncontrol4.scala 367:100 371:22]
  wire [31:0] _GEN_1222 = _T_256 == 32'h4 ? _i_vn_1_T_19 : _GEN_1218; // @[ivncontrol4.scala 367:100 372:22]
  wire [31:0] _GEN_1223 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_872; // @[ivncontrol4.scala 360:98 362:23]
  wire [31:0] _GEN_1224 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1219; // @[ivncontrol4.scala 360:98 363:22]
  wire [31:0] _GEN_1225 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1220; // @[ivncontrol4.scala 360:98 364:22]
  wire [31:0] _GEN_1226 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1221; // @[ivncontrol4.scala 360:98 365:22]
  wire [31:0] _GEN_1227 = _T_256 == 32'h5 ? _i_vn_1_T_19 : _GEN_1222; // @[ivncontrol4.scala 360:98 366:22]
  wire [31:0] _GEN_1228 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_871; // @[ivncontrol4.scala 352:99 354:22]
  wire [31:0] _GEN_1229 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1223; // @[ivncontrol4.scala 352:99 355:21]
  wire [31:0] _GEN_1230 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1224; // @[ivncontrol4.scala 352:99 356:22]
  wire [31:0] _GEN_1231 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1225; // @[ivncontrol4.scala 352:99 357:22]
  wire [31:0] _GEN_1232 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1226; // @[ivncontrol4.scala 352:99 358:22]
  wire [31:0] _GEN_1233 = _T_256 == 32'h6 ? _i_vn_1_T_19 : _GEN_1227; // @[ivncontrol4.scala 352:99 359:22]
  wire [31:0] _GEN_1234 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_870; // @[ivncontrol4.scala 343:94 344:22]
  wire [31:0] _GEN_1235 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1228; // @[ivncontrol4.scala 343:94 345:21]
  wire [31:0] _GEN_1236 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1229; // @[ivncontrol4.scala 343:94 346:21]
  wire [31:0] _GEN_1237 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1230; // @[ivncontrol4.scala 343:94 347:22]
  wire [31:0] _GEN_1238 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1231; // @[ivncontrol4.scala 343:94 348:22]
  wire [31:0] _GEN_1239 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1232; // @[ivncontrol4.scala 343:94 349:22]
  wire [31:0] _GEN_1240 = _T_256 == 32'h7 ? _i_vn_1_T_19 : _GEN_1233; // @[ivncontrol4.scala 343:94 350:22]
  wire [31:0] _GEN_1290 = 4'h1 == _i_vn_1_T_19[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1291 = 4'h2 == _i_vn_1_T_19[3:0] ? rowcount_2 : _GEN_1290; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1292 = 4'h3 == _i_vn_1_T_19[3:0] ? rowcount_3 : _GEN_1291; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1293 = 4'h4 == _i_vn_1_T_19[3:0] ? rowcount_4 : _GEN_1292; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1294 = 4'h5 == _i_vn_1_T_19[3:0] ? rowcount_5 : _GEN_1293; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1295 = 4'h6 == _i_vn_1_T_19[3:0] ? rowcount_6 : _GEN_1294; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1296 = 4'h7 == _i_vn_1_T_19[3:0] ? rowcount_7 : _GEN_1295; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1297 = 4'h8 == _i_vn_1_T_19[3:0] ? rowcount_8 : _GEN_1296; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1298 = 4'h9 == _i_vn_1_T_19[3:0] ? rowcount_9 : _GEN_1297; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1299 = 4'ha == _i_vn_1_T_19[3:0] ? rowcount_10 : _GEN_1298; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1300 = 4'hb == _i_vn_1_T_19[3:0] ? rowcount_11 : _GEN_1299; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1301 = 4'hc == _i_vn_1_T_19[3:0] ? rowcount_12 : _GEN_1300; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1302 = 4'hd == _i_vn_1_T_19[3:0] ? rowcount_13 : _GEN_1301; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1303 = 4'he == _i_vn_1_T_19[3:0] ? rowcount_14 : _GEN_1302; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _GEN_1304 = 4'hf == _i_vn_1_T_19[3:0] ? rowcount_15 : _GEN_1303; // @[ivncontrol4.scala 393:{86,86}]
  wire [31:0] _T_371 = _T_254 + _GEN_1304; // @[ivncontrol4.scala 393:86]
  wire [31:0] _T_373 = 32'h8 - _T_371; // @[ivncontrol4.scala 393:19]
  wire [31:0] _i_vn_1_T_21 = 32'h4 + pin; // @[ivncontrol4.scala 394:29]
  wire [31:0] _GEN_1689 = _T_373 == 32'h1 ? _i_vn_1_T_21 : _GEN_1240; // @[ivncontrol4.scala 436:122 439:22]
  wire [31:0] _GEN_1690 = _T_373 == 32'h2 ? _i_vn_1_T_21 : _GEN_1239; // @[ivncontrol4.scala 430:121 433:22]
  wire [31:0] _GEN_1691 = _T_373 == 32'h2 ? _i_vn_1_T_21 : _GEN_1689; // @[ivncontrol4.scala 430:121 434:22]
  wire [31:0] _GEN_1692 = _T_373 == 32'h3 ? _i_vn_1_T_21 : _GEN_1238; // @[ivncontrol4.scala 423:123 425:23]
  wire [31:0] _GEN_1693 = _T_373 == 32'h3 ? _i_vn_1_T_21 : _GEN_1690; // @[ivncontrol4.scala 423:123 426:22]
  wire [31:0] _GEN_1694 = _T_373 == 32'h3 ? _i_vn_1_T_21 : _GEN_1691; // @[ivncontrol4.scala 423:123 427:22]
  wire [31:0] _GEN_1695 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1237; // @[ivncontrol4.scala 417:122 419:22]
  wire [31:0] _GEN_1696 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1692; // @[ivncontrol4.scala 417:122 420:22]
  wire [31:0] _GEN_1697 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1693; // @[ivncontrol4.scala 417:122 421:22]
  wire [31:0] _GEN_1698 = _T_373 == 32'h4 ? _i_vn_1_T_21 : _GEN_1694; // @[ivncontrol4.scala 417:122 422:22]
  wire [31:0] _GEN_1699 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1236; // @[ivncontrol4.scala 410:121 412:23]
  wire [31:0] _GEN_1700 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1695; // @[ivncontrol4.scala 410:121 413:22]
  wire [31:0] _GEN_1701 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1696; // @[ivncontrol4.scala 410:121 414:22]
  wire [31:0] _GEN_1702 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1697; // @[ivncontrol4.scala 410:121 415:22]
  wire [31:0] _GEN_1703 = _T_373 == 32'h5 ? _i_vn_1_T_21 : _GEN_1698; // @[ivncontrol4.scala 410:121 416:22]
  wire [31:0] _GEN_1704 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1235; // @[ivncontrol4.scala 402:121 404:22]
  wire [31:0] _GEN_1705 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1699; // @[ivncontrol4.scala 402:121 405:21]
  wire [31:0] _GEN_1706 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1700; // @[ivncontrol4.scala 402:121 406:22]
  wire [31:0] _GEN_1707 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1701; // @[ivncontrol4.scala 402:121 407:22]
  wire [31:0] _GEN_1708 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1702; // @[ivncontrol4.scala 402:121 408:22]
  wire [31:0] _GEN_1709 = _T_373 == 32'h6 ? _i_vn_1_T_21 : _GEN_1703; // @[ivncontrol4.scala 402:121 409:22]
  wire [31:0] _GEN_1710 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1234; // @[ivncontrol4.scala 393:118 394:22]
  wire [31:0] _GEN_1711 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1704; // @[ivncontrol4.scala 393:118 395:21]
  wire [31:0] _GEN_1712 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1705; // @[ivncontrol4.scala 393:118 396:21]
  wire [31:0] _GEN_1713 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1706; // @[ivncontrol4.scala 393:118 397:22]
  wire [31:0] _GEN_1714 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1707; // @[ivncontrol4.scala 393:118 398:22]
  wire [31:0] _GEN_1715 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1708; // @[ivncontrol4.scala 393:118 399:22]
  wire [31:0] _GEN_1716 = _T_373 == 32'h7 ? _i_vn_1_T_21 : _GEN_1709; // @[ivncontrol4.scala 393:118 400:22]
  wire [31:0] _GEN_1782 = 4'h1 == _i_vn_1_T_21[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1783 = 4'h2 == _i_vn_1_T_21[3:0] ? rowcount_2 : _GEN_1782; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1784 = 4'h3 == _i_vn_1_T_21[3:0] ? rowcount_3 : _GEN_1783; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1785 = 4'h4 == _i_vn_1_T_21[3:0] ? rowcount_4 : _GEN_1784; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1786 = 4'h5 == _i_vn_1_T_21[3:0] ? rowcount_5 : _GEN_1785; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1787 = 4'h6 == _i_vn_1_T_21[3:0] ? rowcount_6 : _GEN_1786; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1788 = 4'h7 == _i_vn_1_T_21[3:0] ? rowcount_7 : _GEN_1787; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1789 = 4'h8 == _i_vn_1_T_21[3:0] ? rowcount_8 : _GEN_1788; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1790 = 4'h9 == _i_vn_1_T_21[3:0] ? rowcount_9 : _GEN_1789; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1791 = 4'ha == _i_vn_1_T_21[3:0] ? rowcount_10 : _GEN_1790; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1792 = 4'hb == _i_vn_1_T_21[3:0] ? rowcount_11 : _GEN_1791; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1793 = 4'hc == _i_vn_1_T_21[3:0] ? rowcount_12 : _GEN_1792; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1794 = 4'hd == _i_vn_1_T_21[3:0] ? rowcount_13 : _GEN_1793; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1795 = 4'he == _i_vn_1_T_21[3:0] ? rowcount_14 : _GEN_1794; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _GEN_1796 = 4'hf == _i_vn_1_T_21[3:0] ? rowcount_15 : _GEN_1795; // @[ivncontrol4.scala 443:{108,108}]
  wire [31:0] _T_523 = _T_371 + _GEN_1796; // @[ivncontrol4.scala 443:108]
  wire [31:0] _T_525 = 32'h8 - _T_523; // @[ivncontrol4.scala 443:19]
  wire [31:0] _i_vn_1_T_23 = 32'h5 + pin; // @[ivncontrol4.scala 444:29]
  wire [31:0] _GEN_2277 = _T_525 == 32'h1 ? _i_vn_1_T_23 : _GEN_1716; // @[ivncontrol4.scala 486:144 489:22]
  wire [31:0] _GEN_2278 = _T_525 == 32'h2 ? _i_vn_1_T_23 : _GEN_1715; // @[ivncontrol4.scala 480:143 483:22]
  wire [31:0] _GEN_2279 = _T_525 == 32'h2 ? _i_vn_1_T_23 : _GEN_2277; // @[ivncontrol4.scala 480:143 484:22]
  wire [31:0] _GEN_2280 = _T_525 == 32'h3 ? _i_vn_1_T_23 : _GEN_1714; // @[ivncontrol4.scala 473:145 475:23]
  wire [31:0] _GEN_2281 = _T_525 == 32'h3 ? _i_vn_1_T_23 : _GEN_2278; // @[ivncontrol4.scala 473:145 476:22]
  wire [31:0] _GEN_2282 = _T_525 == 32'h3 ? _i_vn_1_T_23 : _GEN_2279; // @[ivncontrol4.scala 473:145 477:22]
  wire [31:0] _GEN_2283 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_1713; // @[ivncontrol4.scala 467:143 469:22]
  wire [31:0] _GEN_2284 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_2280; // @[ivncontrol4.scala 467:143 470:22]
  wire [31:0] _GEN_2285 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_2281; // @[ivncontrol4.scala 467:143 471:22]
  wire [31:0] _GEN_2286 = _T_525 == 32'h4 ? _i_vn_1_T_23 : _GEN_2282; // @[ivncontrol4.scala 467:143 472:22]
  wire [31:0] _GEN_2287 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_1712; // @[ivncontrol4.scala 460:143 462:23]
  wire [31:0] _GEN_2288 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2283; // @[ivncontrol4.scala 460:143 463:22]
  wire [31:0] _GEN_2289 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2284; // @[ivncontrol4.scala 460:143 464:22]
  wire [31:0] _GEN_2290 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2285; // @[ivncontrol4.scala 460:143 465:22]
  wire [31:0] _GEN_2291 = _T_525 == 32'h5 ? _i_vn_1_T_23 : _GEN_2286; // @[ivncontrol4.scala 460:143 466:22]
  wire [31:0] _GEN_2292 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_1711; // @[ivncontrol4.scala 452:143 454:22]
  wire [31:0] _GEN_2293 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2287; // @[ivncontrol4.scala 452:143 455:21]
  wire [31:0] _GEN_2294 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2288; // @[ivncontrol4.scala 452:143 456:22]
  wire [31:0] _GEN_2295 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2289; // @[ivncontrol4.scala 452:143 457:22]
  wire [31:0] _GEN_2296 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2290; // @[ivncontrol4.scala 452:143 458:22]
  wire [31:0] _GEN_2297 = _T_525 == 32'h6 ? _i_vn_1_T_23 : _GEN_2291; // @[ivncontrol4.scala 452:143 459:22]
  wire [31:0] _GEN_2298 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_1710; // @[ivncontrol4.scala 443:140 444:22]
  wire [31:0] _GEN_2299 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2292; // @[ivncontrol4.scala 443:140 445:21]
  wire [31:0] _GEN_2300 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2293; // @[ivncontrol4.scala 443:140 446:21]
  wire [31:0] _GEN_2301 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2294; // @[ivncontrol4.scala 443:140 447:22]
  wire [31:0] _GEN_2302 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2295; // @[ivncontrol4.scala 443:140 448:22]
  wire [31:0] _GEN_2303 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2296; // @[ivncontrol4.scala 443:140 449:22]
  wire [31:0] _GEN_2304 = _T_525 == 32'h7 ? _i_vn_1_T_23 : _GEN_2297; // @[ivncontrol4.scala 443:140 450:22]
  wire [31:0] _GEN_2386 = 4'h1 == _i_vn_1_T_23[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2387 = 4'h2 == _i_vn_1_T_23[3:0] ? rowcount_2 : _GEN_2386; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2388 = 4'h3 == _i_vn_1_T_23[3:0] ? rowcount_3 : _GEN_2387; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2389 = 4'h4 == _i_vn_1_T_23[3:0] ? rowcount_4 : _GEN_2388; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2390 = 4'h5 == _i_vn_1_T_23[3:0] ? rowcount_5 : _GEN_2389; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2391 = 4'h6 == _i_vn_1_T_23[3:0] ? rowcount_6 : _GEN_2390; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2392 = 4'h7 == _i_vn_1_T_23[3:0] ? rowcount_7 : _GEN_2391; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2393 = 4'h8 == _i_vn_1_T_23[3:0] ? rowcount_8 : _GEN_2392; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2394 = 4'h9 == _i_vn_1_T_23[3:0] ? rowcount_9 : _GEN_2393; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2395 = 4'ha == _i_vn_1_T_23[3:0] ? rowcount_10 : _GEN_2394; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2396 = 4'hb == _i_vn_1_T_23[3:0] ? rowcount_11 : _GEN_2395; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2397 = 4'hc == _i_vn_1_T_23[3:0] ? rowcount_12 : _GEN_2396; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2398 = 4'hd == _i_vn_1_T_23[3:0] ? rowcount_13 : _GEN_2397; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2399 = 4'he == _i_vn_1_T_23[3:0] ? rowcount_14 : _GEN_2398; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _GEN_2400 = 4'hf == _i_vn_1_T_23[3:0] ? rowcount_15 : _GEN_2399; // @[ivncontrol4.scala 494:{130,130}]
  wire [31:0] _T_710 = _T_523 + _GEN_2400; // @[ivncontrol4.scala 494:130]
  wire [31:0] _T_712 = 32'h8 - _T_710; // @[ivncontrol4.scala 494:19]
  wire [31:0] _i_vn_1_T_25 = 32'h6 + pin; // @[ivncontrol4.scala 495:29]
  wire [31:0] _GEN_2977 = _T_712 == 32'h1 ? _i_vn_1_T_25 : _GEN_2304; // @[ivncontrol4.scala 537:166 540:22]
  wire [31:0] _GEN_2978 = _T_712 == 32'h2 ? _i_vn_1_T_25 : _GEN_2303; // @[ivncontrol4.scala 531:166 534:22]
  wire [31:0] _GEN_2979 = _T_712 == 32'h2 ? _i_vn_1_T_25 : _GEN_2977; // @[ivncontrol4.scala 531:166 535:22]
  wire [31:0] _GEN_2980 = _T_712 == 32'h3 ? _i_vn_1_T_25 : _GEN_2302; // @[ivncontrol4.scala 524:168 526:23]
  wire [31:0] _GEN_2981 = _T_712 == 32'h3 ? _i_vn_1_T_25 : _GEN_2978; // @[ivncontrol4.scala 524:168 527:22]
  wire [31:0] _GEN_2982 = _T_712 == 32'h3 ? _i_vn_1_T_25 : _GEN_2979; // @[ivncontrol4.scala 524:168 528:22]
  wire [31:0] _GEN_2983 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2301; // @[ivncontrol4.scala 518:166 520:22]
  wire [31:0] _GEN_2984 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2980; // @[ivncontrol4.scala 518:166 521:22]
  wire [31:0] _GEN_2985 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2981; // @[ivncontrol4.scala 518:166 522:22]
  wire [31:0] _GEN_2986 = _T_712 == 32'h4 ? _i_vn_1_T_25 : _GEN_2982; // @[ivncontrol4.scala 518:166 523:22]
  wire [31:0] _GEN_2987 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2300; // @[ivncontrol4.scala 511:166 513:23]
  wire [31:0] _GEN_2988 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2983; // @[ivncontrol4.scala 511:166 514:22]
  wire [31:0] _GEN_2989 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2984; // @[ivncontrol4.scala 511:166 515:22]
  wire [31:0] _GEN_2990 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2985; // @[ivncontrol4.scala 511:166 516:22]
  wire [31:0] _GEN_2991 = _T_712 == 32'h5 ? _i_vn_1_T_25 : _GEN_2986; // @[ivncontrol4.scala 511:166 517:22]
  wire [31:0] _GEN_2992 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2299; // @[ivncontrol4.scala 503:166 505:22]
  wire [31:0] _GEN_2993 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2987; // @[ivncontrol4.scala 503:166 506:21]
  wire [31:0] _GEN_2994 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2988; // @[ivncontrol4.scala 503:166 507:22]
  wire [31:0] _GEN_2995 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2989; // @[ivncontrol4.scala 503:166 508:22]
  wire [31:0] _GEN_2996 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2990; // @[ivncontrol4.scala 503:166 509:22]
  wire [31:0] _GEN_2997 = _T_712 == 32'h6 ? _i_vn_1_T_25 : _GEN_2991; // @[ivncontrol4.scala 503:166 510:22]
  wire [31:0] _GEN_2998 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2298; // @[ivncontrol4.scala 494:162 495:22]
  wire [31:0] _GEN_2999 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2992; // @[ivncontrol4.scala 494:162 496:21]
  wire [31:0] _GEN_3000 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2993; // @[ivncontrol4.scala 494:162 497:21]
  wire [31:0] _GEN_3001 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2994; // @[ivncontrol4.scala 494:162 498:22]
  wire [31:0] _GEN_3002 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2995; // @[ivncontrol4.scala 494:162 499:22]
  wire [31:0] _GEN_3003 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2996; // @[ivncontrol4.scala 494:162 500:22]
  wire [31:0] _GEN_3004 = _T_712 == 32'h7 ? _i_vn_1_T_25 : _GEN_2997; // @[ivncontrol4.scala 494:162 501:22]
  wire [31:0] _GEN_3102 = 4'h1 == _i_vn_1_T_25[3:0] ? rowcount_1 : rowcount_0; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3103 = 4'h2 == _i_vn_1_T_25[3:0] ? rowcount_2 : _GEN_3102; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3104 = 4'h3 == _i_vn_1_T_25[3:0] ? rowcount_3 : _GEN_3103; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3105 = 4'h4 == _i_vn_1_T_25[3:0] ? rowcount_4 : _GEN_3104; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3106 = 4'h5 == _i_vn_1_T_25[3:0] ? rowcount_5 : _GEN_3105; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3107 = 4'h6 == _i_vn_1_T_25[3:0] ? rowcount_6 : _GEN_3106; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3108 = 4'h7 == _i_vn_1_T_25[3:0] ? rowcount_7 : _GEN_3107; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3109 = 4'h8 == _i_vn_1_T_25[3:0] ? rowcount_8 : _GEN_3108; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3110 = 4'h9 == _i_vn_1_T_25[3:0] ? rowcount_9 : _GEN_3109; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3111 = 4'ha == _i_vn_1_T_25[3:0] ? rowcount_10 : _GEN_3110; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3112 = 4'hb == _i_vn_1_T_25[3:0] ? rowcount_11 : _GEN_3111; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3113 = 4'hc == _i_vn_1_T_25[3:0] ? rowcount_12 : _GEN_3112; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3114 = 4'hd == _i_vn_1_T_25[3:0] ? rowcount_13 : _GEN_3113; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3115 = 4'he == _i_vn_1_T_25[3:0] ? rowcount_14 : _GEN_3114; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _GEN_3116 = 4'hf == _i_vn_1_T_25[3:0] ? rowcount_15 : _GEN_3115; // @[ivncontrol4.scala 545:{152,152}]
  wire [31:0] _T_932 = _T_710 + _GEN_3116; // @[ivncontrol4.scala 545:152]
  wire [31:0] _T_934 = 32'h8 - _T_932; // @[ivncontrol4.scala 545:19]
  wire [31:0] _i_vn_1_T_27 = 32'h7 + pin; // @[ivncontrol4.scala 546:29]
  wire [31:0] _GEN_3789 = _T_934 == 32'h1 ? _i_vn_1_T_27 : _GEN_3004; // @[ivncontrol4.scala 588:188 591:22]
  wire [31:0] _GEN_3790 = _T_934 == 32'h2 ? _i_vn_1_T_27 : _GEN_3003; // @[ivncontrol4.scala 582:188 585:22]
  wire [31:0] _GEN_3791 = _T_934 == 32'h2 ? _i_vn_1_T_27 : _GEN_3789; // @[ivncontrol4.scala 582:188 586:22]
  wire [31:0] _GEN_3792 = _T_934 == 32'h3 ? _i_vn_1_T_27 : _GEN_3002; // @[ivncontrol4.scala 575:190 577:23]
  wire [31:0] _GEN_3793 = _T_934 == 32'h3 ? _i_vn_1_T_27 : _GEN_3790; // @[ivncontrol4.scala 575:190 578:22]
  wire [31:0] _GEN_3794 = _T_934 == 32'h3 ? _i_vn_1_T_27 : _GEN_3791; // @[ivncontrol4.scala 575:190 579:22]
  wire [31:0] _GEN_3795 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_3001; // @[ivncontrol4.scala 569:188 571:22]
  wire [31:0] _GEN_3796 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_3792; // @[ivncontrol4.scala 569:188 572:22]
  wire [31:0] _GEN_3797 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_3793; // @[ivncontrol4.scala 569:188 573:22]
  wire [31:0] _GEN_3798 = _T_934 == 32'h4 ? _i_vn_1_T_27 : _GEN_3794; // @[ivncontrol4.scala 569:188 574:22]
  wire [31:0] _GEN_3799 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3000; // @[ivncontrol4.scala 562:188 564:23]
  wire [31:0] _GEN_3800 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3795; // @[ivncontrol4.scala 562:188 565:22]
  wire [31:0] _GEN_3801 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3796; // @[ivncontrol4.scala 562:188 566:22]
  wire [31:0] _GEN_3802 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3797; // @[ivncontrol4.scala 562:188 567:22]
  wire [31:0] _GEN_3803 = _T_934 == 32'h5 ? _i_vn_1_T_27 : _GEN_3798; // @[ivncontrol4.scala 562:188 568:22]
  wire [31:0] _GEN_3804 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_2999; // @[ivncontrol4.scala 554:188 556:22]
  wire [31:0] _GEN_3805 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3799; // @[ivncontrol4.scala 554:188 557:21]
  wire [31:0] _GEN_3806 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3800; // @[ivncontrol4.scala 554:188 558:22]
  wire [31:0] _GEN_3807 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3801; // @[ivncontrol4.scala 554:188 559:22]
  wire [31:0] _GEN_3808 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3802; // @[ivncontrol4.scala 554:188 560:22]
  wire [31:0] _GEN_3809 = _T_934 == 32'h6 ? _i_vn_1_T_27 : _GEN_3803; // @[ivncontrol4.scala 554:188 561:22]
  wire [31:0] _GEN_3810 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_2998; // @[ivncontrol4.scala 545:184 546:22]
  wire [31:0] _GEN_3811 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3804; // @[ivncontrol4.scala 545:184 547:21]
  wire [31:0] _GEN_3812 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3805; // @[ivncontrol4.scala 545:184 548:21]
  wire [31:0] _GEN_3813 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3806; // @[ivncontrol4.scala 545:184 549:22]
  wire [31:0] _GEN_3814 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3807; // @[ivncontrol4.scala 545:184 550:22]
  wire [31:0] _GEN_3815 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3808; // @[ivncontrol4.scala 545:184 551:22]
  wire [31:0] _GEN_3816 = _T_934 == 32'h7 ? _i_vn_1_T_27 : _GEN_3809; // @[ivncontrol4.scala 545:184 552:22]
  wire [31:0] _GEN_3817 = _GEN_312 ? _GEN_477 : 32'h1c; // @[ivncontrol4.scala 142:17 189:28]
  wire [31:0] _GEN_3818 = _GEN_312 ? _GEN_3810 : 32'h11; // @[ivncontrol4.scala 142:17 189:28]
  wire [31:0] _GEN_3819 = _GEN_312 ? _GEN_3811 : 32'hc; // @[ivncontrol4.scala 142:17 189:28]
  wire [31:0] _GEN_3820 = _GEN_312 ? _GEN_3812 : 32'h7; // @[ivncontrol4.scala 142:17 189:28]
  wire [31:0] _GEN_3821 = _GEN_312 ? _GEN_3813 : 32'ha; // @[ivncontrol4.scala 143:18 189:28]
  wire [31:0] _GEN_3822 = _GEN_312 ? _GEN_3814 : 32'h3; // @[ivncontrol4.scala 143:18 189:28]
  wire [31:0] _GEN_3823 = _GEN_312 ? _GEN_3815 : 32'h1b; // @[ivncontrol4.scala 143:18 189:28]
  wire [31:0] _GEN_3824 = _GEN_312 ? _GEN_3816 : 32'h15; // @[ivncontrol4.scala 143:18 189:28]
  wire  valid1 = 1'h0;
  wire [31:0] _GEN_4221 = reset ? 32'h0 : _GEN_3817; // @[ivncontrol4.scala 17:{23,23}]
  wire [31:0] _GEN_4222 = reset ? 32'h0 : _GEN_3818; // @[ivncontrol4.scala 17:{23,23}]
  wire [31:0] _GEN_4223 = reset ? 32'h0 : _GEN_3819; // @[ivncontrol4.scala 17:{23,23}]
  wire [31:0] _GEN_4224 = reset ? 32'h0 : _GEN_3820; // @[ivncontrol4.scala 17:{23,23}]
  wire [31:0] _GEN_4225 = reset ? 32'h0 : _GEN_3821; // @[ivncontrol4.scala 18:{24,24}]
  wire [31:0] _GEN_4226 = reset ? 32'h0 : _GEN_3822; // @[ivncontrol4.scala 18:{24,24}]
  wire [31:0] _GEN_4227 = reset ? 32'h0 : _GEN_3823; // @[ivncontrol4.scala 18:{24,24}]
  wire [31:0] _GEN_4228 = reset ? 32'h0 : _GEN_3824; // @[ivncontrol4.scala 18:{24,24}]
  assign io_o_vn_0 = i_vn_0; // @[ivncontrol4.scala 138:13]
  assign io_o_vn_1 = i_vn_1; // @[ivncontrol4.scala 138:13]
  assign io_o_vn_2 = i_vn_2; // @[ivncontrol4.scala 138:13]
  assign io_o_vn_3 = i_vn_3; // @[ivncontrol4.scala 138:13]
  assign io_o_vn2_0 = i_vn2_0; // @[ivncontrol4.scala 139:14]
  assign io_o_vn2_1 = i_vn2_1; // @[ivncontrol4.scala 139:14]
  assign io_o_vn2_2 = i_vn2_2; // @[ivncontrol4.scala 139:14]
  assign io_o_vn2_3 = i_vn2_3; // @[ivncontrol4.scala 139:14]
  always @(posedge clock) begin
    i_vn_0 <= _GEN_4221[4:0]; // @[ivncontrol4.scala 17:{23,23}]
    i_vn_1 <= _GEN_4222[4:0]; // @[ivncontrol4.scala 17:{23,23}]
    i_vn_2 <= _GEN_4223[4:0]; // @[ivncontrol4.scala 17:{23,23}]
    i_vn_3 <= _GEN_4224[4:0]; // @[ivncontrol4.scala 17:{23,23}]
    i_vn2_0 <= _GEN_4225[4:0]; // @[ivncontrol4.scala 18:{24,24}]
    i_vn2_1 <= _GEN_4226[4:0]; // @[ivncontrol4.scala 18:{24,24}]
    i_vn2_2 <= _GEN_4227[4:0]; // @[ivncontrol4.scala 18:{24,24}]
    i_vn2_3 <= _GEN_4228[4:0]; // @[ivncontrol4.scala 18:{24,24}]
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_0 <= io_Stationary_matrix_0_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_1 <= io_Stationary_matrix_0_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_2 <= io_Stationary_matrix_0_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_3 <= io_Stationary_matrix_0_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_4 <= io_Stationary_matrix_0_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_5 <= io_Stationary_matrix_0_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_6 <= io_Stationary_matrix_0_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_0_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_0_7 <= io_Stationary_matrix_0_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_0 <= io_Stationary_matrix_1_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_1 <= io_Stationary_matrix_1_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_2 <= io_Stationary_matrix_1_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_3 <= io_Stationary_matrix_1_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_4 <= io_Stationary_matrix_1_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_5 <= io_Stationary_matrix_1_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_6 <= io_Stationary_matrix_1_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_1_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_1_7 <= io_Stationary_matrix_1_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_0 <= io_Stationary_matrix_2_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_1 <= io_Stationary_matrix_2_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_2 <= io_Stationary_matrix_2_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_3 <= io_Stationary_matrix_2_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_4 <= io_Stationary_matrix_2_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_5 <= io_Stationary_matrix_2_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_6 <= io_Stationary_matrix_2_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_2_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_2_7 <= io_Stationary_matrix_2_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_0 <= io_Stationary_matrix_3_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_1 <= io_Stationary_matrix_3_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_2 <= io_Stationary_matrix_3_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_3 <= io_Stationary_matrix_3_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_4 <= io_Stationary_matrix_3_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_5 <= io_Stationary_matrix_3_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_6 <= io_Stationary_matrix_3_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_3_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_3_7 <= io_Stationary_matrix_3_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_0 <= io_Stationary_matrix_4_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_1 <= io_Stationary_matrix_4_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_2 <= io_Stationary_matrix_4_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_3 <= io_Stationary_matrix_4_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_4 <= io_Stationary_matrix_4_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_5 <= io_Stationary_matrix_4_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_6 <= io_Stationary_matrix_4_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_4_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_4_7 <= io_Stationary_matrix_4_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_0 <= io_Stationary_matrix_5_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_1 <= io_Stationary_matrix_5_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_2 <= io_Stationary_matrix_5_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_3 <= io_Stationary_matrix_5_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_4 <= io_Stationary_matrix_5_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_5 <= io_Stationary_matrix_5_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_6 <= io_Stationary_matrix_5_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_5_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_5_7 <= io_Stationary_matrix_5_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_0 <= io_Stationary_matrix_6_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_1 <= io_Stationary_matrix_6_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_2 <= io_Stationary_matrix_6_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_3 <= io_Stationary_matrix_6_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_4 <= io_Stationary_matrix_6_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_5 <= io_Stationary_matrix_6_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_6 <= io_Stationary_matrix_6_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_6_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_6_7 <= io_Stationary_matrix_6_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_0 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_0 <= io_Stationary_matrix_7_0; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_1 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_1 <= io_Stationary_matrix_7_1; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_2 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_2 <= io_Stationary_matrix_7_2; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_3 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_3 <= io_Stationary_matrix_7_3; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_4 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_4 <= io_Stationary_matrix_7_4; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_5 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_5 <= io_Stationary_matrix_7_5; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_6 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_6 <= io_Stationary_matrix_7_6; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 21:27]
      solution_7_7 <= 16'h0; // @[ivncontrol4.scala 21:27]
    end else begin
      solution_7_7 <= io_Stationary_matrix_7_7; // @[ivncontrol4.scala 24:28]
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_0 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_0 <= count_0; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_1 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_1 <= count_1; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_2 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_2 <= count_2; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_3 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_3 <= count_3; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_4 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_4 <= count_4; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_5 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_5 <= count_5; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_6 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_6 <= count_6; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_7 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_7 <= count_7; // @[ivncontrol4.scala 85:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_8 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_8 <= 32'h0; // @[ivncontrol4.scala 87:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_9 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_9 <= 32'h0; // @[ivncontrol4.scala 87:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_10 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_10 <= 32'h0; // @[ivncontrol4.scala 87:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_11 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_11 <= 32'h0; // @[ivncontrol4.scala 87:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_12 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_12 <= 32'h0; // @[ivncontrol4.scala 87:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_13 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_13 <= 32'h0; // @[ivncontrol4.scala 87:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_14 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 78:75]
        rowcount_14 <= 32'h0; // @[ivncontrol4.scala 87:19]
      end
    end
    if (reset) begin // @[ivncontrol4.scala 27:27]
      rowcount_15 <= 32'h0; // @[ivncontrol4.scala 27:27]
    end
    if (reset) begin // @[ivncontrol4.scala 37:22]
      pin <= 32'h0; // @[ivncontrol4.scala 37:22]
    end else if (_T_72 & rowcount_6 == 32'h0 & rowcount_7 != 32'h0) begin // @[ivncontrol4.scala 183:192]
      pin <= 32'h7; // @[ivncontrol4.scala 184:13]
    end else if (_T_59 & rowcount_5 == 32'h0 & rowcount_6 != 32'h0) begin // @[ivncontrol4.scala 180:169]
      pin <= 32'h6; // @[ivncontrol4.scala 181:13]
    end else if (_T_48 & rowcount_4 == 32'h0 & rowcount_5 != 32'h0) begin // @[ivncontrol4.scala 177:146]
      pin <= 32'h5; // @[ivncontrol4.scala 178:13]
    end else begin
      pin <= _GEN_317;
    end
    if (reset) begin // @[ivncontrol4.scala 41:20]
      i <= 32'h0; // @[ivncontrol4.scala 41:20]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
        i <= _GEN_247;
      end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
        i <= _GEN_247;
      end else begin
        i <= _GEN_265;
      end
    end
    if (reset) begin // @[ivncontrol4.scala 42:20]
      j <= 32'h0; // @[ivncontrol4.scala 42:20]
    end else if (io_validpin) begin // @[ivncontrol4.scala 46:29]
      if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
        j <= 32'h8; // @[ivncontrol4.scala 116:11]
      end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
        j <= _j_T_1; // @[ivncontrol4.scala 118:11]
      end else begin
        j <= {{28'd0}, _GEN_264};
      end
    end
    if (3'h0 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h0 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h0 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h0 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h0 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h0 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h0 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h0 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_0_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h1 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_1_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h2 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_2_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h3 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_3_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h4 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_4_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h5 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_5_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h6 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_6_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h0 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_0 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h1 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_1 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h2 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_2 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h3 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_3 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h4 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_4 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h5 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_5 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h6 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_6 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (3'h7 == i[2:0] & 3'h7 == j[2:0]) begin // @[ivncontrol4.scala 63:17]
      mat_7_7 <= _mat_T_1_T_2; // @[ivncontrol4.scala 63:17]
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_0 <= _GEN_224;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_0 <= _GEN_224;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h0 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_0 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_0 <= _GEN_224;
      end
    end else begin
      count_0 <= _GEN_224;
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_1 <= _GEN_225;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_1 <= _GEN_225;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h1 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_1 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_1 <= _GEN_225;
      end
    end else begin
      count_1 <= _GEN_225;
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_2 <= _GEN_226;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_2 <= _GEN_226;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h2 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_2 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_2 <= _GEN_226;
      end
    end else begin
      count_2 <= _GEN_226;
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_3 <= _GEN_227;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_3 <= _GEN_227;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h3 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_3 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_3 <= _GEN_227;
      end
    end else begin
      count_3 <= _GEN_227;
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_4 <= _GEN_228;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_4 <= _GEN_228;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h4 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_4 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_4 <= _GEN_228;
      end
    end else begin
      count_4 <= _GEN_228;
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_5 <= _GEN_229;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_5 <= _GEN_229;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h5 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_5 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_5 <= _GEN_229;
      end
    end else begin
      count_5 <= _GEN_229;
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_6 <= _GEN_230;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_6 <= _GEN_230;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h6 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_6 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_6 <= _GEN_230;
      end
    end else begin
      count_6 <= _GEN_230;
    end
    if (_io_ProcessValid_T_2) begin // @[ivncontrol4.scala 115:77]
      count_7 <= _GEN_231;
    end else if (j < 32'h7 & i <= 32'h7) begin // @[ivncontrol4.scala 117:77]
      count_7 <= _GEN_231;
    end else if (_io_ProcessValid_T & j == 32'h8) begin // @[ivncontrol4.scala 120:77]
      if (3'h7 == i[2:0]) begin // @[ivncontrol4.scala 123:18]
        count_7 <= _GEN_207; // @[ivncontrol4.scala 123:18]
      end else begin
        count_7 <= _GEN_231;
      end
    end else begin
      count_7 <= _GEN_231;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  i_vn_0 = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  i_vn_1 = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  i_vn_2 = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  i_vn_3 = _RAND_3[4:0];
  _RAND_4 = {1{`RANDOM}};
  i_vn2_0 = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  i_vn2_1 = _RAND_5[4:0];
  _RAND_6 = {1{`RANDOM}};
  i_vn2_2 = _RAND_6[4:0];
  _RAND_7 = {1{`RANDOM}};
  i_vn2_3 = _RAND_7[4:0];
  _RAND_8 = {1{`RANDOM}};
  solution_0_0 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  solution_0_1 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  solution_0_2 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  solution_0_3 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  solution_0_4 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  solution_0_5 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  solution_0_6 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  solution_0_7 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  solution_1_0 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  solution_1_1 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  solution_1_2 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  solution_1_3 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  solution_1_4 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  solution_1_5 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  solution_1_6 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  solution_1_7 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  solution_2_0 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  solution_2_1 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  solution_2_2 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  solution_2_3 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  solution_2_4 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  solution_2_5 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  solution_2_6 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  solution_2_7 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  solution_3_0 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  solution_3_1 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  solution_3_2 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  solution_3_3 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  solution_3_4 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  solution_3_5 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  solution_3_6 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  solution_3_7 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  solution_4_0 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  solution_4_1 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  solution_4_2 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  solution_4_3 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  solution_4_4 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  solution_4_5 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  solution_4_6 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  solution_4_7 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  solution_5_0 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  solution_5_1 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  solution_5_2 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  solution_5_3 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  solution_5_4 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  solution_5_5 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  solution_5_6 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  solution_5_7 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  solution_6_0 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  solution_6_1 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  solution_6_2 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  solution_6_3 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  solution_6_4 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  solution_6_5 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  solution_6_6 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  solution_6_7 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  solution_7_0 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  solution_7_1 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  solution_7_2 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  solution_7_3 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  solution_7_4 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  solution_7_5 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  solution_7_6 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  solution_7_7 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  rowcount_0 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  rowcount_1 = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  rowcount_2 = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  rowcount_3 = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  rowcount_4 = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  rowcount_5 = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  rowcount_6 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  rowcount_7 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  rowcount_8 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  rowcount_9 = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  rowcount_10 = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  rowcount_11 = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  rowcount_12 = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  rowcount_13 = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  rowcount_14 = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  rowcount_15 = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  pin = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  i = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  j = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  mat_0_0 = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  mat_0_1 = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  mat_0_2 = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  mat_0_3 = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  mat_0_4 = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  mat_0_5 = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  mat_0_6 = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  mat_0_7 = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  mat_1_0 = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  mat_1_1 = _RAND_100[31:0];
  _RAND_101 = {1{`RANDOM}};
  mat_1_2 = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  mat_1_3 = _RAND_102[31:0];
  _RAND_103 = {1{`RANDOM}};
  mat_1_4 = _RAND_103[31:0];
  _RAND_104 = {1{`RANDOM}};
  mat_1_5 = _RAND_104[31:0];
  _RAND_105 = {1{`RANDOM}};
  mat_1_6 = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  mat_1_7 = _RAND_106[31:0];
  _RAND_107 = {1{`RANDOM}};
  mat_2_0 = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  mat_2_1 = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  mat_2_2 = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  mat_2_3 = _RAND_110[31:0];
  _RAND_111 = {1{`RANDOM}};
  mat_2_4 = _RAND_111[31:0];
  _RAND_112 = {1{`RANDOM}};
  mat_2_5 = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  mat_2_6 = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  mat_2_7 = _RAND_114[31:0];
  _RAND_115 = {1{`RANDOM}};
  mat_3_0 = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  mat_3_1 = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  mat_3_2 = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  mat_3_3 = _RAND_118[31:0];
  _RAND_119 = {1{`RANDOM}};
  mat_3_4 = _RAND_119[31:0];
  _RAND_120 = {1{`RANDOM}};
  mat_3_5 = _RAND_120[31:0];
  _RAND_121 = {1{`RANDOM}};
  mat_3_6 = _RAND_121[31:0];
  _RAND_122 = {1{`RANDOM}};
  mat_3_7 = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  mat_4_0 = _RAND_123[31:0];
  _RAND_124 = {1{`RANDOM}};
  mat_4_1 = _RAND_124[31:0];
  _RAND_125 = {1{`RANDOM}};
  mat_4_2 = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  mat_4_3 = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  mat_4_4 = _RAND_127[31:0];
  _RAND_128 = {1{`RANDOM}};
  mat_4_5 = _RAND_128[31:0];
  _RAND_129 = {1{`RANDOM}};
  mat_4_6 = _RAND_129[31:0];
  _RAND_130 = {1{`RANDOM}};
  mat_4_7 = _RAND_130[31:0];
  _RAND_131 = {1{`RANDOM}};
  mat_5_0 = _RAND_131[31:0];
  _RAND_132 = {1{`RANDOM}};
  mat_5_1 = _RAND_132[31:0];
  _RAND_133 = {1{`RANDOM}};
  mat_5_2 = _RAND_133[31:0];
  _RAND_134 = {1{`RANDOM}};
  mat_5_3 = _RAND_134[31:0];
  _RAND_135 = {1{`RANDOM}};
  mat_5_4 = _RAND_135[31:0];
  _RAND_136 = {1{`RANDOM}};
  mat_5_5 = _RAND_136[31:0];
  _RAND_137 = {1{`RANDOM}};
  mat_5_6 = _RAND_137[31:0];
  _RAND_138 = {1{`RANDOM}};
  mat_5_7 = _RAND_138[31:0];
  _RAND_139 = {1{`RANDOM}};
  mat_6_0 = _RAND_139[31:0];
  _RAND_140 = {1{`RANDOM}};
  mat_6_1 = _RAND_140[31:0];
  _RAND_141 = {1{`RANDOM}};
  mat_6_2 = _RAND_141[31:0];
  _RAND_142 = {1{`RANDOM}};
  mat_6_3 = _RAND_142[31:0];
  _RAND_143 = {1{`RANDOM}};
  mat_6_4 = _RAND_143[31:0];
  _RAND_144 = {1{`RANDOM}};
  mat_6_5 = _RAND_144[31:0];
  _RAND_145 = {1{`RANDOM}};
  mat_6_6 = _RAND_145[31:0];
  _RAND_146 = {1{`RANDOM}};
  mat_6_7 = _RAND_146[31:0];
  _RAND_147 = {1{`RANDOM}};
  mat_7_0 = _RAND_147[31:0];
  _RAND_148 = {1{`RANDOM}};
  mat_7_1 = _RAND_148[31:0];
  _RAND_149 = {1{`RANDOM}};
  mat_7_2 = _RAND_149[31:0];
  _RAND_150 = {1{`RANDOM}};
  mat_7_3 = _RAND_150[31:0];
  _RAND_151 = {1{`RANDOM}};
  mat_7_4 = _RAND_151[31:0];
  _RAND_152 = {1{`RANDOM}};
  mat_7_5 = _RAND_152[31:0];
  _RAND_153 = {1{`RANDOM}};
  mat_7_6 = _RAND_153[31:0];
  _RAND_154 = {1{`RANDOM}};
  mat_7_7 = _RAND_154[31:0];
  _RAND_155 = {1{`RANDOM}};
  count_0 = _RAND_155[31:0];
  _RAND_156 = {1{`RANDOM}};
  count_1 = _RAND_156[31:0];
  _RAND_157 = {1{`RANDOM}};
  count_2 = _RAND_157[31:0];
  _RAND_158 = {1{`RANDOM}};
  count_3 = _RAND_158[31:0];
  _RAND_159 = {1{`RANDOM}};
  count_4 = _RAND_159[31:0];
  _RAND_160 = {1{`RANDOM}};
  count_5 = _RAND_160[31:0];
  _RAND_161 = {1{`RANDOM}};
  count_6 = _RAND_161[31:0];
  _RAND_162 = {1{`RANDOM}};
  count_7 = _RAND_162[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ivntop(
  input         clock,
  input         reset,
  output        io_ProcessValid,
  input  [15:0] io_Stationary_matrix_0_0,
  input  [15:0] io_Stationary_matrix_0_1,
  input  [15:0] io_Stationary_matrix_0_2,
  input  [15:0] io_Stationary_matrix_0_3,
  input  [15:0] io_Stationary_matrix_0_4,
  input  [15:0] io_Stationary_matrix_0_5,
  input  [15:0] io_Stationary_matrix_0_6,
  input  [15:0] io_Stationary_matrix_0_7,
  input  [15:0] io_Stationary_matrix_1_0,
  input  [15:0] io_Stationary_matrix_1_1,
  input  [15:0] io_Stationary_matrix_1_2,
  input  [15:0] io_Stationary_matrix_1_3,
  input  [15:0] io_Stationary_matrix_1_4,
  input  [15:0] io_Stationary_matrix_1_5,
  input  [15:0] io_Stationary_matrix_1_6,
  input  [15:0] io_Stationary_matrix_1_7,
  input  [15:0] io_Stationary_matrix_2_0,
  input  [15:0] io_Stationary_matrix_2_1,
  input  [15:0] io_Stationary_matrix_2_2,
  input  [15:0] io_Stationary_matrix_2_3,
  input  [15:0] io_Stationary_matrix_2_4,
  input  [15:0] io_Stationary_matrix_2_5,
  input  [15:0] io_Stationary_matrix_2_6,
  input  [15:0] io_Stationary_matrix_2_7,
  input  [15:0] io_Stationary_matrix_3_0,
  input  [15:0] io_Stationary_matrix_3_1,
  input  [15:0] io_Stationary_matrix_3_2,
  input  [15:0] io_Stationary_matrix_3_3,
  input  [15:0] io_Stationary_matrix_3_4,
  input  [15:0] io_Stationary_matrix_3_5,
  input  [15:0] io_Stationary_matrix_3_6,
  input  [15:0] io_Stationary_matrix_3_7,
  input  [15:0] io_Stationary_matrix_4_0,
  input  [15:0] io_Stationary_matrix_4_1,
  input  [15:0] io_Stationary_matrix_4_2,
  input  [15:0] io_Stationary_matrix_4_3,
  input  [15:0] io_Stationary_matrix_4_4,
  input  [15:0] io_Stationary_matrix_4_5,
  input  [15:0] io_Stationary_matrix_4_6,
  input  [15:0] io_Stationary_matrix_4_7,
  input  [15:0] io_Stationary_matrix_5_0,
  input  [15:0] io_Stationary_matrix_5_1,
  input  [15:0] io_Stationary_matrix_5_2,
  input  [15:0] io_Stationary_matrix_5_3,
  input  [15:0] io_Stationary_matrix_5_4,
  input  [15:0] io_Stationary_matrix_5_5,
  input  [15:0] io_Stationary_matrix_5_6,
  input  [15:0] io_Stationary_matrix_5_7,
  input  [15:0] io_Stationary_matrix_6_0,
  input  [15:0] io_Stationary_matrix_6_1,
  input  [15:0] io_Stationary_matrix_6_2,
  input  [15:0] io_Stationary_matrix_6_3,
  input  [15:0] io_Stationary_matrix_6_4,
  input  [15:0] io_Stationary_matrix_6_5,
  input  [15:0] io_Stationary_matrix_6_6,
  input  [15:0] io_Stationary_matrix_6_7,
  input  [15:0] io_Stationary_matrix_7_0,
  input  [15:0] io_Stationary_matrix_7_1,
  input  [15:0] io_Stationary_matrix_7_2,
  input  [15:0] io_Stationary_matrix_7_3,
  input  [15:0] io_Stationary_matrix_7_4,
  input  [15:0] io_Stationary_matrix_7_5,
  input  [15:0] io_Stationary_matrix_7_6,
  input  [15:0] io_Stationary_matrix_7_7,
  output [4:0]  io_o_vn_0_0,
  output [4:0]  io_o_vn_0_1,
  output [4:0]  io_o_vn_0_2,
  output [4:0]  io_o_vn_0_3,
  output [4:0]  io_o_vn_1_0,
  output [4:0]  io_o_vn_1_1,
  output [4:0]  io_o_vn_1_2,
  output [4:0]  io_o_vn_1_3,
  output [4:0]  io_o_vn_2_0,
  output [4:0]  io_o_vn_2_1,
  output [4:0]  io_o_vn_2_2,
  output [4:0]  io_o_vn_2_3,
  output [4:0]  io_o_vn_3_0,
  output [4:0]  io_o_vn_3_1,
  output [4:0]  io_o_vn_3_2,
  output [4:0]  io_o_vn_3_3,
  output [4:0]  io_o_vn_4_0,
  output [4:0]  io_o_vn_4_1,
  output [4:0]  io_o_vn_4_2,
  output [4:0]  io_o_vn_4_3,
  output [4:0]  io_o_vn_5_0,
  output [4:0]  io_o_vn_5_1,
  output [4:0]  io_o_vn_5_2,
  output [4:0]  io_o_vn_5_3,
  output [4:0]  io_o_vn_6_0,
  output [4:0]  io_o_vn_6_1,
  output [4:0]  io_o_vn_6_2,
  output [4:0]  io_o_vn_6_3,
  output [4:0]  io_o_vn_7_0,
  output [4:0]  io_o_vn_7_1,
  output [4:0]  io_o_vn_7_2,
  output [4:0]  io_o_vn_7_3,
  output [4:0]  io_o_vn_8_0,
  output [4:0]  io_o_vn_8_1,
  output [4:0]  io_o_vn_8_2,
  output [4:0]  io_o_vn_8_3,
  output [4:0]  io_o_vn_9_0,
  output [4:0]  io_o_vn_9_1,
  output [4:0]  io_o_vn_9_2,
  output [4:0]  io_o_vn_9_3,
  output [4:0]  io_o_vn_10_0,
  output [4:0]  io_o_vn_10_1,
  output [4:0]  io_o_vn_10_2,
  output [4:0]  io_o_vn_10_3,
  output [4:0]  io_o_vn_11_0,
  output [4:0]  io_o_vn_11_1,
  output [4:0]  io_o_vn_11_2,
  output [4:0]  io_o_vn_11_3,
  output [4:0]  io_o_vn_12_0,
  output [4:0]  io_o_vn_12_1,
  output [4:0]  io_o_vn_12_2,
  output [4:0]  io_o_vn_12_3,
  output [4:0]  io_o_vn_13_0,
  output [4:0]  io_o_vn_13_1,
  output [4:0]  io_o_vn_13_2,
  output [4:0]  io_o_vn_13_3,
  output [4:0]  io_o_vn_14_0,
  output [4:0]  io_o_vn_14_1,
  output [4:0]  io_o_vn_14_2,
  output [4:0]  io_o_vn_14_3,
  output [4:0]  io_o_vn_15_0,
  output [4:0]  io_o_vn_15_1,
  output [4:0]  io_o_vn_15_2,
  output [4:0]  io_o_vn_15_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
`endif // RANDOMIZE_REG_INIT
  wire  my_stationary_clock; // @[ivntop.scala 29:31]
  wire  my_stationary_reset; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_0_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_0_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_0_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_0_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_0_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_0_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_0_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_0_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_1_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_1_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_1_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_1_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_1_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_1_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_1_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_1_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_2_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_2_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_2_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_2_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_2_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_2_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_2_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_2_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_3_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_3_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_3_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_3_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_3_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_3_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_3_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_3_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_4_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_4_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_4_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_4_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_4_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_4_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_4_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_4_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_5_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_5_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_5_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_5_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_5_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_5_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_5_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_5_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_6_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_6_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_6_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_6_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_6_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_6_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_6_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_6_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_7_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_7_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_7_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_7_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_7_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_7_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_7_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_Stationary_matrix_7_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_0_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_0_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_0_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_0_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_0_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_0_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_0_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_0_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_1_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_1_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_1_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_1_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_1_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_1_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_1_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_1_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_2_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_2_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_2_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_2_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_2_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_2_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_2_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_2_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_3_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_3_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_3_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_3_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_3_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_3_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_3_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_3_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_4_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_4_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_4_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_4_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_4_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_4_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_4_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_4_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_5_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_5_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_5_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_5_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_5_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_5_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_5_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_5_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_6_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_6_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_6_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_6_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_6_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_6_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_6_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_6_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_7_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_7_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_7_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_7_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_7_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_7_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_7_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix1_7_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_0_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_0_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_0_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_0_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_0_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_0_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_0_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_0_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_1_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_1_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_1_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_1_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_1_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_1_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_1_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_1_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_2_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_2_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_2_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_2_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_2_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_2_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_2_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_2_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_3_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_3_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_3_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_3_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_3_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_3_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_3_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_3_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_4_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_4_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_4_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_4_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_4_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_4_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_4_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_4_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_5_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_5_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_5_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_5_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_5_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_5_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_5_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_5_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_6_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_6_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_6_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_6_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_6_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_6_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_6_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_6_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_7_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_7_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_7_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_7_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_7_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_7_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_7_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix2_7_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_0_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_0_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_0_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_0_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_0_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_0_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_0_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_0_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_1_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_1_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_1_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_1_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_1_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_1_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_1_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_1_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_2_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_2_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_2_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_2_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_2_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_2_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_2_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_2_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_3_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_3_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_3_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_3_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_3_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_3_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_3_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_3_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_4_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_4_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_4_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_4_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_4_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_4_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_4_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_4_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_5_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_5_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_5_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_5_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_5_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_5_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_5_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_5_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_6_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_6_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_6_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_6_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_6_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_6_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_6_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_6_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_7_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_7_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_7_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_7_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_7_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_7_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_7_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix3_7_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_0_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_0_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_0_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_0_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_0_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_0_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_0_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_0_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_1_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_1_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_1_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_1_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_1_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_1_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_1_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_1_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_2_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_2_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_2_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_2_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_2_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_2_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_2_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_2_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_3_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_3_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_3_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_3_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_3_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_3_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_3_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_3_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_4_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_4_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_4_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_4_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_4_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_4_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_4_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_4_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_5_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_5_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_5_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_5_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_5_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_5_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_5_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_5_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_6_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_6_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_6_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_6_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_6_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_6_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_6_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_6_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_7_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_7_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_7_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_7_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_7_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_7_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_7_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix4_7_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_0_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_0_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_0_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_0_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_0_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_0_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_0_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_0_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_1_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_1_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_1_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_1_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_1_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_1_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_1_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_1_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_2_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_2_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_2_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_2_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_2_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_2_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_2_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_2_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_3_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_3_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_3_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_3_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_3_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_3_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_3_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_3_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_4_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_4_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_4_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_4_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_4_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_4_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_4_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_4_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_5_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_5_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_5_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_5_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_5_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_5_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_5_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_5_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_6_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_6_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_6_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_6_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_6_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_6_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_6_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_6_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_7_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_7_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_7_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_7_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_7_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_7_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_7_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix5_7_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_0_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_0_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_0_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_0_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_0_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_0_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_0_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_0_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_1_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_1_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_1_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_1_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_1_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_1_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_1_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_1_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_2_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_2_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_2_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_2_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_2_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_2_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_2_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_2_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_3_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_3_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_3_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_3_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_3_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_3_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_3_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_3_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_4_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_4_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_4_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_4_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_4_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_4_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_4_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_4_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_5_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_5_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_5_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_5_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_5_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_5_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_5_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_5_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_6_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_6_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_6_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_6_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_6_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_6_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_6_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_6_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_7_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_7_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_7_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_7_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_7_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_7_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_7_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix6_7_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_0_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_0_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_0_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_0_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_0_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_0_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_0_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_0_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_1_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_1_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_1_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_1_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_1_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_1_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_1_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_1_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_2_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_2_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_2_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_2_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_2_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_2_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_2_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_2_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_3_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_3_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_3_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_3_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_3_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_3_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_3_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_3_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_4_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_4_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_4_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_4_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_4_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_4_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_4_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_4_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_5_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_5_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_5_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_5_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_5_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_5_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_5_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_5_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_6_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_6_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_6_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_6_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_6_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_6_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_6_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_6_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_7_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_7_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_7_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_7_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_7_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_7_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_7_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix7_7_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_0_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_0_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_0_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_0_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_0_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_0_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_0_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_0_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_1_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_1_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_1_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_1_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_1_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_1_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_1_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_1_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_2_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_2_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_2_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_2_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_2_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_2_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_2_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_2_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_3_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_3_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_3_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_3_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_3_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_3_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_3_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_3_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_4_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_4_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_4_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_4_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_4_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_4_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_4_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_4_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_5_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_5_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_5_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_5_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_5_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_5_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_5_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_5_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_6_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_6_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_6_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_6_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_6_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_6_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_6_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_6_7; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_7_0; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_7_1; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_7_2; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_7_3; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_7_4; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_7_5; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_7_6; // @[ivntop.scala 29:31]
  wire [15:0] my_stationary_io_o_Stationary_matrix8_7_7; // @[ivntop.scala 29:31]
  wire  my_ivn1_clock; // @[ivntop.scala 69:24]
  wire  my_ivn1_reset; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_0_0; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_0_1; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_0_2; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_0_3; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_0_4; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_0_5; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_0_6; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_0_7; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_1_0; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_1_1; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_1_2; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_1_3; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_1_4; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_1_5; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_1_6; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_1_7; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_2_0; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_2_1; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_2_2; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_2_3; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_2_4; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_2_5; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_2_6; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_2_7; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_3_0; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_3_1; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_3_2; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_3_3; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_3_4; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_3_5; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_3_6; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_3_7; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_4_0; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_4_1; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_4_2; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_4_3; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_4_4; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_4_5; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_4_6; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_4_7; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_5_0; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_5_1; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_5_2; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_5_3; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_5_4; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_5_5; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_5_6; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_5_7; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_6_0; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_6_1; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_6_2; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_6_3; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_6_4; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_6_5; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_6_6; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_6_7; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_7_0; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_7_1; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_7_2; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_7_3; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_7_4; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_7_5; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_7_6; // @[ivntop.scala 69:24]
  wire [15:0] my_ivn1_io_Stationary_matrix_7_7; // @[ivntop.scala 69:24]
  wire [4:0] my_ivn1_io_o_vn_0; // @[ivntop.scala 69:24]
  wire [4:0] my_ivn1_io_o_vn_1; // @[ivntop.scala 69:24]
  wire [4:0] my_ivn1_io_o_vn_2; // @[ivntop.scala 69:24]
  wire [4:0] my_ivn1_io_o_vn_3; // @[ivntop.scala 69:24]
  wire [4:0] my_ivn1_io_o_vn2_0; // @[ivntop.scala 69:24]
  wire [4:0] my_ivn1_io_o_vn2_1; // @[ivntop.scala 69:24]
  wire [4:0] my_ivn1_io_o_vn2_2; // @[ivntop.scala 69:24]
  wire [4:0] my_ivn1_io_o_vn2_3; // @[ivntop.scala 69:24]
  wire  my_ivn1_io_ProcessValid; // @[ivntop.scala 69:24]
  wire  my_ivn1_io_validpin; // @[ivntop.scala 69:24]
  wire  my_ivn2_clock; // @[ivntop.scala 78:24]
  wire  my_ivn2_reset; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_0_0; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_0_1; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_0_2; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_0_3; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_0_4; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_0_5; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_0_6; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_0_7; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_1_0; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_1_1; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_1_2; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_1_3; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_1_4; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_1_5; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_1_6; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_1_7; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_2_0; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_2_1; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_2_2; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_2_3; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_2_4; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_2_5; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_2_6; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_2_7; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_3_0; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_3_1; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_3_2; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_3_3; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_3_4; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_3_5; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_3_6; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_3_7; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_4_0; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_4_1; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_4_2; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_4_3; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_4_4; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_4_5; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_4_6; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_4_7; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_5_0; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_5_1; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_5_2; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_5_3; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_5_4; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_5_5; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_5_6; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_5_7; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_6_0; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_6_1; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_6_2; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_6_3; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_6_4; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_6_5; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_6_6; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_6_7; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_7_0; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_7_1; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_7_2; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_7_3; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_7_4; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_7_5; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_7_6; // @[ivntop.scala 78:24]
  wire [15:0] my_ivn2_io_Stationary_matrix_7_7; // @[ivntop.scala 78:24]
  wire [4:0] my_ivn2_io_o_vn_0; // @[ivntop.scala 78:24]
  wire [4:0] my_ivn2_io_o_vn_1; // @[ivntop.scala 78:24]
  wire [4:0] my_ivn2_io_o_vn_2; // @[ivntop.scala 78:24]
  wire [4:0] my_ivn2_io_o_vn_3; // @[ivntop.scala 78:24]
  wire [4:0] my_ivn2_io_o_vn2_0; // @[ivntop.scala 78:24]
  wire [4:0] my_ivn2_io_o_vn2_1; // @[ivntop.scala 78:24]
  wire [4:0] my_ivn2_io_o_vn2_2; // @[ivntop.scala 78:24]
  wire [4:0] my_ivn2_io_o_vn2_3; // @[ivntop.scala 78:24]
  wire  my_ivn2_io_validpin; // @[ivntop.scala 78:24]
  wire  my_ivn3_clock; // @[ivntop.scala 86:25]
  wire  my_ivn3_reset; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_0_0; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_0_1; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_0_2; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_0_3; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_0_4; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_0_5; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_0_6; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_0_7; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_1_0; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_1_1; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_1_2; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_1_3; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_1_4; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_1_5; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_1_6; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_1_7; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_2_0; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_2_1; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_2_2; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_2_3; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_2_4; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_2_5; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_2_6; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_2_7; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_3_0; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_3_1; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_3_2; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_3_3; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_3_4; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_3_5; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_3_6; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_3_7; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_4_0; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_4_1; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_4_2; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_4_3; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_4_4; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_4_5; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_4_6; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_4_7; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_5_0; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_5_1; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_5_2; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_5_3; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_5_4; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_5_5; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_5_6; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_5_7; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_6_0; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_6_1; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_6_2; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_6_3; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_6_4; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_6_5; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_6_6; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_6_7; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_7_0; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_7_1; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_7_2; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_7_3; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_7_4; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_7_5; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_7_6; // @[ivntop.scala 86:25]
  wire [15:0] my_ivn3_io_Stationary_matrix_7_7; // @[ivntop.scala 86:25]
  wire [4:0] my_ivn3_io_o_vn_0; // @[ivntop.scala 86:25]
  wire [4:0] my_ivn3_io_o_vn_1; // @[ivntop.scala 86:25]
  wire [4:0] my_ivn3_io_o_vn_2; // @[ivntop.scala 86:25]
  wire [4:0] my_ivn3_io_o_vn_3; // @[ivntop.scala 86:25]
  wire [4:0] my_ivn3_io_o_vn2_0; // @[ivntop.scala 86:25]
  wire [4:0] my_ivn3_io_o_vn2_1; // @[ivntop.scala 86:25]
  wire [4:0] my_ivn3_io_o_vn2_2; // @[ivntop.scala 86:25]
  wire [4:0] my_ivn3_io_o_vn2_3; // @[ivntop.scala 86:25]
  wire  my_ivn3_io_validpin; // @[ivntop.scala 86:25]
  wire  my_ivn4_clock; // @[ivntop.scala 93:25]
  wire  my_ivn4_reset; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_0_0; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_0_1; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_0_2; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_0_3; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_0_4; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_0_5; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_0_6; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_0_7; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_1_0; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_1_1; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_1_2; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_1_3; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_1_4; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_1_5; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_1_6; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_1_7; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_2_0; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_2_1; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_2_2; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_2_3; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_2_4; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_2_5; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_2_6; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_2_7; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_3_0; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_3_1; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_3_2; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_3_3; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_3_4; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_3_5; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_3_6; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_3_7; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_4_0; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_4_1; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_4_2; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_4_3; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_4_4; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_4_5; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_4_6; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_4_7; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_5_0; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_5_1; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_5_2; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_5_3; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_5_4; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_5_5; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_5_6; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_5_7; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_6_0; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_6_1; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_6_2; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_6_3; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_6_4; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_6_5; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_6_6; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_6_7; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_7_0; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_7_1; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_7_2; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_7_3; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_7_4; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_7_5; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_7_6; // @[ivntop.scala 93:25]
  wire [15:0] my_ivn4_io_Stationary_matrix_7_7; // @[ivntop.scala 93:25]
  wire [4:0] my_ivn4_io_o_vn_0; // @[ivntop.scala 93:25]
  wire [4:0] my_ivn4_io_o_vn_1; // @[ivntop.scala 93:25]
  wire [4:0] my_ivn4_io_o_vn_2; // @[ivntop.scala 93:25]
  wire [4:0] my_ivn4_io_o_vn_3; // @[ivntop.scala 93:25]
  wire [4:0] my_ivn4_io_o_vn2_0; // @[ivntop.scala 93:25]
  wire [4:0] my_ivn4_io_o_vn2_1; // @[ivntop.scala 93:25]
  wire [4:0] my_ivn4_io_o_vn2_2; // @[ivntop.scala 93:25]
  wire [4:0] my_ivn4_io_o_vn2_3; // @[ivntop.scala 93:25]
  wire  my_ivn4_io_validpin; // @[ivntop.scala 93:25]
  wire  my_ivn5_clock; // @[ivntop.scala 100:25]
  wire  my_ivn5_reset; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_0_0; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_0_1; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_0_2; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_0_3; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_0_4; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_0_5; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_0_6; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_0_7; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_1_0; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_1_1; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_1_2; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_1_3; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_1_4; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_1_5; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_1_6; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_1_7; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_2_0; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_2_1; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_2_2; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_2_3; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_2_4; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_2_5; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_2_6; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_2_7; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_3_0; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_3_1; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_3_2; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_3_3; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_3_4; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_3_5; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_3_6; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_3_7; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_4_0; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_4_1; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_4_2; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_4_3; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_4_4; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_4_5; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_4_6; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_4_7; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_5_0; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_5_1; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_5_2; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_5_3; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_5_4; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_5_5; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_5_6; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_5_7; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_6_0; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_6_1; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_6_2; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_6_3; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_6_4; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_6_5; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_6_6; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_6_7; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_7_0; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_7_1; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_7_2; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_7_3; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_7_4; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_7_5; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_7_6; // @[ivntop.scala 100:25]
  wire [15:0] my_ivn5_io_Stationary_matrix_7_7; // @[ivntop.scala 100:25]
  wire [4:0] my_ivn5_io_o_vn_0; // @[ivntop.scala 100:25]
  wire [4:0] my_ivn5_io_o_vn_1; // @[ivntop.scala 100:25]
  wire [4:0] my_ivn5_io_o_vn_2; // @[ivntop.scala 100:25]
  wire [4:0] my_ivn5_io_o_vn_3; // @[ivntop.scala 100:25]
  wire [4:0] my_ivn5_io_o_vn2_0; // @[ivntop.scala 100:25]
  wire [4:0] my_ivn5_io_o_vn2_1; // @[ivntop.scala 100:25]
  wire [4:0] my_ivn5_io_o_vn2_2; // @[ivntop.scala 100:25]
  wire [4:0] my_ivn5_io_o_vn2_3; // @[ivntop.scala 100:25]
  wire  my_ivn5_io_validpin; // @[ivntop.scala 100:25]
  wire  my_ivn6_clock; // @[ivntop.scala 107:25]
  wire  my_ivn6_reset; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_0_0; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_0_1; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_0_2; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_0_3; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_0_4; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_0_5; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_0_6; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_0_7; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_1_0; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_1_1; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_1_2; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_1_3; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_1_4; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_1_5; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_1_6; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_1_7; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_2_0; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_2_1; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_2_2; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_2_3; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_2_4; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_2_5; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_2_6; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_2_7; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_3_0; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_3_1; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_3_2; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_3_3; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_3_4; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_3_5; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_3_6; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_3_7; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_4_0; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_4_1; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_4_2; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_4_3; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_4_4; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_4_5; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_4_6; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_4_7; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_5_0; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_5_1; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_5_2; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_5_3; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_5_4; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_5_5; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_5_6; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_5_7; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_6_0; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_6_1; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_6_2; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_6_3; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_6_4; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_6_5; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_6_6; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_6_7; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_7_0; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_7_1; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_7_2; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_7_3; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_7_4; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_7_5; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_7_6; // @[ivntop.scala 107:25]
  wire [15:0] my_ivn6_io_Stationary_matrix_7_7; // @[ivntop.scala 107:25]
  wire [4:0] my_ivn6_io_o_vn_0; // @[ivntop.scala 107:25]
  wire [4:0] my_ivn6_io_o_vn_1; // @[ivntop.scala 107:25]
  wire [4:0] my_ivn6_io_o_vn_2; // @[ivntop.scala 107:25]
  wire [4:0] my_ivn6_io_o_vn_3; // @[ivntop.scala 107:25]
  wire [4:0] my_ivn6_io_o_vn2_0; // @[ivntop.scala 107:25]
  wire [4:0] my_ivn6_io_o_vn2_1; // @[ivntop.scala 107:25]
  wire [4:0] my_ivn6_io_o_vn2_2; // @[ivntop.scala 107:25]
  wire [4:0] my_ivn6_io_o_vn2_3; // @[ivntop.scala 107:25]
  wire  my_ivn6_io_validpin; // @[ivntop.scala 107:25]
  wire  my_ivn7_clock; // @[ivntop.scala 114:25]
  wire  my_ivn7_reset; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_0_0; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_0_1; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_0_2; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_0_3; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_0_4; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_0_5; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_0_6; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_0_7; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_1_0; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_1_1; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_1_2; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_1_3; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_1_4; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_1_5; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_1_6; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_1_7; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_2_0; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_2_1; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_2_2; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_2_3; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_2_4; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_2_5; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_2_6; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_2_7; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_3_0; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_3_1; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_3_2; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_3_3; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_3_4; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_3_5; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_3_6; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_3_7; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_4_0; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_4_1; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_4_2; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_4_3; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_4_4; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_4_5; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_4_6; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_4_7; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_5_0; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_5_1; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_5_2; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_5_3; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_5_4; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_5_5; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_5_6; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_5_7; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_6_0; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_6_1; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_6_2; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_6_3; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_6_4; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_6_5; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_6_6; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_6_7; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_7_0; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_7_1; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_7_2; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_7_3; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_7_4; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_7_5; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_7_6; // @[ivntop.scala 114:25]
  wire [15:0] my_ivn7_io_Stationary_matrix_7_7; // @[ivntop.scala 114:25]
  wire [4:0] my_ivn7_io_o_vn_0; // @[ivntop.scala 114:25]
  wire [4:0] my_ivn7_io_o_vn_1; // @[ivntop.scala 114:25]
  wire [4:0] my_ivn7_io_o_vn_2; // @[ivntop.scala 114:25]
  wire [4:0] my_ivn7_io_o_vn_3; // @[ivntop.scala 114:25]
  wire [4:0] my_ivn7_io_o_vn2_0; // @[ivntop.scala 114:25]
  wire [4:0] my_ivn7_io_o_vn2_1; // @[ivntop.scala 114:25]
  wire [4:0] my_ivn7_io_o_vn2_2; // @[ivntop.scala 114:25]
  wire [4:0] my_ivn7_io_o_vn2_3; // @[ivntop.scala 114:25]
  wire  my_ivn7_io_validpin; // @[ivntop.scala 114:25]
  wire  my_ivn8_clock; // @[ivntop.scala 121:25]
  wire  my_ivn8_reset; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_0_0; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_0_1; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_0_2; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_0_3; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_0_4; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_0_5; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_0_6; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_0_7; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_1_0; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_1_1; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_1_2; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_1_3; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_1_4; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_1_5; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_1_6; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_1_7; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_2_0; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_2_1; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_2_2; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_2_3; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_2_4; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_2_5; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_2_6; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_2_7; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_3_0; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_3_1; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_3_2; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_3_3; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_3_4; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_3_5; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_3_6; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_3_7; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_4_0; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_4_1; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_4_2; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_4_3; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_4_4; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_4_5; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_4_6; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_4_7; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_5_0; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_5_1; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_5_2; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_5_3; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_5_4; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_5_5; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_5_6; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_5_7; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_6_0; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_6_1; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_6_2; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_6_3; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_6_4; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_6_5; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_6_6; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_6_7; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_7_0; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_7_1; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_7_2; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_7_3; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_7_4; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_7_5; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_7_6; // @[ivntop.scala 121:25]
  wire [15:0] my_ivn8_io_Stationary_matrix_7_7; // @[ivntop.scala 121:25]
  wire [4:0] my_ivn8_io_o_vn_0; // @[ivntop.scala 121:25]
  wire [4:0] my_ivn8_io_o_vn_1; // @[ivntop.scala 121:25]
  wire [4:0] my_ivn8_io_o_vn_2; // @[ivntop.scala 121:25]
  wire [4:0] my_ivn8_io_o_vn_3; // @[ivntop.scala 121:25]
  wire [4:0] my_ivn8_io_o_vn2_0; // @[ivntop.scala 121:25]
  wire [4:0] my_ivn8_io_o_vn2_1; // @[ivntop.scala 121:25]
  wire [4:0] my_ivn8_io_o_vn2_2; // @[ivntop.scala 121:25]
  wire [4:0] my_ivn8_io_o_vn2_3; // @[ivntop.scala 121:25]
  wire  my_ivn8_io_validpin; // @[ivntop.scala 121:25]
  reg [4:0] i_vn_0_0; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_0_1; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_0_2; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_0_3; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_1_0; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_1_1; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_1_2; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_1_3; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_2_0; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_2_1; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_2_2; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_2_3; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_3_0; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_3_1; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_3_2; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_3_3; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_4_0; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_4_1; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_4_2; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_4_3; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_5_0; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_5_1; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_5_2; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_5_3; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_6_0; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_6_1; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_6_2; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_6_3; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_7_0; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_7_1; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_7_2; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_7_3; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_8_0; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_8_1; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_8_2; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_8_3; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_9_0; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_9_1; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_9_2; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_9_3; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_10_0; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_10_1; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_10_2; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_10_3; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_11_0; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_11_1; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_11_2; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_11_3; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_12_0; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_12_1; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_12_2; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_12_3; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_13_0; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_13_1; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_13_2; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_13_3; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_14_0; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_14_1; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_14_2; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_14_3; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_15_0; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_15_1; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_15_2; // @[ivntop.scala 15:17]
  reg [4:0] i_vn_15_3; // @[ivntop.scala 15:17]
  reg [31:0] counter; // @[ivntop.scala 27:26]
  wire  _T = 1'h1; // @[ivntop.scala 40:16]
  wire [31:0] _counter_T_1 = counter + 32'h1; // @[ivntop.scala 156:22]
  wire  valid = 1'h1; // @[ivntop.scala 40:22 41:11]
  stationary my_stationary ( // @[ivntop.scala 29:31]
    .clock(my_stationary_clock),
    .reset(my_stationary_reset),
    .io_Stationary_matrix_0_0(my_stationary_io_Stationary_matrix_0_0),
    .io_Stationary_matrix_0_1(my_stationary_io_Stationary_matrix_0_1),
    .io_Stationary_matrix_0_2(my_stationary_io_Stationary_matrix_0_2),
    .io_Stationary_matrix_0_3(my_stationary_io_Stationary_matrix_0_3),
    .io_Stationary_matrix_0_4(my_stationary_io_Stationary_matrix_0_4),
    .io_Stationary_matrix_0_5(my_stationary_io_Stationary_matrix_0_5),
    .io_Stationary_matrix_0_6(my_stationary_io_Stationary_matrix_0_6),
    .io_Stationary_matrix_0_7(my_stationary_io_Stationary_matrix_0_7),
    .io_Stationary_matrix_1_0(my_stationary_io_Stationary_matrix_1_0),
    .io_Stationary_matrix_1_1(my_stationary_io_Stationary_matrix_1_1),
    .io_Stationary_matrix_1_2(my_stationary_io_Stationary_matrix_1_2),
    .io_Stationary_matrix_1_3(my_stationary_io_Stationary_matrix_1_3),
    .io_Stationary_matrix_1_4(my_stationary_io_Stationary_matrix_1_4),
    .io_Stationary_matrix_1_5(my_stationary_io_Stationary_matrix_1_5),
    .io_Stationary_matrix_1_6(my_stationary_io_Stationary_matrix_1_6),
    .io_Stationary_matrix_1_7(my_stationary_io_Stationary_matrix_1_7),
    .io_Stationary_matrix_2_0(my_stationary_io_Stationary_matrix_2_0),
    .io_Stationary_matrix_2_1(my_stationary_io_Stationary_matrix_2_1),
    .io_Stationary_matrix_2_2(my_stationary_io_Stationary_matrix_2_2),
    .io_Stationary_matrix_2_3(my_stationary_io_Stationary_matrix_2_3),
    .io_Stationary_matrix_2_4(my_stationary_io_Stationary_matrix_2_4),
    .io_Stationary_matrix_2_5(my_stationary_io_Stationary_matrix_2_5),
    .io_Stationary_matrix_2_6(my_stationary_io_Stationary_matrix_2_6),
    .io_Stationary_matrix_2_7(my_stationary_io_Stationary_matrix_2_7),
    .io_Stationary_matrix_3_0(my_stationary_io_Stationary_matrix_3_0),
    .io_Stationary_matrix_3_1(my_stationary_io_Stationary_matrix_3_1),
    .io_Stationary_matrix_3_2(my_stationary_io_Stationary_matrix_3_2),
    .io_Stationary_matrix_3_3(my_stationary_io_Stationary_matrix_3_3),
    .io_Stationary_matrix_3_4(my_stationary_io_Stationary_matrix_3_4),
    .io_Stationary_matrix_3_5(my_stationary_io_Stationary_matrix_3_5),
    .io_Stationary_matrix_3_6(my_stationary_io_Stationary_matrix_3_6),
    .io_Stationary_matrix_3_7(my_stationary_io_Stationary_matrix_3_7),
    .io_Stationary_matrix_4_0(my_stationary_io_Stationary_matrix_4_0),
    .io_Stationary_matrix_4_1(my_stationary_io_Stationary_matrix_4_1),
    .io_Stationary_matrix_4_2(my_stationary_io_Stationary_matrix_4_2),
    .io_Stationary_matrix_4_3(my_stationary_io_Stationary_matrix_4_3),
    .io_Stationary_matrix_4_4(my_stationary_io_Stationary_matrix_4_4),
    .io_Stationary_matrix_4_5(my_stationary_io_Stationary_matrix_4_5),
    .io_Stationary_matrix_4_6(my_stationary_io_Stationary_matrix_4_6),
    .io_Stationary_matrix_4_7(my_stationary_io_Stationary_matrix_4_7),
    .io_Stationary_matrix_5_0(my_stationary_io_Stationary_matrix_5_0),
    .io_Stationary_matrix_5_1(my_stationary_io_Stationary_matrix_5_1),
    .io_Stationary_matrix_5_2(my_stationary_io_Stationary_matrix_5_2),
    .io_Stationary_matrix_5_3(my_stationary_io_Stationary_matrix_5_3),
    .io_Stationary_matrix_5_4(my_stationary_io_Stationary_matrix_5_4),
    .io_Stationary_matrix_5_5(my_stationary_io_Stationary_matrix_5_5),
    .io_Stationary_matrix_5_6(my_stationary_io_Stationary_matrix_5_6),
    .io_Stationary_matrix_5_7(my_stationary_io_Stationary_matrix_5_7),
    .io_Stationary_matrix_6_0(my_stationary_io_Stationary_matrix_6_0),
    .io_Stationary_matrix_6_1(my_stationary_io_Stationary_matrix_6_1),
    .io_Stationary_matrix_6_2(my_stationary_io_Stationary_matrix_6_2),
    .io_Stationary_matrix_6_3(my_stationary_io_Stationary_matrix_6_3),
    .io_Stationary_matrix_6_4(my_stationary_io_Stationary_matrix_6_4),
    .io_Stationary_matrix_6_5(my_stationary_io_Stationary_matrix_6_5),
    .io_Stationary_matrix_6_6(my_stationary_io_Stationary_matrix_6_6),
    .io_Stationary_matrix_6_7(my_stationary_io_Stationary_matrix_6_7),
    .io_Stationary_matrix_7_0(my_stationary_io_Stationary_matrix_7_0),
    .io_Stationary_matrix_7_1(my_stationary_io_Stationary_matrix_7_1),
    .io_Stationary_matrix_7_2(my_stationary_io_Stationary_matrix_7_2),
    .io_Stationary_matrix_7_3(my_stationary_io_Stationary_matrix_7_3),
    .io_Stationary_matrix_7_4(my_stationary_io_Stationary_matrix_7_4),
    .io_Stationary_matrix_7_5(my_stationary_io_Stationary_matrix_7_5),
    .io_Stationary_matrix_7_6(my_stationary_io_Stationary_matrix_7_6),
    .io_Stationary_matrix_7_7(my_stationary_io_Stationary_matrix_7_7),
    .io_o_Stationary_matrix1_0_0(my_stationary_io_o_Stationary_matrix1_0_0),
    .io_o_Stationary_matrix1_0_1(my_stationary_io_o_Stationary_matrix1_0_1),
    .io_o_Stationary_matrix1_0_2(my_stationary_io_o_Stationary_matrix1_0_2),
    .io_o_Stationary_matrix1_0_3(my_stationary_io_o_Stationary_matrix1_0_3),
    .io_o_Stationary_matrix1_0_4(my_stationary_io_o_Stationary_matrix1_0_4),
    .io_o_Stationary_matrix1_0_5(my_stationary_io_o_Stationary_matrix1_0_5),
    .io_o_Stationary_matrix1_0_6(my_stationary_io_o_Stationary_matrix1_0_6),
    .io_o_Stationary_matrix1_0_7(my_stationary_io_o_Stationary_matrix1_0_7),
    .io_o_Stationary_matrix1_1_0(my_stationary_io_o_Stationary_matrix1_1_0),
    .io_o_Stationary_matrix1_1_1(my_stationary_io_o_Stationary_matrix1_1_1),
    .io_o_Stationary_matrix1_1_2(my_stationary_io_o_Stationary_matrix1_1_2),
    .io_o_Stationary_matrix1_1_3(my_stationary_io_o_Stationary_matrix1_1_3),
    .io_o_Stationary_matrix1_1_4(my_stationary_io_o_Stationary_matrix1_1_4),
    .io_o_Stationary_matrix1_1_5(my_stationary_io_o_Stationary_matrix1_1_5),
    .io_o_Stationary_matrix1_1_6(my_stationary_io_o_Stationary_matrix1_1_6),
    .io_o_Stationary_matrix1_1_7(my_stationary_io_o_Stationary_matrix1_1_7),
    .io_o_Stationary_matrix1_2_0(my_stationary_io_o_Stationary_matrix1_2_0),
    .io_o_Stationary_matrix1_2_1(my_stationary_io_o_Stationary_matrix1_2_1),
    .io_o_Stationary_matrix1_2_2(my_stationary_io_o_Stationary_matrix1_2_2),
    .io_o_Stationary_matrix1_2_3(my_stationary_io_o_Stationary_matrix1_2_3),
    .io_o_Stationary_matrix1_2_4(my_stationary_io_o_Stationary_matrix1_2_4),
    .io_o_Stationary_matrix1_2_5(my_stationary_io_o_Stationary_matrix1_2_5),
    .io_o_Stationary_matrix1_2_6(my_stationary_io_o_Stationary_matrix1_2_6),
    .io_o_Stationary_matrix1_2_7(my_stationary_io_o_Stationary_matrix1_2_7),
    .io_o_Stationary_matrix1_3_0(my_stationary_io_o_Stationary_matrix1_3_0),
    .io_o_Stationary_matrix1_3_1(my_stationary_io_o_Stationary_matrix1_3_1),
    .io_o_Stationary_matrix1_3_2(my_stationary_io_o_Stationary_matrix1_3_2),
    .io_o_Stationary_matrix1_3_3(my_stationary_io_o_Stationary_matrix1_3_3),
    .io_o_Stationary_matrix1_3_4(my_stationary_io_o_Stationary_matrix1_3_4),
    .io_o_Stationary_matrix1_3_5(my_stationary_io_o_Stationary_matrix1_3_5),
    .io_o_Stationary_matrix1_3_6(my_stationary_io_o_Stationary_matrix1_3_6),
    .io_o_Stationary_matrix1_3_7(my_stationary_io_o_Stationary_matrix1_3_7),
    .io_o_Stationary_matrix1_4_0(my_stationary_io_o_Stationary_matrix1_4_0),
    .io_o_Stationary_matrix1_4_1(my_stationary_io_o_Stationary_matrix1_4_1),
    .io_o_Stationary_matrix1_4_2(my_stationary_io_o_Stationary_matrix1_4_2),
    .io_o_Stationary_matrix1_4_3(my_stationary_io_o_Stationary_matrix1_4_3),
    .io_o_Stationary_matrix1_4_4(my_stationary_io_o_Stationary_matrix1_4_4),
    .io_o_Stationary_matrix1_4_5(my_stationary_io_o_Stationary_matrix1_4_5),
    .io_o_Stationary_matrix1_4_6(my_stationary_io_o_Stationary_matrix1_4_6),
    .io_o_Stationary_matrix1_4_7(my_stationary_io_o_Stationary_matrix1_4_7),
    .io_o_Stationary_matrix1_5_0(my_stationary_io_o_Stationary_matrix1_5_0),
    .io_o_Stationary_matrix1_5_1(my_stationary_io_o_Stationary_matrix1_5_1),
    .io_o_Stationary_matrix1_5_2(my_stationary_io_o_Stationary_matrix1_5_2),
    .io_o_Stationary_matrix1_5_3(my_stationary_io_o_Stationary_matrix1_5_3),
    .io_o_Stationary_matrix1_5_4(my_stationary_io_o_Stationary_matrix1_5_4),
    .io_o_Stationary_matrix1_5_5(my_stationary_io_o_Stationary_matrix1_5_5),
    .io_o_Stationary_matrix1_5_6(my_stationary_io_o_Stationary_matrix1_5_6),
    .io_o_Stationary_matrix1_5_7(my_stationary_io_o_Stationary_matrix1_5_7),
    .io_o_Stationary_matrix1_6_0(my_stationary_io_o_Stationary_matrix1_6_0),
    .io_o_Stationary_matrix1_6_1(my_stationary_io_o_Stationary_matrix1_6_1),
    .io_o_Stationary_matrix1_6_2(my_stationary_io_o_Stationary_matrix1_6_2),
    .io_o_Stationary_matrix1_6_3(my_stationary_io_o_Stationary_matrix1_6_3),
    .io_o_Stationary_matrix1_6_4(my_stationary_io_o_Stationary_matrix1_6_4),
    .io_o_Stationary_matrix1_6_5(my_stationary_io_o_Stationary_matrix1_6_5),
    .io_o_Stationary_matrix1_6_6(my_stationary_io_o_Stationary_matrix1_6_6),
    .io_o_Stationary_matrix1_6_7(my_stationary_io_o_Stationary_matrix1_6_7),
    .io_o_Stationary_matrix1_7_0(my_stationary_io_o_Stationary_matrix1_7_0),
    .io_o_Stationary_matrix1_7_1(my_stationary_io_o_Stationary_matrix1_7_1),
    .io_o_Stationary_matrix1_7_2(my_stationary_io_o_Stationary_matrix1_7_2),
    .io_o_Stationary_matrix1_7_3(my_stationary_io_o_Stationary_matrix1_7_3),
    .io_o_Stationary_matrix1_7_4(my_stationary_io_o_Stationary_matrix1_7_4),
    .io_o_Stationary_matrix1_7_5(my_stationary_io_o_Stationary_matrix1_7_5),
    .io_o_Stationary_matrix1_7_6(my_stationary_io_o_Stationary_matrix1_7_6),
    .io_o_Stationary_matrix1_7_7(my_stationary_io_o_Stationary_matrix1_7_7),
    .io_o_Stationary_matrix2_0_0(my_stationary_io_o_Stationary_matrix2_0_0),
    .io_o_Stationary_matrix2_0_1(my_stationary_io_o_Stationary_matrix2_0_1),
    .io_o_Stationary_matrix2_0_2(my_stationary_io_o_Stationary_matrix2_0_2),
    .io_o_Stationary_matrix2_0_3(my_stationary_io_o_Stationary_matrix2_0_3),
    .io_o_Stationary_matrix2_0_4(my_stationary_io_o_Stationary_matrix2_0_4),
    .io_o_Stationary_matrix2_0_5(my_stationary_io_o_Stationary_matrix2_0_5),
    .io_o_Stationary_matrix2_0_6(my_stationary_io_o_Stationary_matrix2_0_6),
    .io_o_Stationary_matrix2_0_7(my_stationary_io_o_Stationary_matrix2_0_7),
    .io_o_Stationary_matrix2_1_0(my_stationary_io_o_Stationary_matrix2_1_0),
    .io_o_Stationary_matrix2_1_1(my_stationary_io_o_Stationary_matrix2_1_1),
    .io_o_Stationary_matrix2_1_2(my_stationary_io_o_Stationary_matrix2_1_2),
    .io_o_Stationary_matrix2_1_3(my_stationary_io_o_Stationary_matrix2_1_3),
    .io_o_Stationary_matrix2_1_4(my_stationary_io_o_Stationary_matrix2_1_4),
    .io_o_Stationary_matrix2_1_5(my_stationary_io_o_Stationary_matrix2_1_5),
    .io_o_Stationary_matrix2_1_6(my_stationary_io_o_Stationary_matrix2_1_6),
    .io_o_Stationary_matrix2_1_7(my_stationary_io_o_Stationary_matrix2_1_7),
    .io_o_Stationary_matrix2_2_0(my_stationary_io_o_Stationary_matrix2_2_0),
    .io_o_Stationary_matrix2_2_1(my_stationary_io_o_Stationary_matrix2_2_1),
    .io_o_Stationary_matrix2_2_2(my_stationary_io_o_Stationary_matrix2_2_2),
    .io_o_Stationary_matrix2_2_3(my_stationary_io_o_Stationary_matrix2_2_3),
    .io_o_Stationary_matrix2_2_4(my_stationary_io_o_Stationary_matrix2_2_4),
    .io_o_Stationary_matrix2_2_5(my_stationary_io_o_Stationary_matrix2_2_5),
    .io_o_Stationary_matrix2_2_6(my_stationary_io_o_Stationary_matrix2_2_6),
    .io_o_Stationary_matrix2_2_7(my_stationary_io_o_Stationary_matrix2_2_7),
    .io_o_Stationary_matrix2_3_0(my_stationary_io_o_Stationary_matrix2_3_0),
    .io_o_Stationary_matrix2_3_1(my_stationary_io_o_Stationary_matrix2_3_1),
    .io_o_Stationary_matrix2_3_2(my_stationary_io_o_Stationary_matrix2_3_2),
    .io_o_Stationary_matrix2_3_3(my_stationary_io_o_Stationary_matrix2_3_3),
    .io_o_Stationary_matrix2_3_4(my_stationary_io_o_Stationary_matrix2_3_4),
    .io_o_Stationary_matrix2_3_5(my_stationary_io_o_Stationary_matrix2_3_5),
    .io_o_Stationary_matrix2_3_6(my_stationary_io_o_Stationary_matrix2_3_6),
    .io_o_Stationary_matrix2_3_7(my_stationary_io_o_Stationary_matrix2_3_7),
    .io_o_Stationary_matrix2_4_0(my_stationary_io_o_Stationary_matrix2_4_0),
    .io_o_Stationary_matrix2_4_1(my_stationary_io_o_Stationary_matrix2_4_1),
    .io_o_Stationary_matrix2_4_2(my_stationary_io_o_Stationary_matrix2_4_2),
    .io_o_Stationary_matrix2_4_3(my_stationary_io_o_Stationary_matrix2_4_3),
    .io_o_Stationary_matrix2_4_4(my_stationary_io_o_Stationary_matrix2_4_4),
    .io_o_Stationary_matrix2_4_5(my_stationary_io_o_Stationary_matrix2_4_5),
    .io_o_Stationary_matrix2_4_6(my_stationary_io_o_Stationary_matrix2_4_6),
    .io_o_Stationary_matrix2_4_7(my_stationary_io_o_Stationary_matrix2_4_7),
    .io_o_Stationary_matrix2_5_0(my_stationary_io_o_Stationary_matrix2_5_0),
    .io_o_Stationary_matrix2_5_1(my_stationary_io_o_Stationary_matrix2_5_1),
    .io_o_Stationary_matrix2_5_2(my_stationary_io_o_Stationary_matrix2_5_2),
    .io_o_Stationary_matrix2_5_3(my_stationary_io_o_Stationary_matrix2_5_3),
    .io_o_Stationary_matrix2_5_4(my_stationary_io_o_Stationary_matrix2_5_4),
    .io_o_Stationary_matrix2_5_5(my_stationary_io_o_Stationary_matrix2_5_5),
    .io_o_Stationary_matrix2_5_6(my_stationary_io_o_Stationary_matrix2_5_6),
    .io_o_Stationary_matrix2_5_7(my_stationary_io_o_Stationary_matrix2_5_7),
    .io_o_Stationary_matrix2_6_0(my_stationary_io_o_Stationary_matrix2_6_0),
    .io_o_Stationary_matrix2_6_1(my_stationary_io_o_Stationary_matrix2_6_1),
    .io_o_Stationary_matrix2_6_2(my_stationary_io_o_Stationary_matrix2_6_2),
    .io_o_Stationary_matrix2_6_3(my_stationary_io_o_Stationary_matrix2_6_3),
    .io_o_Stationary_matrix2_6_4(my_stationary_io_o_Stationary_matrix2_6_4),
    .io_o_Stationary_matrix2_6_5(my_stationary_io_o_Stationary_matrix2_6_5),
    .io_o_Stationary_matrix2_6_6(my_stationary_io_o_Stationary_matrix2_6_6),
    .io_o_Stationary_matrix2_6_7(my_stationary_io_o_Stationary_matrix2_6_7),
    .io_o_Stationary_matrix2_7_0(my_stationary_io_o_Stationary_matrix2_7_0),
    .io_o_Stationary_matrix2_7_1(my_stationary_io_o_Stationary_matrix2_7_1),
    .io_o_Stationary_matrix2_7_2(my_stationary_io_o_Stationary_matrix2_7_2),
    .io_o_Stationary_matrix2_7_3(my_stationary_io_o_Stationary_matrix2_7_3),
    .io_o_Stationary_matrix2_7_4(my_stationary_io_o_Stationary_matrix2_7_4),
    .io_o_Stationary_matrix2_7_5(my_stationary_io_o_Stationary_matrix2_7_5),
    .io_o_Stationary_matrix2_7_6(my_stationary_io_o_Stationary_matrix2_7_6),
    .io_o_Stationary_matrix2_7_7(my_stationary_io_o_Stationary_matrix2_7_7),
    .io_o_Stationary_matrix3_0_0(my_stationary_io_o_Stationary_matrix3_0_0),
    .io_o_Stationary_matrix3_0_1(my_stationary_io_o_Stationary_matrix3_0_1),
    .io_o_Stationary_matrix3_0_2(my_stationary_io_o_Stationary_matrix3_0_2),
    .io_o_Stationary_matrix3_0_3(my_stationary_io_o_Stationary_matrix3_0_3),
    .io_o_Stationary_matrix3_0_4(my_stationary_io_o_Stationary_matrix3_0_4),
    .io_o_Stationary_matrix3_0_5(my_stationary_io_o_Stationary_matrix3_0_5),
    .io_o_Stationary_matrix3_0_6(my_stationary_io_o_Stationary_matrix3_0_6),
    .io_o_Stationary_matrix3_0_7(my_stationary_io_o_Stationary_matrix3_0_7),
    .io_o_Stationary_matrix3_1_0(my_stationary_io_o_Stationary_matrix3_1_0),
    .io_o_Stationary_matrix3_1_1(my_stationary_io_o_Stationary_matrix3_1_1),
    .io_o_Stationary_matrix3_1_2(my_stationary_io_o_Stationary_matrix3_1_2),
    .io_o_Stationary_matrix3_1_3(my_stationary_io_o_Stationary_matrix3_1_3),
    .io_o_Stationary_matrix3_1_4(my_stationary_io_o_Stationary_matrix3_1_4),
    .io_o_Stationary_matrix3_1_5(my_stationary_io_o_Stationary_matrix3_1_5),
    .io_o_Stationary_matrix3_1_6(my_stationary_io_o_Stationary_matrix3_1_6),
    .io_o_Stationary_matrix3_1_7(my_stationary_io_o_Stationary_matrix3_1_7),
    .io_o_Stationary_matrix3_2_0(my_stationary_io_o_Stationary_matrix3_2_0),
    .io_o_Stationary_matrix3_2_1(my_stationary_io_o_Stationary_matrix3_2_1),
    .io_o_Stationary_matrix3_2_2(my_stationary_io_o_Stationary_matrix3_2_2),
    .io_o_Stationary_matrix3_2_3(my_stationary_io_o_Stationary_matrix3_2_3),
    .io_o_Stationary_matrix3_2_4(my_stationary_io_o_Stationary_matrix3_2_4),
    .io_o_Stationary_matrix3_2_5(my_stationary_io_o_Stationary_matrix3_2_5),
    .io_o_Stationary_matrix3_2_6(my_stationary_io_o_Stationary_matrix3_2_6),
    .io_o_Stationary_matrix3_2_7(my_stationary_io_o_Stationary_matrix3_2_7),
    .io_o_Stationary_matrix3_3_0(my_stationary_io_o_Stationary_matrix3_3_0),
    .io_o_Stationary_matrix3_3_1(my_stationary_io_o_Stationary_matrix3_3_1),
    .io_o_Stationary_matrix3_3_2(my_stationary_io_o_Stationary_matrix3_3_2),
    .io_o_Stationary_matrix3_3_3(my_stationary_io_o_Stationary_matrix3_3_3),
    .io_o_Stationary_matrix3_3_4(my_stationary_io_o_Stationary_matrix3_3_4),
    .io_o_Stationary_matrix3_3_5(my_stationary_io_o_Stationary_matrix3_3_5),
    .io_o_Stationary_matrix3_3_6(my_stationary_io_o_Stationary_matrix3_3_6),
    .io_o_Stationary_matrix3_3_7(my_stationary_io_o_Stationary_matrix3_3_7),
    .io_o_Stationary_matrix3_4_0(my_stationary_io_o_Stationary_matrix3_4_0),
    .io_o_Stationary_matrix3_4_1(my_stationary_io_o_Stationary_matrix3_4_1),
    .io_o_Stationary_matrix3_4_2(my_stationary_io_o_Stationary_matrix3_4_2),
    .io_o_Stationary_matrix3_4_3(my_stationary_io_o_Stationary_matrix3_4_3),
    .io_o_Stationary_matrix3_4_4(my_stationary_io_o_Stationary_matrix3_4_4),
    .io_o_Stationary_matrix3_4_5(my_stationary_io_o_Stationary_matrix3_4_5),
    .io_o_Stationary_matrix3_4_6(my_stationary_io_o_Stationary_matrix3_4_6),
    .io_o_Stationary_matrix3_4_7(my_stationary_io_o_Stationary_matrix3_4_7),
    .io_o_Stationary_matrix3_5_0(my_stationary_io_o_Stationary_matrix3_5_0),
    .io_o_Stationary_matrix3_5_1(my_stationary_io_o_Stationary_matrix3_5_1),
    .io_o_Stationary_matrix3_5_2(my_stationary_io_o_Stationary_matrix3_5_2),
    .io_o_Stationary_matrix3_5_3(my_stationary_io_o_Stationary_matrix3_5_3),
    .io_o_Stationary_matrix3_5_4(my_stationary_io_o_Stationary_matrix3_5_4),
    .io_o_Stationary_matrix3_5_5(my_stationary_io_o_Stationary_matrix3_5_5),
    .io_o_Stationary_matrix3_5_6(my_stationary_io_o_Stationary_matrix3_5_6),
    .io_o_Stationary_matrix3_5_7(my_stationary_io_o_Stationary_matrix3_5_7),
    .io_o_Stationary_matrix3_6_0(my_stationary_io_o_Stationary_matrix3_6_0),
    .io_o_Stationary_matrix3_6_1(my_stationary_io_o_Stationary_matrix3_6_1),
    .io_o_Stationary_matrix3_6_2(my_stationary_io_o_Stationary_matrix3_6_2),
    .io_o_Stationary_matrix3_6_3(my_stationary_io_o_Stationary_matrix3_6_3),
    .io_o_Stationary_matrix3_6_4(my_stationary_io_o_Stationary_matrix3_6_4),
    .io_o_Stationary_matrix3_6_5(my_stationary_io_o_Stationary_matrix3_6_5),
    .io_o_Stationary_matrix3_6_6(my_stationary_io_o_Stationary_matrix3_6_6),
    .io_o_Stationary_matrix3_6_7(my_stationary_io_o_Stationary_matrix3_6_7),
    .io_o_Stationary_matrix3_7_0(my_stationary_io_o_Stationary_matrix3_7_0),
    .io_o_Stationary_matrix3_7_1(my_stationary_io_o_Stationary_matrix3_7_1),
    .io_o_Stationary_matrix3_7_2(my_stationary_io_o_Stationary_matrix3_7_2),
    .io_o_Stationary_matrix3_7_3(my_stationary_io_o_Stationary_matrix3_7_3),
    .io_o_Stationary_matrix3_7_4(my_stationary_io_o_Stationary_matrix3_7_4),
    .io_o_Stationary_matrix3_7_5(my_stationary_io_o_Stationary_matrix3_7_5),
    .io_o_Stationary_matrix3_7_6(my_stationary_io_o_Stationary_matrix3_7_6),
    .io_o_Stationary_matrix3_7_7(my_stationary_io_o_Stationary_matrix3_7_7),
    .io_o_Stationary_matrix4_0_0(my_stationary_io_o_Stationary_matrix4_0_0),
    .io_o_Stationary_matrix4_0_1(my_stationary_io_o_Stationary_matrix4_0_1),
    .io_o_Stationary_matrix4_0_2(my_stationary_io_o_Stationary_matrix4_0_2),
    .io_o_Stationary_matrix4_0_3(my_stationary_io_o_Stationary_matrix4_0_3),
    .io_o_Stationary_matrix4_0_4(my_stationary_io_o_Stationary_matrix4_0_4),
    .io_o_Stationary_matrix4_0_5(my_stationary_io_o_Stationary_matrix4_0_5),
    .io_o_Stationary_matrix4_0_6(my_stationary_io_o_Stationary_matrix4_0_6),
    .io_o_Stationary_matrix4_0_7(my_stationary_io_o_Stationary_matrix4_0_7),
    .io_o_Stationary_matrix4_1_0(my_stationary_io_o_Stationary_matrix4_1_0),
    .io_o_Stationary_matrix4_1_1(my_stationary_io_o_Stationary_matrix4_1_1),
    .io_o_Stationary_matrix4_1_2(my_stationary_io_o_Stationary_matrix4_1_2),
    .io_o_Stationary_matrix4_1_3(my_stationary_io_o_Stationary_matrix4_1_3),
    .io_o_Stationary_matrix4_1_4(my_stationary_io_o_Stationary_matrix4_1_4),
    .io_o_Stationary_matrix4_1_5(my_stationary_io_o_Stationary_matrix4_1_5),
    .io_o_Stationary_matrix4_1_6(my_stationary_io_o_Stationary_matrix4_1_6),
    .io_o_Stationary_matrix4_1_7(my_stationary_io_o_Stationary_matrix4_1_7),
    .io_o_Stationary_matrix4_2_0(my_stationary_io_o_Stationary_matrix4_2_0),
    .io_o_Stationary_matrix4_2_1(my_stationary_io_o_Stationary_matrix4_2_1),
    .io_o_Stationary_matrix4_2_2(my_stationary_io_o_Stationary_matrix4_2_2),
    .io_o_Stationary_matrix4_2_3(my_stationary_io_o_Stationary_matrix4_2_3),
    .io_o_Stationary_matrix4_2_4(my_stationary_io_o_Stationary_matrix4_2_4),
    .io_o_Stationary_matrix4_2_5(my_stationary_io_o_Stationary_matrix4_2_5),
    .io_o_Stationary_matrix4_2_6(my_stationary_io_o_Stationary_matrix4_2_6),
    .io_o_Stationary_matrix4_2_7(my_stationary_io_o_Stationary_matrix4_2_7),
    .io_o_Stationary_matrix4_3_0(my_stationary_io_o_Stationary_matrix4_3_0),
    .io_o_Stationary_matrix4_3_1(my_stationary_io_o_Stationary_matrix4_3_1),
    .io_o_Stationary_matrix4_3_2(my_stationary_io_o_Stationary_matrix4_3_2),
    .io_o_Stationary_matrix4_3_3(my_stationary_io_o_Stationary_matrix4_3_3),
    .io_o_Stationary_matrix4_3_4(my_stationary_io_o_Stationary_matrix4_3_4),
    .io_o_Stationary_matrix4_3_5(my_stationary_io_o_Stationary_matrix4_3_5),
    .io_o_Stationary_matrix4_3_6(my_stationary_io_o_Stationary_matrix4_3_6),
    .io_o_Stationary_matrix4_3_7(my_stationary_io_o_Stationary_matrix4_3_7),
    .io_o_Stationary_matrix4_4_0(my_stationary_io_o_Stationary_matrix4_4_0),
    .io_o_Stationary_matrix4_4_1(my_stationary_io_o_Stationary_matrix4_4_1),
    .io_o_Stationary_matrix4_4_2(my_stationary_io_o_Stationary_matrix4_4_2),
    .io_o_Stationary_matrix4_4_3(my_stationary_io_o_Stationary_matrix4_4_3),
    .io_o_Stationary_matrix4_4_4(my_stationary_io_o_Stationary_matrix4_4_4),
    .io_o_Stationary_matrix4_4_5(my_stationary_io_o_Stationary_matrix4_4_5),
    .io_o_Stationary_matrix4_4_6(my_stationary_io_o_Stationary_matrix4_4_6),
    .io_o_Stationary_matrix4_4_7(my_stationary_io_o_Stationary_matrix4_4_7),
    .io_o_Stationary_matrix4_5_0(my_stationary_io_o_Stationary_matrix4_5_0),
    .io_o_Stationary_matrix4_5_1(my_stationary_io_o_Stationary_matrix4_5_1),
    .io_o_Stationary_matrix4_5_2(my_stationary_io_o_Stationary_matrix4_5_2),
    .io_o_Stationary_matrix4_5_3(my_stationary_io_o_Stationary_matrix4_5_3),
    .io_o_Stationary_matrix4_5_4(my_stationary_io_o_Stationary_matrix4_5_4),
    .io_o_Stationary_matrix4_5_5(my_stationary_io_o_Stationary_matrix4_5_5),
    .io_o_Stationary_matrix4_5_6(my_stationary_io_o_Stationary_matrix4_5_6),
    .io_o_Stationary_matrix4_5_7(my_stationary_io_o_Stationary_matrix4_5_7),
    .io_o_Stationary_matrix4_6_0(my_stationary_io_o_Stationary_matrix4_6_0),
    .io_o_Stationary_matrix4_6_1(my_stationary_io_o_Stationary_matrix4_6_1),
    .io_o_Stationary_matrix4_6_2(my_stationary_io_o_Stationary_matrix4_6_2),
    .io_o_Stationary_matrix4_6_3(my_stationary_io_o_Stationary_matrix4_6_3),
    .io_o_Stationary_matrix4_6_4(my_stationary_io_o_Stationary_matrix4_6_4),
    .io_o_Stationary_matrix4_6_5(my_stationary_io_o_Stationary_matrix4_6_5),
    .io_o_Stationary_matrix4_6_6(my_stationary_io_o_Stationary_matrix4_6_6),
    .io_o_Stationary_matrix4_6_7(my_stationary_io_o_Stationary_matrix4_6_7),
    .io_o_Stationary_matrix4_7_0(my_stationary_io_o_Stationary_matrix4_7_0),
    .io_o_Stationary_matrix4_7_1(my_stationary_io_o_Stationary_matrix4_7_1),
    .io_o_Stationary_matrix4_7_2(my_stationary_io_o_Stationary_matrix4_7_2),
    .io_o_Stationary_matrix4_7_3(my_stationary_io_o_Stationary_matrix4_7_3),
    .io_o_Stationary_matrix4_7_4(my_stationary_io_o_Stationary_matrix4_7_4),
    .io_o_Stationary_matrix4_7_5(my_stationary_io_o_Stationary_matrix4_7_5),
    .io_o_Stationary_matrix4_7_6(my_stationary_io_o_Stationary_matrix4_7_6),
    .io_o_Stationary_matrix4_7_7(my_stationary_io_o_Stationary_matrix4_7_7),
    .io_o_Stationary_matrix5_0_0(my_stationary_io_o_Stationary_matrix5_0_0),
    .io_o_Stationary_matrix5_0_1(my_stationary_io_o_Stationary_matrix5_0_1),
    .io_o_Stationary_matrix5_0_2(my_stationary_io_o_Stationary_matrix5_0_2),
    .io_o_Stationary_matrix5_0_3(my_stationary_io_o_Stationary_matrix5_0_3),
    .io_o_Stationary_matrix5_0_4(my_stationary_io_o_Stationary_matrix5_0_4),
    .io_o_Stationary_matrix5_0_5(my_stationary_io_o_Stationary_matrix5_0_5),
    .io_o_Stationary_matrix5_0_6(my_stationary_io_o_Stationary_matrix5_0_6),
    .io_o_Stationary_matrix5_0_7(my_stationary_io_o_Stationary_matrix5_0_7),
    .io_o_Stationary_matrix5_1_0(my_stationary_io_o_Stationary_matrix5_1_0),
    .io_o_Stationary_matrix5_1_1(my_stationary_io_o_Stationary_matrix5_1_1),
    .io_o_Stationary_matrix5_1_2(my_stationary_io_o_Stationary_matrix5_1_2),
    .io_o_Stationary_matrix5_1_3(my_stationary_io_o_Stationary_matrix5_1_3),
    .io_o_Stationary_matrix5_1_4(my_stationary_io_o_Stationary_matrix5_1_4),
    .io_o_Stationary_matrix5_1_5(my_stationary_io_o_Stationary_matrix5_1_5),
    .io_o_Stationary_matrix5_1_6(my_stationary_io_o_Stationary_matrix5_1_6),
    .io_o_Stationary_matrix5_1_7(my_stationary_io_o_Stationary_matrix5_1_7),
    .io_o_Stationary_matrix5_2_0(my_stationary_io_o_Stationary_matrix5_2_0),
    .io_o_Stationary_matrix5_2_1(my_stationary_io_o_Stationary_matrix5_2_1),
    .io_o_Stationary_matrix5_2_2(my_stationary_io_o_Stationary_matrix5_2_2),
    .io_o_Stationary_matrix5_2_3(my_stationary_io_o_Stationary_matrix5_2_3),
    .io_o_Stationary_matrix5_2_4(my_stationary_io_o_Stationary_matrix5_2_4),
    .io_o_Stationary_matrix5_2_5(my_stationary_io_o_Stationary_matrix5_2_5),
    .io_o_Stationary_matrix5_2_6(my_stationary_io_o_Stationary_matrix5_2_6),
    .io_o_Stationary_matrix5_2_7(my_stationary_io_o_Stationary_matrix5_2_7),
    .io_o_Stationary_matrix5_3_0(my_stationary_io_o_Stationary_matrix5_3_0),
    .io_o_Stationary_matrix5_3_1(my_stationary_io_o_Stationary_matrix5_3_1),
    .io_o_Stationary_matrix5_3_2(my_stationary_io_o_Stationary_matrix5_3_2),
    .io_o_Stationary_matrix5_3_3(my_stationary_io_o_Stationary_matrix5_3_3),
    .io_o_Stationary_matrix5_3_4(my_stationary_io_o_Stationary_matrix5_3_4),
    .io_o_Stationary_matrix5_3_5(my_stationary_io_o_Stationary_matrix5_3_5),
    .io_o_Stationary_matrix5_3_6(my_stationary_io_o_Stationary_matrix5_3_6),
    .io_o_Stationary_matrix5_3_7(my_stationary_io_o_Stationary_matrix5_3_7),
    .io_o_Stationary_matrix5_4_0(my_stationary_io_o_Stationary_matrix5_4_0),
    .io_o_Stationary_matrix5_4_1(my_stationary_io_o_Stationary_matrix5_4_1),
    .io_o_Stationary_matrix5_4_2(my_stationary_io_o_Stationary_matrix5_4_2),
    .io_o_Stationary_matrix5_4_3(my_stationary_io_o_Stationary_matrix5_4_3),
    .io_o_Stationary_matrix5_4_4(my_stationary_io_o_Stationary_matrix5_4_4),
    .io_o_Stationary_matrix5_4_5(my_stationary_io_o_Stationary_matrix5_4_5),
    .io_o_Stationary_matrix5_4_6(my_stationary_io_o_Stationary_matrix5_4_6),
    .io_o_Stationary_matrix5_4_7(my_stationary_io_o_Stationary_matrix5_4_7),
    .io_o_Stationary_matrix5_5_0(my_stationary_io_o_Stationary_matrix5_5_0),
    .io_o_Stationary_matrix5_5_1(my_stationary_io_o_Stationary_matrix5_5_1),
    .io_o_Stationary_matrix5_5_2(my_stationary_io_o_Stationary_matrix5_5_2),
    .io_o_Stationary_matrix5_5_3(my_stationary_io_o_Stationary_matrix5_5_3),
    .io_o_Stationary_matrix5_5_4(my_stationary_io_o_Stationary_matrix5_5_4),
    .io_o_Stationary_matrix5_5_5(my_stationary_io_o_Stationary_matrix5_5_5),
    .io_o_Stationary_matrix5_5_6(my_stationary_io_o_Stationary_matrix5_5_6),
    .io_o_Stationary_matrix5_5_7(my_stationary_io_o_Stationary_matrix5_5_7),
    .io_o_Stationary_matrix5_6_0(my_stationary_io_o_Stationary_matrix5_6_0),
    .io_o_Stationary_matrix5_6_1(my_stationary_io_o_Stationary_matrix5_6_1),
    .io_o_Stationary_matrix5_6_2(my_stationary_io_o_Stationary_matrix5_6_2),
    .io_o_Stationary_matrix5_6_3(my_stationary_io_o_Stationary_matrix5_6_3),
    .io_o_Stationary_matrix5_6_4(my_stationary_io_o_Stationary_matrix5_6_4),
    .io_o_Stationary_matrix5_6_5(my_stationary_io_o_Stationary_matrix5_6_5),
    .io_o_Stationary_matrix5_6_6(my_stationary_io_o_Stationary_matrix5_6_6),
    .io_o_Stationary_matrix5_6_7(my_stationary_io_o_Stationary_matrix5_6_7),
    .io_o_Stationary_matrix5_7_0(my_stationary_io_o_Stationary_matrix5_7_0),
    .io_o_Stationary_matrix5_7_1(my_stationary_io_o_Stationary_matrix5_7_1),
    .io_o_Stationary_matrix5_7_2(my_stationary_io_o_Stationary_matrix5_7_2),
    .io_o_Stationary_matrix5_7_3(my_stationary_io_o_Stationary_matrix5_7_3),
    .io_o_Stationary_matrix5_7_4(my_stationary_io_o_Stationary_matrix5_7_4),
    .io_o_Stationary_matrix5_7_5(my_stationary_io_o_Stationary_matrix5_7_5),
    .io_o_Stationary_matrix5_7_6(my_stationary_io_o_Stationary_matrix5_7_6),
    .io_o_Stationary_matrix5_7_7(my_stationary_io_o_Stationary_matrix5_7_7),
    .io_o_Stationary_matrix6_0_0(my_stationary_io_o_Stationary_matrix6_0_0),
    .io_o_Stationary_matrix6_0_1(my_stationary_io_o_Stationary_matrix6_0_1),
    .io_o_Stationary_matrix6_0_2(my_stationary_io_o_Stationary_matrix6_0_2),
    .io_o_Stationary_matrix6_0_3(my_stationary_io_o_Stationary_matrix6_0_3),
    .io_o_Stationary_matrix6_0_4(my_stationary_io_o_Stationary_matrix6_0_4),
    .io_o_Stationary_matrix6_0_5(my_stationary_io_o_Stationary_matrix6_0_5),
    .io_o_Stationary_matrix6_0_6(my_stationary_io_o_Stationary_matrix6_0_6),
    .io_o_Stationary_matrix6_0_7(my_stationary_io_o_Stationary_matrix6_0_7),
    .io_o_Stationary_matrix6_1_0(my_stationary_io_o_Stationary_matrix6_1_0),
    .io_o_Stationary_matrix6_1_1(my_stationary_io_o_Stationary_matrix6_1_1),
    .io_o_Stationary_matrix6_1_2(my_stationary_io_o_Stationary_matrix6_1_2),
    .io_o_Stationary_matrix6_1_3(my_stationary_io_o_Stationary_matrix6_1_3),
    .io_o_Stationary_matrix6_1_4(my_stationary_io_o_Stationary_matrix6_1_4),
    .io_o_Stationary_matrix6_1_5(my_stationary_io_o_Stationary_matrix6_1_5),
    .io_o_Stationary_matrix6_1_6(my_stationary_io_o_Stationary_matrix6_1_6),
    .io_o_Stationary_matrix6_1_7(my_stationary_io_o_Stationary_matrix6_1_7),
    .io_o_Stationary_matrix6_2_0(my_stationary_io_o_Stationary_matrix6_2_0),
    .io_o_Stationary_matrix6_2_1(my_stationary_io_o_Stationary_matrix6_2_1),
    .io_o_Stationary_matrix6_2_2(my_stationary_io_o_Stationary_matrix6_2_2),
    .io_o_Stationary_matrix6_2_3(my_stationary_io_o_Stationary_matrix6_2_3),
    .io_o_Stationary_matrix6_2_4(my_stationary_io_o_Stationary_matrix6_2_4),
    .io_o_Stationary_matrix6_2_5(my_stationary_io_o_Stationary_matrix6_2_5),
    .io_o_Stationary_matrix6_2_6(my_stationary_io_o_Stationary_matrix6_2_6),
    .io_o_Stationary_matrix6_2_7(my_stationary_io_o_Stationary_matrix6_2_7),
    .io_o_Stationary_matrix6_3_0(my_stationary_io_o_Stationary_matrix6_3_0),
    .io_o_Stationary_matrix6_3_1(my_stationary_io_o_Stationary_matrix6_3_1),
    .io_o_Stationary_matrix6_3_2(my_stationary_io_o_Stationary_matrix6_3_2),
    .io_o_Stationary_matrix6_3_3(my_stationary_io_o_Stationary_matrix6_3_3),
    .io_o_Stationary_matrix6_3_4(my_stationary_io_o_Stationary_matrix6_3_4),
    .io_o_Stationary_matrix6_3_5(my_stationary_io_o_Stationary_matrix6_3_5),
    .io_o_Stationary_matrix6_3_6(my_stationary_io_o_Stationary_matrix6_3_6),
    .io_o_Stationary_matrix6_3_7(my_stationary_io_o_Stationary_matrix6_3_7),
    .io_o_Stationary_matrix6_4_0(my_stationary_io_o_Stationary_matrix6_4_0),
    .io_o_Stationary_matrix6_4_1(my_stationary_io_o_Stationary_matrix6_4_1),
    .io_o_Stationary_matrix6_4_2(my_stationary_io_o_Stationary_matrix6_4_2),
    .io_o_Stationary_matrix6_4_3(my_stationary_io_o_Stationary_matrix6_4_3),
    .io_o_Stationary_matrix6_4_4(my_stationary_io_o_Stationary_matrix6_4_4),
    .io_o_Stationary_matrix6_4_5(my_stationary_io_o_Stationary_matrix6_4_5),
    .io_o_Stationary_matrix6_4_6(my_stationary_io_o_Stationary_matrix6_4_6),
    .io_o_Stationary_matrix6_4_7(my_stationary_io_o_Stationary_matrix6_4_7),
    .io_o_Stationary_matrix6_5_0(my_stationary_io_o_Stationary_matrix6_5_0),
    .io_o_Stationary_matrix6_5_1(my_stationary_io_o_Stationary_matrix6_5_1),
    .io_o_Stationary_matrix6_5_2(my_stationary_io_o_Stationary_matrix6_5_2),
    .io_o_Stationary_matrix6_5_3(my_stationary_io_o_Stationary_matrix6_5_3),
    .io_o_Stationary_matrix6_5_4(my_stationary_io_o_Stationary_matrix6_5_4),
    .io_o_Stationary_matrix6_5_5(my_stationary_io_o_Stationary_matrix6_5_5),
    .io_o_Stationary_matrix6_5_6(my_stationary_io_o_Stationary_matrix6_5_6),
    .io_o_Stationary_matrix6_5_7(my_stationary_io_o_Stationary_matrix6_5_7),
    .io_o_Stationary_matrix6_6_0(my_stationary_io_o_Stationary_matrix6_6_0),
    .io_o_Stationary_matrix6_6_1(my_stationary_io_o_Stationary_matrix6_6_1),
    .io_o_Stationary_matrix6_6_2(my_stationary_io_o_Stationary_matrix6_6_2),
    .io_o_Stationary_matrix6_6_3(my_stationary_io_o_Stationary_matrix6_6_3),
    .io_o_Stationary_matrix6_6_4(my_stationary_io_o_Stationary_matrix6_6_4),
    .io_o_Stationary_matrix6_6_5(my_stationary_io_o_Stationary_matrix6_6_5),
    .io_o_Stationary_matrix6_6_6(my_stationary_io_o_Stationary_matrix6_6_6),
    .io_o_Stationary_matrix6_6_7(my_stationary_io_o_Stationary_matrix6_6_7),
    .io_o_Stationary_matrix6_7_0(my_stationary_io_o_Stationary_matrix6_7_0),
    .io_o_Stationary_matrix6_7_1(my_stationary_io_o_Stationary_matrix6_7_1),
    .io_o_Stationary_matrix6_7_2(my_stationary_io_o_Stationary_matrix6_7_2),
    .io_o_Stationary_matrix6_7_3(my_stationary_io_o_Stationary_matrix6_7_3),
    .io_o_Stationary_matrix6_7_4(my_stationary_io_o_Stationary_matrix6_7_4),
    .io_o_Stationary_matrix6_7_5(my_stationary_io_o_Stationary_matrix6_7_5),
    .io_o_Stationary_matrix6_7_6(my_stationary_io_o_Stationary_matrix6_7_6),
    .io_o_Stationary_matrix6_7_7(my_stationary_io_o_Stationary_matrix6_7_7),
    .io_o_Stationary_matrix7_0_0(my_stationary_io_o_Stationary_matrix7_0_0),
    .io_o_Stationary_matrix7_0_1(my_stationary_io_o_Stationary_matrix7_0_1),
    .io_o_Stationary_matrix7_0_2(my_stationary_io_o_Stationary_matrix7_0_2),
    .io_o_Stationary_matrix7_0_3(my_stationary_io_o_Stationary_matrix7_0_3),
    .io_o_Stationary_matrix7_0_4(my_stationary_io_o_Stationary_matrix7_0_4),
    .io_o_Stationary_matrix7_0_5(my_stationary_io_o_Stationary_matrix7_0_5),
    .io_o_Stationary_matrix7_0_6(my_stationary_io_o_Stationary_matrix7_0_6),
    .io_o_Stationary_matrix7_0_7(my_stationary_io_o_Stationary_matrix7_0_7),
    .io_o_Stationary_matrix7_1_0(my_stationary_io_o_Stationary_matrix7_1_0),
    .io_o_Stationary_matrix7_1_1(my_stationary_io_o_Stationary_matrix7_1_1),
    .io_o_Stationary_matrix7_1_2(my_stationary_io_o_Stationary_matrix7_1_2),
    .io_o_Stationary_matrix7_1_3(my_stationary_io_o_Stationary_matrix7_1_3),
    .io_o_Stationary_matrix7_1_4(my_stationary_io_o_Stationary_matrix7_1_4),
    .io_o_Stationary_matrix7_1_5(my_stationary_io_o_Stationary_matrix7_1_5),
    .io_o_Stationary_matrix7_1_6(my_stationary_io_o_Stationary_matrix7_1_6),
    .io_o_Stationary_matrix7_1_7(my_stationary_io_o_Stationary_matrix7_1_7),
    .io_o_Stationary_matrix7_2_0(my_stationary_io_o_Stationary_matrix7_2_0),
    .io_o_Stationary_matrix7_2_1(my_stationary_io_o_Stationary_matrix7_2_1),
    .io_o_Stationary_matrix7_2_2(my_stationary_io_o_Stationary_matrix7_2_2),
    .io_o_Stationary_matrix7_2_3(my_stationary_io_o_Stationary_matrix7_2_3),
    .io_o_Stationary_matrix7_2_4(my_stationary_io_o_Stationary_matrix7_2_4),
    .io_o_Stationary_matrix7_2_5(my_stationary_io_o_Stationary_matrix7_2_5),
    .io_o_Stationary_matrix7_2_6(my_stationary_io_o_Stationary_matrix7_2_6),
    .io_o_Stationary_matrix7_2_7(my_stationary_io_o_Stationary_matrix7_2_7),
    .io_o_Stationary_matrix7_3_0(my_stationary_io_o_Stationary_matrix7_3_0),
    .io_o_Stationary_matrix7_3_1(my_stationary_io_o_Stationary_matrix7_3_1),
    .io_o_Stationary_matrix7_3_2(my_stationary_io_o_Stationary_matrix7_3_2),
    .io_o_Stationary_matrix7_3_3(my_stationary_io_o_Stationary_matrix7_3_3),
    .io_o_Stationary_matrix7_3_4(my_stationary_io_o_Stationary_matrix7_3_4),
    .io_o_Stationary_matrix7_3_5(my_stationary_io_o_Stationary_matrix7_3_5),
    .io_o_Stationary_matrix7_3_6(my_stationary_io_o_Stationary_matrix7_3_6),
    .io_o_Stationary_matrix7_3_7(my_stationary_io_o_Stationary_matrix7_3_7),
    .io_o_Stationary_matrix7_4_0(my_stationary_io_o_Stationary_matrix7_4_0),
    .io_o_Stationary_matrix7_4_1(my_stationary_io_o_Stationary_matrix7_4_1),
    .io_o_Stationary_matrix7_4_2(my_stationary_io_o_Stationary_matrix7_4_2),
    .io_o_Stationary_matrix7_4_3(my_stationary_io_o_Stationary_matrix7_4_3),
    .io_o_Stationary_matrix7_4_4(my_stationary_io_o_Stationary_matrix7_4_4),
    .io_o_Stationary_matrix7_4_5(my_stationary_io_o_Stationary_matrix7_4_5),
    .io_o_Stationary_matrix7_4_6(my_stationary_io_o_Stationary_matrix7_4_6),
    .io_o_Stationary_matrix7_4_7(my_stationary_io_o_Stationary_matrix7_4_7),
    .io_o_Stationary_matrix7_5_0(my_stationary_io_o_Stationary_matrix7_5_0),
    .io_o_Stationary_matrix7_5_1(my_stationary_io_o_Stationary_matrix7_5_1),
    .io_o_Stationary_matrix7_5_2(my_stationary_io_o_Stationary_matrix7_5_2),
    .io_o_Stationary_matrix7_5_3(my_stationary_io_o_Stationary_matrix7_5_3),
    .io_o_Stationary_matrix7_5_4(my_stationary_io_o_Stationary_matrix7_5_4),
    .io_o_Stationary_matrix7_5_5(my_stationary_io_o_Stationary_matrix7_5_5),
    .io_o_Stationary_matrix7_5_6(my_stationary_io_o_Stationary_matrix7_5_6),
    .io_o_Stationary_matrix7_5_7(my_stationary_io_o_Stationary_matrix7_5_7),
    .io_o_Stationary_matrix7_6_0(my_stationary_io_o_Stationary_matrix7_6_0),
    .io_o_Stationary_matrix7_6_1(my_stationary_io_o_Stationary_matrix7_6_1),
    .io_o_Stationary_matrix7_6_2(my_stationary_io_o_Stationary_matrix7_6_2),
    .io_o_Stationary_matrix7_6_3(my_stationary_io_o_Stationary_matrix7_6_3),
    .io_o_Stationary_matrix7_6_4(my_stationary_io_o_Stationary_matrix7_6_4),
    .io_o_Stationary_matrix7_6_5(my_stationary_io_o_Stationary_matrix7_6_5),
    .io_o_Stationary_matrix7_6_6(my_stationary_io_o_Stationary_matrix7_6_6),
    .io_o_Stationary_matrix7_6_7(my_stationary_io_o_Stationary_matrix7_6_7),
    .io_o_Stationary_matrix7_7_0(my_stationary_io_o_Stationary_matrix7_7_0),
    .io_o_Stationary_matrix7_7_1(my_stationary_io_o_Stationary_matrix7_7_1),
    .io_o_Stationary_matrix7_7_2(my_stationary_io_o_Stationary_matrix7_7_2),
    .io_o_Stationary_matrix7_7_3(my_stationary_io_o_Stationary_matrix7_7_3),
    .io_o_Stationary_matrix7_7_4(my_stationary_io_o_Stationary_matrix7_7_4),
    .io_o_Stationary_matrix7_7_5(my_stationary_io_o_Stationary_matrix7_7_5),
    .io_o_Stationary_matrix7_7_6(my_stationary_io_o_Stationary_matrix7_7_6),
    .io_o_Stationary_matrix7_7_7(my_stationary_io_o_Stationary_matrix7_7_7),
    .io_o_Stationary_matrix8_0_0(my_stationary_io_o_Stationary_matrix8_0_0),
    .io_o_Stationary_matrix8_0_1(my_stationary_io_o_Stationary_matrix8_0_1),
    .io_o_Stationary_matrix8_0_2(my_stationary_io_o_Stationary_matrix8_0_2),
    .io_o_Stationary_matrix8_0_3(my_stationary_io_o_Stationary_matrix8_0_3),
    .io_o_Stationary_matrix8_0_4(my_stationary_io_o_Stationary_matrix8_0_4),
    .io_o_Stationary_matrix8_0_5(my_stationary_io_o_Stationary_matrix8_0_5),
    .io_o_Stationary_matrix8_0_6(my_stationary_io_o_Stationary_matrix8_0_6),
    .io_o_Stationary_matrix8_0_7(my_stationary_io_o_Stationary_matrix8_0_7),
    .io_o_Stationary_matrix8_1_0(my_stationary_io_o_Stationary_matrix8_1_0),
    .io_o_Stationary_matrix8_1_1(my_stationary_io_o_Stationary_matrix8_1_1),
    .io_o_Stationary_matrix8_1_2(my_stationary_io_o_Stationary_matrix8_1_2),
    .io_o_Stationary_matrix8_1_3(my_stationary_io_o_Stationary_matrix8_1_3),
    .io_o_Stationary_matrix8_1_4(my_stationary_io_o_Stationary_matrix8_1_4),
    .io_o_Stationary_matrix8_1_5(my_stationary_io_o_Stationary_matrix8_1_5),
    .io_o_Stationary_matrix8_1_6(my_stationary_io_o_Stationary_matrix8_1_6),
    .io_o_Stationary_matrix8_1_7(my_stationary_io_o_Stationary_matrix8_1_7),
    .io_o_Stationary_matrix8_2_0(my_stationary_io_o_Stationary_matrix8_2_0),
    .io_o_Stationary_matrix8_2_1(my_stationary_io_o_Stationary_matrix8_2_1),
    .io_o_Stationary_matrix8_2_2(my_stationary_io_o_Stationary_matrix8_2_2),
    .io_o_Stationary_matrix8_2_3(my_stationary_io_o_Stationary_matrix8_2_3),
    .io_o_Stationary_matrix8_2_4(my_stationary_io_o_Stationary_matrix8_2_4),
    .io_o_Stationary_matrix8_2_5(my_stationary_io_o_Stationary_matrix8_2_5),
    .io_o_Stationary_matrix8_2_6(my_stationary_io_o_Stationary_matrix8_2_6),
    .io_o_Stationary_matrix8_2_7(my_stationary_io_o_Stationary_matrix8_2_7),
    .io_o_Stationary_matrix8_3_0(my_stationary_io_o_Stationary_matrix8_3_0),
    .io_o_Stationary_matrix8_3_1(my_stationary_io_o_Stationary_matrix8_3_1),
    .io_o_Stationary_matrix8_3_2(my_stationary_io_o_Stationary_matrix8_3_2),
    .io_o_Stationary_matrix8_3_3(my_stationary_io_o_Stationary_matrix8_3_3),
    .io_o_Stationary_matrix8_3_4(my_stationary_io_o_Stationary_matrix8_3_4),
    .io_o_Stationary_matrix8_3_5(my_stationary_io_o_Stationary_matrix8_3_5),
    .io_o_Stationary_matrix8_3_6(my_stationary_io_o_Stationary_matrix8_3_6),
    .io_o_Stationary_matrix8_3_7(my_stationary_io_o_Stationary_matrix8_3_7),
    .io_o_Stationary_matrix8_4_0(my_stationary_io_o_Stationary_matrix8_4_0),
    .io_o_Stationary_matrix8_4_1(my_stationary_io_o_Stationary_matrix8_4_1),
    .io_o_Stationary_matrix8_4_2(my_stationary_io_o_Stationary_matrix8_4_2),
    .io_o_Stationary_matrix8_4_3(my_stationary_io_o_Stationary_matrix8_4_3),
    .io_o_Stationary_matrix8_4_4(my_stationary_io_o_Stationary_matrix8_4_4),
    .io_o_Stationary_matrix8_4_5(my_stationary_io_o_Stationary_matrix8_4_5),
    .io_o_Stationary_matrix8_4_6(my_stationary_io_o_Stationary_matrix8_4_6),
    .io_o_Stationary_matrix8_4_7(my_stationary_io_o_Stationary_matrix8_4_7),
    .io_o_Stationary_matrix8_5_0(my_stationary_io_o_Stationary_matrix8_5_0),
    .io_o_Stationary_matrix8_5_1(my_stationary_io_o_Stationary_matrix8_5_1),
    .io_o_Stationary_matrix8_5_2(my_stationary_io_o_Stationary_matrix8_5_2),
    .io_o_Stationary_matrix8_5_3(my_stationary_io_o_Stationary_matrix8_5_3),
    .io_o_Stationary_matrix8_5_4(my_stationary_io_o_Stationary_matrix8_5_4),
    .io_o_Stationary_matrix8_5_5(my_stationary_io_o_Stationary_matrix8_5_5),
    .io_o_Stationary_matrix8_5_6(my_stationary_io_o_Stationary_matrix8_5_6),
    .io_o_Stationary_matrix8_5_7(my_stationary_io_o_Stationary_matrix8_5_7),
    .io_o_Stationary_matrix8_6_0(my_stationary_io_o_Stationary_matrix8_6_0),
    .io_o_Stationary_matrix8_6_1(my_stationary_io_o_Stationary_matrix8_6_1),
    .io_o_Stationary_matrix8_6_2(my_stationary_io_o_Stationary_matrix8_6_2),
    .io_o_Stationary_matrix8_6_3(my_stationary_io_o_Stationary_matrix8_6_3),
    .io_o_Stationary_matrix8_6_4(my_stationary_io_o_Stationary_matrix8_6_4),
    .io_o_Stationary_matrix8_6_5(my_stationary_io_o_Stationary_matrix8_6_5),
    .io_o_Stationary_matrix8_6_6(my_stationary_io_o_Stationary_matrix8_6_6),
    .io_o_Stationary_matrix8_6_7(my_stationary_io_o_Stationary_matrix8_6_7),
    .io_o_Stationary_matrix8_7_0(my_stationary_io_o_Stationary_matrix8_7_0),
    .io_o_Stationary_matrix8_7_1(my_stationary_io_o_Stationary_matrix8_7_1),
    .io_o_Stationary_matrix8_7_2(my_stationary_io_o_Stationary_matrix8_7_2),
    .io_o_Stationary_matrix8_7_3(my_stationary_io_o_Stationary_matrix8_7_3),
    .io_o_Stationary_matrix8_7_4(my_stationary_io_o_Stationary_matrix8_7_4),
    .io_o_Stationary_matrix8_7_5(my_stationary_io_o_Stationary_matrix8_7_5),
    .io_o_Stationary_matrix8_7_6(my_stationary_io_o_Stationary_matrix8_7_6),
    .io_o_Stationary_matrix8_7_7(my_stationary_io_o_Stationary_matrix8_7_7)
  );
  ivncontrol4 my_ivn1 ( // @[ivntop.scala 69:24]
    .clock(my_ivn1_clock),
    .reset(my_ivn1_reset),
    .io_Stationary_matrix_0_0(my_ivn1_io_Stationary_matrix_0_0),
    .io_Stationary_matrix_0_1(my_ivn1_io_Stationary_matrix_0_1),
    .io_Stationary_matrix_0_2(my_ivn1_io_Stationary_matrix_0_2),
    .io_Stationary_matrix_0_3(my_ivn1_io_Stationary_matrix_0_3),
    .io_Stationary_matrix_0_4(my_ivn1_io_Stationary_matrix_0_4),
    .io_Stationary_matrix_0_5(my_ivn1_io_Stationary_matrix_0_5),
    .io_Stationary_matrix_0_6(my_ivn1_io_Stationary_matrix_0_6),
    .io_Stationary_matrix_0_7(my_ivn1_io_Stationary_matrix_0_7),
    .io_Stationary_matrix_1_0(my_ivn1_io_Stationary_matrix_1_0),
    .io_Stationary_matrix_1_1(my_ivn1_io_Stationary_matrix_1_1),
    .io_Stationary_matrix_1_2(my_ivn1_io_Stationary_matrix_1_2),
    .io_Stationary_matrix_1_3(my_ivn1_io_Stationary_matrix_1_3),
    .io_Stationary_matrix_1_4(my_ivn1_io_Stationary_matrix_1_4),
    .io_Stationary_matrix_1_5(my_ivn1_io_Stationary_matrix_1_5),
    .io_Stationary_matrix_1_6(my_ivn1_io_Stationary_matrix_1_6),
    .io_Stationary_matrix_1_7(my_ivn1_io_Stationary_matrix_1_7),
    .io_Stationary_matrix_2_0(my_ivn1_io_Stationary_matrix_2_0),
    .io_Stationary_matrix_2_1(my_ivn1_io_Stationary_matrix_2_1),
    .io_Stationary_matrix_2_2(my_ivn1_io_Stationary_matrix_2_2),
    .io_Stationary_matrix_2_3(my_ivn1_io_Stationary_matrix_2_3),
    .io_Stationary_matrix_2_4(my_ivn1_io_Stationary_matrix_2_4),
    .io_Stationary_matrix_2_5(my_ivn1_io_Stationary_matrix_2_5),
    .io_Stationary_matrix_2_6(my_ivn1_io_Stationary_matrix_2_6),
    .io_Stationary_matrix_2_7(my_ivn1_io_Stationary_matrix_2_7),
    .io_Stationary_matrix_3_0(my_ivn1_io_Stationary_matrix_3_0),
    .io_Stationary_matrix_3_1(my_ivn1_io_Stationary_matrix_3_1),
    .io_Stationary_matrix_3_2(my_ivn1_io_Stationary_matrix_3_2),
    .io_Stationary_matrix_3_3(my_ivn1_io_Stationary_matrix_3_3),
    .io_Stationary_matrix_3_4(my_ivn1_io_Stationary_matrix_3_4),
    .io_Stationary_matrix_3_5(my_ivn1_io_Stationary_matrix_3_5),
    .io_Stationary_matrix_3_6(my_ivn1_io_Stationary_matrix_3_6),
    .io_Stationary_matrix_3_7(my_ivn1_io_Stationary_matrix_3_7),
    .io_Stationary_matrix_4_0(my_ivn1_io_Stationary_matrix_4_0),
    .io_Stationary_matrix_4_1(my_ivn1_io_Stationary_matrix_4_1),
    .io_Stationary_matrix_4_2(my_ivn1_io_Stationary_matrix_4_2),
    .io_Stationary_matrix_4_3(my_ivn1_io_Stationary_matrix_4_3),
    .io_Stationary_matrix_4_4(my_ivn1_io_Stationary_matrix_4_4),
    .io_Stationary_matrix_4_5(my_ivn1_io_Stationary_matrix_4_5),
    .io_Stationary_matrix_4_6(my_ivn1_io_Stationary_matrix_4_6),
    .io_Stationary_matrix_4_7(my_ivn1_io_Stationary_matrix_4_7),
    .io_Stationary_matrix_5_0(my_ivn1_io_Stationary_matrix_5_0),
    .io_Stationary_matrix_5_1(my_ivn1_io_Stationary_matrix_5_1),
    .io_Stationary_matrix_5_2(my_ivn1_io_Stationary_matrix_5_2),
    .io_Stationary_matrix_5_3(my_ivn1_io_Stationary_matrix_5_3),
    .io_Stationary_matrix_5_4(my_ivn1_io_Stationary_matrix_5_4),
    .io_Stationary_matrix_5_5(my_ivn1_io_Stationary_matrix_5_5),
    .io_Stationary_matrix_5_6(my_ivn1_io_Stationary_matrix_5_6),
    .io_Stationary_matrix_5_7(my_ivn1_io_Stationary_matrix_5_7),
    .io_Stationary_matrix_6_0(my_ivn1_io_Stationary_matrix_6_0),
    .io_Stationary_matrix_6_1(my_ivn1_io_Stationary_matrix_6_1),
    .io_Stationary_matrix_6_2(my_ivn1_io_Stationary_matrix_6_2),
    .io_Stationary_matrix_6_3(my_ivn1_io_Stationary_matrix_6_3),
    .io_Stationary_matrix_6_4(my_ivn1_io_Stationary_matrix_6_4),
    .io_Stationary_matrix_6_5(my_ivn1_io_Stationary_matrix_6_5),
    .io_Stationary_matrix_6_6(my_ivn1_io_Stationary_matrix_6_6),
    .io_Stationary_matrix_6_7(my_ivn1_io_Stationary_matrix_6_7),
    .io_Stationary_matrix_7_0(my_ivn1_io_Stationary_matrix_7_0),
    .io_Stationary_matrix_7_1(my_ivn1_io_Stationary_matrix_7_1),
    .io_Stationary_matrix_7_2(my_ivn1_io_Stationary_matrix_7_2),
    .io_Stationary_matrix_7_3(my_ivn1_io_Stationary_matrix_7_3),
    .io_Stationary_matrix_7_4(my_ivn1_io_Stationary_matrix_7_4),
    .io_Stationary_matrix_7_5(my_ivn1_io_Stationary_matrix_7_5),
    .io_Stationary_matrix_7_6(my_ivn1_io_Stationary_matrix_7_6),
    .io_Stationary_matrix_7_7(my_ivn1_io_Stationary_matrix_7_7),
    .io_o_vn_0(my_ivn1_io_o_vn_0),
    .io_o_vn_1(my_ivn1_io_o_vn_1),
    .io_o_vn_2(my_ivn1_io_o_vn_2),
    .io_o_vn_3(my_ivn1_io_o_vn_3),
    .io_o_vn2_0(my_ivn1_io_o_vn2_0),
    .io_o_vn2_1(my_ivn1_io_o_vn2_1),
    .io_o_vn2_2(my_ivn1_io_o_vn2_2),
    .io_o_vn2_3(my_ivn1_io_o_vn2_3),
    .io_ProcessValid(my_ivn1_io_ProcessValid),
    .io_validpin(my_ivn1_io_validpin)
  );
  ivncontrol4_1 my_ivn2 ( // @[ivntop.scala 78:24]
    .clock(my_ivn2_clock),
    .reset(my_ivn2_reset),
    .io_Stationary_matrix_0_0(my_ivn2_io_Stationary_matrix_0_0),
    .io_Stationary_matrix_0_1(my_ivn2_io_Stationary_matrix_0_1),
    .io_Stationary_matrix_0_2(my_ivn2_io_Stationary_matrix_0_2),
    .io_Stationary_matrix_0_3(my_ivn2_io_Stationary_matrix_0_3),
    .io_Stationary_matrix_0_4(my_ivn2_io_Stationary_matrix_0_4),
    .io_Stationary_matrix_0_5(my_ivn2_io_Stationary_matrix_0_5),
    .io_Stationary_matrix_0_6(my_ivn2_io_Stationary_matrix_0_6),
    .io_Stationary_matrix_0_7(my_ivn2_io_Stationary_matrix_0_7),
    .io_Stationary_matrix_1_0(my_ivn2_io_Stationary_matrix_1_0),
    .io_Stationary_matrix_1_1(my_ivn2_io_Stationary_matrix_1_1),
    .io_Stationary_matrix_1_2(my_ivn2_io_Stationary_matrix_1_2),
    .io_Stationary_matrix_1_3(my_ivn2_io_Stationary_matrix_1_3),
    .io_Stationary_matrix_1_4(my_ivn2_io_Stationary_matrix_1_4),
    .io_Stationary_matrix_1_5(my_ivn2_io_Stationary_matrix_1_5),
    .io_Stationary_matrix_1_6(my_ivn2_io_Stationary_matrix_1_6),
    .io_Stationary_matrix_1_7(my_ivn2_io_Stationary_matrix_1_7),
    .io_Stationary_matrix_2_0(my_ivn2_io_Stationary_matrix_2_0),
    .io_Stationary_matrix_2_1(my_ivn2_io_Stationary_matrix_2_1),
    .io_Stationary_matrix_2_2(my_ivn2_io_Stationary_matrix_2_2),
    .io_Stationary_matrix_2_3(my_ivn2_io_Stationary_matrix_2_3),
    .io_Stationary_matrix_2_4(my_ivn2_io_Stationary_matrix_2_4),
    .io_Stationary_matrix_2_5(my_ivn2_io_Stationary_matrix_2_5),
    .io_Stationary_matrix_2_6(my_ivn2_io_Stationary_matrix_2_6),
    .io_Stationary_matrix_2_7(my_ivn2_io_Stationary_matrix_2_7),
    .io_Stationary_matrix_3_0(my_ivn2_io_Stationary_matrix_3_0),
    .io_Stationary_matrix_3_1(my_ivn2_io_Stationary_matrix_3_1),
    .io_Stationary_matrix_3_2(my_ivn2_io_Stationary_matrix_3_2),
    .io_Stationary_matrix_3_3(my_ivn2_io_Stationary_matrix_3_3),
    .io_Stationary_matrix_3_4(my_ivn2_io_Stationary_matrix_3_4),
    .io_Stationary_matrix_3_5(my_ivn2_io_Stationary_matrix_3_5),
    .io_Stationary_matrix_3_6(my_ivn2_io_Stationary_matrix_3_6),
    .io_Stationary_matrix_3_7(my_ivn2_io_Stationary_matrix_3_7),
    .io_Stationary_matrix_4_0(my_ivn2_io_Stationary_matrix_4_0),
    .io_Stationary_matrix_4_1(my_ivn2_io_Stationary_matrix_4_1),
    .io_Stationary_matrix_4_2(my_ivn2_io_Stationary_matrix_4_2),
    .io_Stationary_matrix_4_3(my_ivn2_io_Stationary_matrix_4_3),
    .io_Stationary_matrix_4_4(my_ivn2_io_Stationary_matrix_4_4),
    .io_Stationary_matrix_4_5(my_ivn2_io_Stationary_matrix_4_5),
    .io_Stationary_matrix_4_6(my_ivn2_io_Stationary_matrix_4_6),
    .io_Stationary_matrix_4_7(my_ivn2_io_Stationary_matrix_4_7),
    .io_Stationary_matrix_5_0(my_ivn2_io_Stationary_matrix_5_0),
    .io_Stationary_matrix_5_1(my_ivn2_io_Stationary_matrix_5_1),
    .io_Stationary_matrix_5_2(my_ivn2_io_Stationary_matrix_5_2),
    .io_Stationary_matrix_5_3(my_ivn2_io_Stationary_matrix_5_3),
    .io_Stationary_matrix_5_4(my_ivn2_io_Stationary_matrix_5_4),
    .io_Stationary_matrix_5_5(my_ivn2_io_Stationary_matrix_5_5),
    .io_Stationary_matrix_5_6(my_ivn2_io_Stationary_matrix_5_6),
    .io_Stationary_matrix_5_7(my_ivn2_io_Stationary_matrix_5_7),
    .io_Stationary_matrix_6_0(my_ivn2_io_Stationary_matrix_6_0),
    .io_Stationary_matrix_6_1(my_ivn2_io_Stationary_matrix_6_1),
    .io_Stationary_matrix_6_2(my_ivn2_io_Stationary_matrix_6_2),
    .io_Stationary_matrix_6_3(my_ivn2_io_Stationary_matrix_6_3),
    .io_Stationary_matrix_6_4(my_ivn2_io_Stationary_matrix_6_4),
    .io_Stationary_matrix_6_5(my_ivn2_io_Stationary_matrix_6_5),
    .io_Stationary_matrix_6_6(my_ivn2_io_Stationary_matrix_6_6),
    .io_Stationary_matrix_6_7(my_ivn2_io_Stationary_matrix_6_7),
    .io_Stationary_matrix_7_0(my_ivn2_io_Stationary_matrix_7_0),
    .io_Stationary_matrix_7_1(my_ivn2_io_Stationary_matrix_7_1),
    .io_Stationary_matrix_7_2(my_ivn2_io_Stationary_matrix_7_2),
    .io_Stationary_matrix_7_3(my_ivn2_io_Stationary_matrix_7_3),
    .io_Stationary_matrix_7_4(my_ivn2_io_Stationary_matrix_7_4),
    .io_Stationary_matrix_7_5(my_ivn2_io_Stationary_matrix_7_5),
    .io_Stationary_matrix_7_6(my_ivn2_io_Stationary_matrix_7_6),
    .io_Stationary_matrix_7_7(my_ivn2_io_Stationary_matrix_7_7),
    .io_o_vn_0(my_ivn2_io_o_vn_0),
    .io_o_vn_1(my_ivn2_io_o_vn_1),
    .io_o_vn_2(my_ivn2_io_o_vn_2),
    .io_o_vn_3(my_ivn2_io_o_vn_3),
    .io_o_vn2_0(my_ivn2_io_o_vn2_0),
    .io_o_vn2_1(my_ivn2_io_o_vn2_1),
    .io_o_vn2_2(my_ivn2_io_o_vn2_2),
    .io_o_vn2_3(my_ivn2_io_o_vn2_3),
    .io_validpin(my_ivn2_io_validpin)
  );
  ivncontrol4_2 my_ivn3 ( // @[ivntop.scala 86:25]
    .clock(my_ivn3_clock),
    .reset(my_ivn3_reset),
    .io_Stationary_matrix_0_0(my_ivn3_io_Stationary_matrix_0_0),
    .io_Stationary_matrix_0_1(my_ivn3_io_Stationary_matrix_0_1),
    .io_Stationary_matrix_0_2(my_ivn3_io_Stationary_matrix_0_2),
    .io_Stationary_matrix_0_3(my_ivn3_io_Stationary_matrix_0_3),
    .io_Stationary_matrix_0_4(my_ivn3_io_Stationary_matrix_0_4),
    .io_Stationary_matrix_0_5(my_ivn3_io_Stationary_matrix_0_5),
    .io_Stationary_matrix_0_6(my_ivn3_io_Stationary_matrix_0_6),
    .io_Stationary_matrix_0_7(my_ivn3_io_Stationary_matrix_0_7),
    .io_Stationary_matrix_1_0(my_ivn3_io_Stationary_matrix_1_0),
    .io_Stationary_matrix_1_1(my_ivn3_io_Stationary_matrix_1_1),
    .io_Stationary_matrix_1_2(my_ivn3_io_Stationary_matrix_1_2),
    .io_Stationary_matrix_1_3(my_ivn3_io_Stationary_matrix_1_3),
    .io_Stationary_matrix_1_4(my_ivn3_io_Stationary_matrix_1_4),
    .io_Stationary_matrix_1_5(my_ivn3_io_Stationary_matrix_1_5),
    .io_Stationary_matrix_1_6(my_ivn3_io_Stationary_matrix_1_6),
    .io_Stationary_matrix_1_7(my_ivn3_io_Stationary_matrix_1_7),
    .io_Stationary_matrix_2_0(my_ivn3_io_Stationary_matrix_2_0),
    .io_Stationary_matrix_2_1(my_ivn3_io_Stationary_matrix_2_1),
    .io_Stationary_matrix_2_2(my_ivn3_io_Stationary_matrix_2_2),
    .io_Stationary_matrix_2_3(my_ivn3_io_Stationary_matrix_2_3),
    .io_Stationary_matrix_2_4(my_ivn3_io_Stationary_matrix_2_4),
    .io_Stationary_matrix_2_5(my_ivn3_io_Stationary_matrix_2_5),
    .io_Stationary_matrix_2_6(my_ivn3_io_Stationary_matrix_2_6),
    .io_Stationary_matrix_2_7(my_ivn3_io_Stationary_matrix_2_7),
    .io_Stationary_matrix_3_0(my_ivn3_io_Stationary_matrix_3_0),
    .io_Stationary_matrix_3_1(my_ivn3_io_Stationary_matrix_3_1),
    .io_Stationary_matrix_3_2(my_ivn3_io_Stationary_matrix_3_2),
    .io_Stationary_matrix_3_3(my_ivn3_io_Stationary_matrix_3_3),
    .io_Stationary_matrix_3_4(my_ivn3_io_Stationary_matrix_3_4),
    .io_Stationary_matrix_3_5(my_ivn3_io_Stationary_matrix_3_5),
    .io_Stationary_matrix_3_6(my_ivn3_io_Stationary_matrix_3_6),
    .io_Stationary_matrix_3_7(my_ivn3_io_Stationary_matrix_3_7),
    .io_Stationary_matrix_4_0(my_ivn3_io_Stationary_matrix_4_0),
    .io_Stationary_matrix_4_1(my_ivn3_io_Stationary_matrix_4_1),
    .io_Stationary_matrix_4_2(my_ivn3_io_Stationary_matrix_4_2),
    .io_Stationary_matrix_4_3(my_ivn3_io_Stationary_matrix_4_3),
    .io_Stationary_matrix_4_4(my_ivn3_io_Stationary_matrix_4_4),
    .io_Stationary_matrix_4_5(my_ivn3_io_Stationary_matrix_4_5),
    .io_Stationary_matrix_4_6(my_ivn3_io_Stationary_matrix_4_6),
    .io_Stationary_matrix_4_7(my_ivn3_io_Stationary_matrix_4_7),
    .io_Stationary_matrix_5_0(my_ivn3_io_Stationary_matrix_5_0),
    .io_Stationary_matrix_5_1(my_ivn3_io_Stationary_matrix_5_1),
    .io_Stationary_matrix_5_2(my_ivn3_io_Stationary_matrix_5_2),
    .io_Stationary_matrix_5_3(my_ivn3_io_Stationary_matrix_5_3),
    .io_Stationary_matrix_5_4(my_ivn3_io_Stationary_matrix_5_4),
    .io_Stationary_matrix_5_5(my_ivn3_io_Stationary_matrix_5_5),
    .io_Stationary_matrix_5_6(my_ivn3_io_Stationary_matrix_5_6),
    .io_Stationary_matrix_5_7(my_ivn3_io_Stationary_matrix_5_7),
    .io_Stationary_matrix_6_0(my_ivn3_io_Stationary_matrix_6_0),
    .io_Stationary_matrix_6_1(my_ivn3_io_Stationary_matrix_6_1),
    .io_Stationary_matrix_6_2(my_ivn3_io_Stationary_matrix_6_2),
    .io_Stationary_matrix_6_3(my_ivn3_io_Stationary_matrix_6_3),
    .io_Stationary_matrix_6_4(my_ivn3_io_Stationary_matrix_6_4),
    .io_Stationary_matrix_6_5(my_ivn3_io_Stationary_matrix_6_5),
    .io_Stationary_matrix_6_6(my_ivn3_io_Stationary_matrix_6_6),
    .io_Stationary_matrix_6_7(my_ivn3_io_Stationary_matrix_6_7),
    .io_Stationary_matrix_7_0(my_ivn3_io_Stationary_matrix_7_0),
    .io_Stationary_matrix_7_1(my_ivn3_io_Stationary_matrix_7_1),
    .io_Stationary_matrix_7_2(my_ivn3_io_Stationary_matrix_7_2),
    .io_Stationary_matrix_7_3(my_ivn3_io_Stationary_matrix_7_3),
    .io_Stationary_matrix_7_4(my_ivn3_io_Stationary_matrix_7_4),
    .io_Stationary_matrix_7_5(my_ivn3_io_Stationary_matrix_7_5),
    .io_Stationary_matrix_7_6(my_ivn3_io_Stationary_matrix_7_6),
    .io_Stationary_matrix_7_7(my_ivn3_io_Stationary_matrix_7_7),
    .io_o_vn_0(my_ivn3_io_o_vn_0),
    .io_o_vn_1(my_ivn3_io_o_vn_1),
    .io_o_vn_2(my_ivn3_io_o_vn_2),
    .io_o_vn_3(my_ivn3_io_o_vn_3),
    .io_o_vn2_0(my_ivn3_io_o_vn2_0),
    .io_o_vn2_1(my_ivn3_io_o_vn2_1),
    .io_o_vn2_2(my_ivn3_io_o_vn2_2),
    .io_o_vn2_3(my_ivn3_io_o_vn2_3),
    .io_validpin(my_ivn3_io_validpin)
  );
  ivncontrol4_3 my_ivn4 ( // @[ivntop.scala 93:25]
    .clock(my_ivn4_clock),
    .reset(my_ivn4_reset),
    .io_Stationary_matrix_0_0(my_ivn4_io_Stationary_matrix_0_0),
    .io_Stationary_matrix_0_1(my_ivn4_io_Stationary_matrix_0_1),
    .io_Stationary_matrix_0_2(my_ivn4_io_Stationary_matrix_0_2),
    .io_Stationary_matrix_0_3(my_ivn4_io_Stationary_matrix_0_3),
    .io_Stationary_matrix_0_4(my_ivn4_io_Stationary_matrix_0_4),
    .io_Stationary_matrix_0_5(my_ivn4_io_Stationary_matrix_0_5),
    .io_Stationary_matrix_0_6(my_ivn4_io_Stationary_matrix_0_6),
    .io_Stationary_matrix_0_7(my_ivn4_io_Stationary_matrix_0_7),
    .io_Stationary_matrix_1_0(my_ivn4_io_Stationary_matrix_1_0),
    .io_Stationary_matrix_1_1(my_ivn4_io_Stationary_matrix_1_1),
    .io_Stationary_matrix_1_2(my_ivn4_io_Stationary_matrix_1_2),
    .io_Stationary_matrix_1_3(my_ivn4_io_Stationary_matrix_1_3),
    .io_Stationary_matrix_1_4(my_ivn4_io_Stationary_matrix_1_4),
    .io_Stationary_matrix_1_5(my_ivn4_io_Stationary_matrix_1_5),
    .io_Stationary_matrix_1_6(my_ivn4_io_Stationary_matrix_1_6),
    .io_Stationary_matrix_1_7(my_ivn4_io_Stationary_matrix_1_7),
    .io_Stationary_matrix_2_0(my_ivn4_io_Stationary_matrix_2_0),
    .io_Stationary_matrix_2_1(my_ivn4_io_Stationary_matrix_2_1),
    .io_Stationary_matrix_2_2(my_ivn4_io_Stationary_matrix_2_2),
    .io_Stationary_matrix_2_3(my_ivn4_io_Stationary_matrix_2_3),
    .io_Stationary_matrix_2_4(my_ivn4_io_Stationary_matrix_2_4),
    .io_Stationary_matrix_2_5(my_ivn4_io_Stationary_matrix_2_5),
    .io_Stationary_matrix_2_6(my_ivn4_io_Stationary_matrix_2_6),
    .io_Stationary_matrix_2_7(my_ivn4_io_Stationary_matrix_2_7),
    .io_Stationary_matrix_3_0(my_ivn4_io_Stationary_matrix_3_0),
    .io_Stationary_matrix_3_1(my_ivn4_io_Stationary_matrix_3_1),
    .io_Stationary_matrix_3_2(my_ivn4_io_Stationary_matrix_3_2),
    .io_Stationary_matrix_3_3(my_ivn4_io_Stationary_matrix_3_3),
    .io_Stationary_matrix_3_4(my_ivn4_io_Stationary_matrix_3_4),
    .io_Stationary_matrix_3_5(my_ivn4_io_Stationary_matrix_3_5),
    .io_Stationary_matrix_3_6(my_ivn4_io_Stationary_matrix_3_6),
    .io_Stationary_matrix_3_7(my_ivn4_io_Stationary_matrix_3_7),
    .io_Stationary_matrix_4_0(my_ivn4_io_Stationary_matrix_4_0),
    .io_Stationary_matrix_4_1(my_ivn4_io_Stationary_matrix_4_1),
    .io_Stationary_matrix_4_2(my_ivn4_io_Stationary_matrix_4_2),
    .io_Stationary_matrix_4_3(my_ivn4_io_Stationary_matrix_4_3),
    .io_Stationary_matrix_4_4(my_ivn4_io_Stationary_matrix_4_4),
    .io_Stationary_matrix_4_5(my_ivn4_io_Stationary_matrix_4_5),
    .io_Stationary_matrix_4_6(my_ivn4_io_Stationary_matrix_4_6),
    .io_Stationary_matrix_4_7(my_ivn4_io_Stationary_matrix_4_7),
    .io_Stationary_matrix_5_0(my_ivn4_io_Stationary_matrix_5_0),
    .io_Stationary_matrix_5_1(my_ivn4_io_Stationary_matrix_5_1),
    .io_Stationary_matrix_5_2(my_ivn4_io_Stationary_matrix_5_2),
    .io_Stationary_matrix_5_3(my_ivn4_io_Stationary_matrix_5_3),
    .io_Stationary_matrix_5_4(my_ivn4_io_Stationary_matrix_5_4),
    .io_Stationary_matrix_5_5(my_ivn4_io_Stationary_matrix_5_5),
    .io_Stationary_matrix_5_6(my_ivn4_io_Stationary_matrix_5_6),
    .io_Stationary_matrix_5_7(my_ivn4_io_Stationary_matrix_5_7),
    .io_Stationary_matrix_6_0(my_ivn4_io_Stationary_matrix_6_0),
    .io_Stationary_matrix_6_1(my_ivn4_io_Stationary_matrix_6_1),
    .io_Stationary_matrix_6_2(my_ivn4_io_Stationary_matrix_6_2),
    .io_Stationary_matrix_6_3(my_ivn4_io_Stationary_matrix_6_3),
    .io_Stationary_matrix_6_4(my_ivn4_io_Stationary_matrix_6_4),
    .io_Stationary_matrix_6_5(my_ivn4_io_Stationary_matrix_6_5),
    .io_Stationary_matrix_6_6(my_ivn4_io_Stationary_matrix_6_6),
    .io_Stationary_matrix_6_7(my_ivn4_io_Stationary_matrix_6_7),
    .io_Stationary_matrix_7_0(my_ivn4_io_Stationary_matrix_7_0),
    .io_Stationary_matrix_7_1(my_ivn4_io_Stationary_matrix_7_1),
    .io_Stationary_matrix_7_2(my_ivn4_io_Stationary_matrix_7_2),
    .io_Stationary_matrix_7_3(my_ivn4_io_Stationary_matrix_7_3),
    .io_Stationary_matrix_7_4(my_ivn4_io_Stationary_matrix_7_4),
    .io_Stationary_matrix_7_5(my_ivn4_io_Stationary_matrix_7_5),
    .io_Stationary_matrix_7_6(my_ivn4_io_Stationary_matrix_7_6),
    .io_Stationary_matrix_7_7(my_ivn4_io_Stationary_matrix_7_7),
    .io_o_vn_0(my_ivn4_io_o_vn_0),
    .io_o_vn_1(my_ivn4_io_o_vn_1),
    .io_o_vn_2(my_ivn4_io_o_vn_2),
    .io_o_vn_3(my_ivn4_io_o_vn_3),
    .io_o_vn2_0(my_ivn4_io_o_vn2_0),
    .io_o_vn2_1(my_ivn4_io_o_vn2_1),
    .io_o_vn2_2(my_ivn4_io_o_vn2_2),
    .io_o_vn2_3(my_ivn4_io_o_vn2_3),
    .io_validpin(my_ivn4_io_validpin)
  );
  ivncontrol4_4 my_ivn5 ( // @[ivntop.scala 100:25]
    .clock(my_ivn5_clock),
    .reset(my_ivn5_reset),
    .io_Stationary_matrix_0_0(my_ivn5_io_Stationary_matrix_0_0),
    .io_Stationary_matrix_0_1(my_ivn5_io_Stationary_matrix_0_1),
    .io_Stationary_matrix_0_2(my_ivn5_io_Stationary_matrix_0_2),
    .io_Stationary_matrix_0_3(my_ivn5_io_Stationary_matrix_0_3),
    .io_Stationary_matrix_0_4(my_ivn5_io_Stationary_matrix_0_4),
    .io_Stationary_matrix_0_5(my_ivn5_io_Stationary_matrix_0_5),
    .io_Stationary_matrix_0_6(my_ivn5_io_Stationary_matrix_0_6),
    .io_Stationary_matrix_0_7(my_ivn5_io_Stationary_matrix_0_7),
    .io_Stationary_matrix_1_0(my_ivn5_io_Stationary_matrix_1_0),
    .io_Stationary_matrix_1_1(my_ivn5_io_Stationary_matrix_1_1),
    .io_Stationary_matrix_1_2(my_ivn5_io_Stationary_matrix_1_2),
    .io_Stationary_matrix_1_3(my_ivn5_io_Stationary_matrix_1_3),
    .io_Stationary_matrix_1_4(my_ivn5_io_Stationary_matrix_1_4),
    .io_Stationary_matrix_1_5(my_ivn5_io_Stationary_matrix_1_5),
    .io_Stationary_matrix_1_6(my_ivn5_io_Stationary_matrix_1_6),
    .io_Stationary_matrix_1_7(my_ivn5_io_Stationary_matrix_1_7),
    .io_Stationary_matrix_2_0(my_ivn5_io_Stationary_matrix_2_0),
    .io_Stationary_matrix_2_1(my_ivn5_io_Stationary_matrix_2_1),
    .io_Stationary_matrix_2_2(my_ivn5_io_Stationary_matrix_2_2),
    .io_Stationary_matrix_2_3(my_ivn5_io_Stationary_matrix_2_3),
    .io_Stationary_matrix_2_4(my_ivn5_io_Stationary_matrix_2_4),
    .io_Stationary_matrix_2_5(my_ivn5_io_Stationary_matrix_2_5),
    .io_Stationary_matrix_2_6(my_ivn5_io_Stationary_matrix_2_6),
    .io_Stationary_matrix_2_7(my_ivn5_io_Stationary_matrix_2_7),
    .io_Stationary_matrix_3_0(my_ivn5_io_Stationary_matrix_3_0),
    .io_Stationary_matrix_3_1(my_ivn5_io_Stationary_matrix_3_1),
    .io_Stationary_matrix_3_2(my_ivn5_io_Stationary_matrix_3_2),
    .io_Stationary_matrix_3_3(my_ivn5_io_Stationary_matrix_3_3),
    .io_Stationary_matrix_3_4(my_ivn5_io_Stationary_matrix_3_4),
    .io_Stationary_matrix_3_5(my_ivn5_io_Stationary_matrix_3_5),
    .io_Stationary_matrix_3_6(my_ivn5_io_Stationary_matrix_3_6),
    .io_Stationary_matrix_3_7(my_ivn5_io_Stationary_matrix_3_7),
    .io_Stationary_matrix_4_0(my_ivn5_io_Stationary_matrix_4_0),
    .io_Stationary_matrix_4_1(my_ivn5_io_Stationary_matrix_4_1),
    .io_Stationary_matrix_4_2(my_ivn5_io_Stationary_matrix_4_2),
    .io_Stationary_matrix_4_3(my_ivn5_io_Stationary_matrix_4_3),
    .io_Stationary_matrix_4_4(my_ivn5_io_Stationary_matrix_4_4),
    .io_Stationary_matrix_4_5(my_ivn5_io_Stationary_matrix_4_5),
    .io_Stationary_matrix_4_6(my_ivn5_io_Stationary_matrix_4_6),
    .io_Stationary_matrix_4_7(my_ivn5_io_Stationary_matrix_4_7),
    .io_Stationary_matrix_5_0(my_ivn5_io_Stationary_matrix_5_0),
    .io_Stationary_matrix_5_1(my_ivn5_io_Stationary_matrix_5_1),
    .io_Stationary_matrix_5_2(my_ivn5_io_Stationary_matrix_5_2),
    .io_Stationary_matrix_5_3(my_ivn5_io_Stationary_matrix_5_3),
    .io_Stationary_matrix_5_4(my_ivn5_io_Stationary_matrix_5_4),
    .io_Stationary_matrix_5_5(my_ivn5_io_Stationary_matrix_5_5),
    .io_Stationary_matrix_5_6(my_ivn5_io_Stationary_matrix_5_6),
    .io_Stationary_matrix_5_7(my_ivn5_io_Stationary_matrix_5_7),
    .io_Stationary_matrix_6_0(my_ivn5_io_Stationary_matrix_6_0),
    .io_Stationary_matrix_6_1(my_ivn5_io_Stationary_matrix_6_1),
    .io_Stationary_matrix_6_2(my_ivn5_io_Stationary_matrix_6_2),
    .io_Stationary_matrix_6_3(my_ivn5_io_Stationary_matrix_6_3),
    .io_Stationary_matrix_6_4(my_ivn5_io_Stationary_matrix_6_4),
    .io_Stationary_matrix_6_5(my_ivn5_io_Stationary_matrix_6_5),
    .io_Stationary_matrix_6_6(my_ivn5_io_Stationary_matrix_6_6),
    .io_Stationary_matrix_6_7(my_ivn5_io_Stationary_matrix_6_7),
    .io_Stationary_matrix_7_0(my_ivn5_io_Stationary_matrix_7_0),
    .io_Stationary_matrix_7_1(my_ivn5_io_Stationary_matrix_7_1),
    .io_Stationary_matrix_7_2(my_ivn5_io_Stationary_matrix_7_2),
    .io_Stationary_matrix_7_3(my_ivn5_io_Stationary_matrix_7_3),
    .io_Stationary_matrix_7_4(my_ivn5_io_Stationary_matrix_7_4),
    .io_Stationary_matrix_7_5(my_ivn5_io_Stationary_matrix_7_5),
    .io_Stationary_matrix_7_6(my_ivn5_io_Stationary_matrix_7_6),
    .io_Stationary_matrix_7_7(my_ivn5_io_Stationary_matrix_7_7),
    .io_o_vn_0(my_ivn5_io_o_vn_0),
    .io_o_vn_1(my_ivn5_io_o_vn_1),
    .io_o_vn_2(my_ivn5_io_o_vn_2),
    .io_o_vn_3(my_ivn5_io_o_vn_3),
    .io_o_vn2_0(my_ivn5_io_o_vn2_0),
    .io_o_vn2_1(my_ivn5_io_o_vn2_1),
    .io_o_vn2_2(my_ivn5_io_o_vn2_2),
    .io_o_vn2_3(my_ivn5_io_o_vn2_3),
    .io_validpin(my_ivn5_io_validpin)
  );
  ivncontrol4_5 my_ivn6 ( // @[ivntop.scala 107:25]
    .clock(my_ivn6_clock),
    .reset(my_ivn6_reset),
    .io_Stationary_matrix_0_0(my_ivn6_io_Stationary_matrix_0_0),
    .io_Stationary_matrix_0_1(my_ivn6_io_Stationary_matrix_0_1),
    .io_Stationary_matrix_0_2(my_ivn6_io_Stationary_matrix_0_2),
    .io_Stationary_matrix_0_3(my_ivn6_io_Stationary_matrix_0_3),
    .io_Stationary_matrix_0_4(my_ivn6_io_Stationary_matrix_0_4),
    .io_Stationary_matrix_0_5(my_ivn6_io_Stationary_matrix_0_5),
    .io_Stationary_matrix_0_6(my_ivn6_io_Stationary_matrix_0_6),
    .io_Stationary_matrix_0_7(my_ivn6_io_Stationary_matrix_0_7),
    .io_Stationary_matrix_1_0(my_ivn6_io_Stationary_matrix_1_0),
    .io_Stationary_matrix_1_1(my_ivn6_io_Stationary_matrix_1_1),
    .io_Stationary_matrix_1_2(my_ivn6_io_Stationary_matrix_1_2),
    .io_Stationary_matrix_1_3(my_ivn6_io_Stationary_matrix_1_3),
    .io_Stationary_matrix_1_4(my_ivn6_io_Stationary_matrix_1_4),
    .io_Stationary_matrix_1_5(my_ivn6_io_Stationary_matrix_1_5),
    .io_Stationary_matrix_1_6(my_ivn6_io_Stationary_matrix_1_6),
    .io_Stationary_matrix_1_7(my_ivn6_io_Stationary_matrix_1_7),
    .io_Stationary_matrix_2_0(my_ivn6_io_Stationary_matrix_2_0),
    .io_Stationary_matrix_2_1(my_ivn6_io_Stationary_matrix_2_1),
    .io_Stationary_matrix_2_2(my_ivn6_io_Stationary_matrix_2_2),
    .io_Stationary_matrix_2_3(my_ivn6_io_Stationary_matrix_2_3),
    .io_Stationary_matrix_2_4(my_ivn6_io_Stationary_matrix_2_4),
    .io_Stationary_matrix_2_5(my_ivn6_io_Stationary_matrix_2_5),
    .io_Stationary_matrix_2_6(my_ivn6_io_Stationary_matrix_2_6),
    .io_Stationary_matrix_2_7(my_ivn6_io_Stationary_matrix_2_7),
    .io_Stationary_matrix_3_0(my_ivn6_io_Stationary_matrix_3_0),
    .io_Stationary_matrix_3_1(my_ivn6_io_Stationary_matrix_3_1),
    .io_Stationary_matrix_3_2(my_ivn6_io_Stationary_matrix_3_2),
    .io_Stationary_matrix_3_3(my_ivn6_io_Stationary_matrix_3_3),
    .io_Stationary_matrix_3_4(my_ivn6_io_Stationary_matrix_3_4),
    .io_Stationary_matrix_3_5(my_ivn6_io_Stationary_matrix_3_5),
    .io_Stationary_matrix_3_6(my_ivn6_io_Stationary_matrix_3_6),
    .io_Stationary_matrix_3_7(my_ivn6_io_Stationary_matrix_3_7),
    .io_Stationary_matrix_4_0(my_ivn6_io_Stationary_matrix_4_0),
    .io_Stationary_matrix_4_1(my_ivn6_io_Stationary_matrix_4_1),
    .io_Stationary_matrix_4_2(my_ivn6_io_Stationary_matrix_4_2),
    .io_Stationary_matrix_4_3(my_ivn6_io_Stationary_matrix_4_3),
    .io_Stationary_matrix_4_4(my_ivn6_io_Stationary_matrix_4_4),
    .io_Stationary_matrix_4_5(my_ivn6_io_Stationary_matrix_4_5),
    .io_Stationary_matrix_4_6(my_ivn6_io_Stationary_matrix_4_6),
    .io_Stationary_matrix_4_7(my_ivn6_io_Stationary_matrix_4_7),
    .io_Stationary_matrix_5_0(my_ivn6_io_Stationary_matrix_5_0),
    .io_Stationary_matrix_5_1(my_ivn6_io_Stationary_matrix_5_1),
    .io_Stationary_matrix_5_2(my_ivn6_io_Stationary_matrix_5_2),
    .io_Stationary_matrix_5_3(my_ivn6_io_Stationary_matrix_5_3),
    .io_Stationary_matrix_5_4(my_ivn6_io_Stationary_matrix_5_4),
    .io_Stationary_matrix_5_5(my_ivn6_io_Stationary_matrix_5_5),
    .io_Stationary_matrix_5_6(my_ivn6_io_Stationary_matrix_5_6),
    .io_Stationary_matrix_5_7(my_ivn6_io_Stationary_matrix_5_7),
    .io_Stationary_matrix_6_0(my_ivn6_io_Stationary_matrix_6_0),
    .io_Stationary_matrix_6_1(my_ivn6_io_Stationary_matrix_6_1),
    .io_Stationary_matrix_6_2(my_ivn6_io_Stationary_matrix_6_2),
    .io_Stationary_matrix_6_3(my_ivn6_io_Stationary_matrix_6_3),
    .io_Stationary_matrix_6_4(my_ivn6_io_Stationary_matrix_6_4),
    .io_Stationary_matrix_6_5(my_ivn6_io_Stationary_matrix_6_5),
    .io_Stationary_matrix_6_6(my_ivn6_io_Stationary_matrix_6_6),
    .io_Stationary_matrix_6_7(my_ivn6_io_Stationary_matrix_6_7),
    .io_Stationary_matrix_7_0(my_ivn6_io_Stationary_matrix_7_0),
    .io_Stationary_matrix_7_1(my_ivn6_io_Stationary_matrix_7_1),
    .io_Stationary_matrix_7_2(my_ivn6_io_Stationary_matrix_7_2),
    .io_Stationary_matrix_7_3(my_ivn6_io_Stationary_matrix_7_3),
    .io_Stationary_matrix_7_4(my_ivn6_io_Stationary_matrix_7_4),
    .io_Stationary_matrix_7_5(my_ivn6_io_Stationary_matrix_7_5),
    .io_Stationary_matrix_7_6(my_ivn6_io_Stationary_matrix_7_6),
    .io_Stationary_matrix_7_7(my_ivn6_io_Stationary_matrix_7_7),
    .io_o_vn_0(my_ivn6_io_o_vn_0),
    .io_o_vn_1(my_ivn6_io_o_vn_1),
    .io_o_vn_2(my_ivn6_io_o_vn_2),
    .io_o_vn_3(my_ivn6_io_o_vn_3),
    .io_o_vn2_0(my_ivn6_io_o_vn2_0),
    .io_o_vn2_1(my_ivn6_io_o_vn2_1),
    .io_o_vn2_2(my_ivn6_io_o_vn2_2),
    .io_o_vn2_3(my_ivn6_io_o_vn2_3),
    .io_validpin(my_ivn6_io_validpin)
  );
  ivncontrol4_6 my_ivn7 ( // @[ivntop.scala 114:25]
    .clock(my_ivn7_clock),
    .reset(my_ivn7_reset),
    .io_Stationary_matrix_0_0(my_ivn7_io_Stationary_matrix_0_0),
    .io_Stationary_matrix_0_1(my_ivn7_io_Stationary_matrix_0_1),
    .io_Stationary_matrix_0_2(my_ivn7_io_Stationary_matrix_0_2),
    .io_Stationary_matrix_0_3(my_ivn7_io_Stationary_matrix_0_3),
    .io_Stationary_matrix_0_4(my_ivn7_io_Stationary_matrix_0_4),
    .io_Stationary_matrix_0_5(my_ivn7_io_Stationary_matrix_0_5),
    .io_Stationary_matrix_0_6(my_ivn7_io_Stationary_matrix_0_6),
    .io_Stationary_matrix_0_7(my_ivn7_io_Stationary_matrix_0_7),
    .io_Stationary_matrix_1_0(my_ivn7_io_Stationary_matrix_1_0),
    .io_Stationary_matrix_1_1(my_ivn7_io_Stationary_matrix_1_1),
    .io_Stationary_matrix_1_2(my_ivn7_io_Stationary_matrix_1_2),
    .io_Stationary_matrix_1_3(my_ivn7_io_Stationary_matrix_1_3),
    .io_Stationary_matrix_1_4(my_ivn7_io_Stationary_matrix_1_4),
    .io_Stationary_matrix_1_5(my_ivn7_io_Stationary_matrix_1_5),
    .io_Stationary_matrix_1_6(my_ivn7_io_Stationary_matrix_1_6),
    .io_Stationary_matrix_1_7(my_ivn7_io_Stationary_matrix_1_7),
    .io_Stationary_matrix_2_0(my_ivn7_io_Stationary_matrix_2_0),
    .io_Stationary_matrix_2_1(my_ivn7_io_Stationary_matrix_2_1),
    .io_Stationary_matrix_2_2(my_ivn7_io_Stationary_matrix_2_2),
    .io_Stationary_matrix_2_3(my_ivn7_io_Stationary_matrix_2_3),
    .io_Stationary_matrix_2_4(my_ivn7_io_Stationary_matrix_2_4),
    .io_Stationary_matrix_2_5(my_ivn7_io_Stationary_matrix_2_5),
    .io_Stationary_matrix_2_6(my_ivn7_io_Stationary_matrix_2_6),
    .io_Stationary_matrix_2_7(my_ivn7_io_Stationary_matrix_2_7),
    .io_Stationary_matrix_3_0(my_ivn7_io_Stationary_matrix_3_0),
    .io_Stationary_matrix_3_1(my_ivn7_io_Stationary_matrix_3_1),
    .io_Stationary_matrix_3_2(my_ivn7_io_Stationary_matrix_3_2),
    .io_Stationary_matrix_3_3(my_ivn7_io_Stationary_matrix_3_3),
    .io_Stationary_matrix_3_4(my_ivn7_io_Stationary_matrix_3_4),
    .io_Stationary_matrix_3_5(my_ivn7_io_Stationary_matrix_3_5),
    .io_Stationary_matrix_3_6(my_ivn7_io_Stationary_matrix_3_6),
    .io_Stationary_matrix_3_7(my_ivn7_io_Stationary_matrix_3_7),
    .io_Stationary_matrix_4_0(my_ivn7_io_Stationary_matrix_4_0),
    .io_Stationary_matrix_4_1(my_ivn7_io_Stationary_matrix_4_1),
    .io_Stationary_matrix_4_2(my_ivn7_io_Stationary_matrix_4_2),
    .io_Stationary_matrix_4_3(my_ivn7_io_Stationary_matrix_4_3),
    .io_Stationary_matrix_4_4(my_ivn7_io_Stationary_matrix_4_4),
    .io_Stationary_matrix_4_5(my_ivn7_io_Stationary_matrix_4_5),
    .io_Stationary_matrix_4_6(my_ivn7_io_Stationary_matrix_4_6),
    .io_Stationary_matrix_4_7(my_ivn7_io_Stationary_matrix_4_7),
    .io_Stationary_matrix_5_0(my_ivn7_io_Stationary_matrix_5_0),
    .io_Stationary_matrix_5_1(my_ivn7_io_Stationary_matrix_5_1),
    .io_Stationary_matrix_5_2(my_ivn7_io_Stationary_matrix_5_2),
    .io_Stationary_matrix_5_3(my_ivn7_io_Stationary_matrix_5_3),
    .io_Stationary_matrix_5_4(my_ivn7_io_Stationary_matrix_5_4),
    .io_Stationary_matrix_5_5(my_ivn7_io_Stationary_matrix_5_5),
    .io_Stationary_matrix_5_6(my_ivn7_io_Stationary_matrix_5_6),
    .io_Stationary_matrix_5_7(my_ivn7_io_Stationary_matrix_5_7),
    .io_Stationary_matrix_6_0(my_ivn7_io_Stationary_matrix_6_0),
    .io_Stationary_matrix_6_1(my_ivn7_io_Stationary_matrix_6_1),
    .io_Stationary_matrix_6_2(my_ivn7_io_Stationary_matrix_6_2),
    .io_Stationary_matrix_6_3(my_ivn7_io_Stationary_matrix_6_3),
    .io_Stationary_matrix_6_4(my_ivn7_io_Stationary_matrix_6_4),
    .io_Stationary_matrix_6_5(my_ivn7_io_Stationary_matrix_6_5),
    .io_Stationary_matrix_6_6(my_ivn7_io_Stationary_matrix_6_6),
    .io_Stationary_matrix_6_7(my_ivn7_io_Stationary_matrix_6_7),
    .io_Stationary_matrix_7_0(my_ivn7_io_Stationary_matrix_7_0),
    .io_Stationary_matrix_7_1(my_ivn7_io_Stationary_matrix_7_1),
    .io_Stationary_matrix_7_2(my_ivn7_io_Stationary_matrix_7_2),
    .io_Stationary_matrix_7_3(my_ivn7_io_Stationary_matrix_7_3),
    .io_Stationary_matrix_7_4(my_ivn7_io_Stationary_matrix_7_4),
    .io_Stationary_matrix_7_5(my_ivn7_io_Stationary_matrix_7_5),
    .io_Stationary_matrix_7_6(my_ivn7_io_Stationary_matrix_7_6),
    .io_Stationary_matrix_7_7(my_ivn7_io_Stationary_matrix_7_7),
    .io_o_vn_0(my_ivn7_io_o_vn_0),
    .io_o_vn_1(my_ivn7_io_o_vn_1),
    .io_o_vn_2(my_ivn7_io_o_vn_2),
    .io_o_vn_3(my_ivn7_io_o_vn_3),
    .io_o_vn2_0(my_ivn7_io_o_vn2_0),
    .io_o_vn2_1(my_ivn7_io_o_vn2_1),
    .io_o_vn2_2(my_ivn7_io_o_vn2_2),
    .io_o_vn2_3(my_ivn7_io_o_vn2_3),
    .io_validpin(my_ivn7_io_validpin)
  );
  ivncontrol4_7 my_ivn8 ( // @[ivntop.scala 121:25]
    .clock(my_ivn8_clock),
    .reset(my_ivn8_reset),
    .io_Stationary_matrix_0_0(my_ivn8_io_Stationary_matrix_0_0),
    .io_Stationary_matrix_0_1(my_ivn8_io_Stationary_matrix_0_1),
    .io_Stationary_matrix_0_2(my_ivn8_io_Stationary_matrix_0_2),
    .io_Stationary_matrix_0_3(my_ivn8_io_Stationary_matrix_0_3),
    .io_Stationary_matrix_0_4(my_ivn8_io_Stationary_matrix_0_4),
    .io_Stationary_matrix_0_5(my_ivn8_io_Stationary_matrix_0_5),
    .io_Stationary_matrix_0_6(my_ivn8_io_Stationary_matrix_0_6),
    .io_Stationary_matrix_0_7(my_ivn8_io_Stationary_matrix_0_7),
    .io_Stationary_matrix_1_0(my_ivn8_io_Stationary_matrix_1_0),
    .io_Stationary_matrix_1_1(my_ivn8_io_Stationary_matrix_1_1),
    .io_Stationary_matrix_1_2(my_ivn8_io_Stationary_matrix_1_2),
    .io_Stationary_matrix_1_3(my_ivn8_io_Stationary_matrix_1_3),
    .io_Stationary_matrix_1_4(my_ivn8_io_Stationary_matrix_1_4),
    .io_Stationary_matrix_1_5(my_ivn8_io_Stationary_matrix_1_5),
    .io_Stationary_matrix_1_6(my_ivn8_io_Stationary_matrix_1_6),
    .io_Stationary_matrix_1_7(my_ivn8_io_Stationary_matrix_1_7),
    .io_Stationary_matrix_2_0(my_ivn8_io_Stationary_matrix_2_0),
    .io_Stationary_matrix_2_1(my_ivn8_io_Stationary_matrix_2_1),
    .io_Stationary_matrix_2_2(my_ivn8_io_Stationary_matrix_2_2),
    .io_Stationary_matrix_2_3(my_ivn8_io_Stationary_matrix_2_3),
    .io_Stationary_matrix_2_4(my_ivn8_io_Stationary_matrix_2_4),
    .io_Stationary_matrix_2_5(my_ivn8_io_Stationary_matrix_2_5),
    .io_Stationary_matrix_2_6(my_ivn8_io_Stationary_matrix_2_6),
    .io_Stationary_matrix_2_7(my_ivn8_io_Stationary_matrix_2_7),
    .io_Stationary_matrix_3_0(my_ivn8_io_Stationary_matrix_3_0),
    .io_Stationary_matrix_3_1(my_ivn8_io_Stationary_matrix_3_1),
    .io_Stationary_matrix_3_2(my_ivn8_io_Stationary_matrix_3_2),
    .io_Stationary_matrix_3_3(my_ivn8_io_Stationary_matrix_3_3),
    .io_Stationary_matrix_3_4(my_ivn8_io_Stationary_matrix_3_4),
    .io_Stationary_matrix_3_5(my_ivn8_io_Stationary_matrix_3_5),
    .io_Stationary_matrix_3_6(my_ivn8_io_Stationary_matrix_3_6),
    .io_Stationary_matrix_3_7(my_ivn8_io_Stationary_matrix_3_7),
    .io_Stationary_matrix_4_0(my_ivn8_io_Stationary_matrix_4_0),
    .io_Stationary_matrix_4_1(my_ivn8_io_Stationary_matrix_4_1),
    .io_Stationary_matrix_4_2(my_ivn8_io_Stationary_matrix_4_2),
    .io_Stationary_matrix_4_3(my_ivn8_io_Stationary_matrix_4_3),
    .io_Stationary_matrix_4_4(my_ivn8_io_Stationary_matrix_4_4),
    .io_Stationary_matrix_4_5(my_ivn8_io_Stationary_matrix_4_5),
    .io_Stationary_matrix_4_6(my_ivn8_io_Stationary_matrix_4_6),
    .io_Stationary_matrix_4_7(my_ivn8_io_Stationary_matrix_4_7),
    .io_Stationary_matrix_5_0(my_ivn8_io_Stationary_matrix_5_0),
    .io_Stationary_matrix_5_1(my_ivn8_io_Stationary_matrix_5_1),
    .io_Stationary_matrix_5_2(my_ivn8_io_Stationary_matrix_5_2),
    .io_Stationary_matrix_5_3(my_ivn8_io_Stationary_matrix_5_3),
    .io_Stationary_matrix_5_4(my_ivn8_io_Stationary_matrix_5_4),
    .io_Stationary_matrix_5_5(my_ivn8_io_Stationary_matrix_5_5),
    .io_Stationary_matrix_5_6(my_ivn8_io_Stationary_matrix_5_6),
    .io_Stationary_matrix_5_7(my_ivn8_io_Stationary_matrix_5_7),
    .io_Stationary_matrix_6_0(my_ivn8_io_Stationary_matrix_6_0),
    .io_Stationary_matrix_6_1(my_ivn8_io_Stationary_matrix_6_1),
    .io_Stationary_matrix_6_2(my_ivn8_io_Stationary_matrix_6_2),
    .io_Stationary_matrix_6_3(my_ivn8_io_Stationary_matrix_6_3),
    .io_Stationary_matrix_6_4(my_ivn8_io_Stationary_matrix_6_4),
    .io_Stationary_matrix_6_5(my_ivn8_io_Stationary_matrix_6_5),
    .io_Stationary_matrix_6_6(my_ivn8_io_Stationary_matrix_6_6),
    .io_Stationary_matrix_6_7(my_ivn8_io_Stationary_matrix_6_7),
    .io_Stationary_matrix_7_0(my_ivn8_io_Stationary_matrix_7_0),
    .io_Stationary_matrix_7_1(my_ivn8_io_Stationary_matrix_7_1),
    .io_Stationary_matrix_7_2(my_ivn8_io_Stationary_matrix_7_2),
    .io_Stationary_matrix_7_3(my_ivn8_io_Stationary_matrix_7_3),
    .io_Stationary_matrix_7_4(my_ivn8_io_Stationary_matrix_7_4),
    .io_Stationary_matrix_7_5(my_ivn8_io_Stationary_matrix_7_5),
    .io_Stationary_matrix_7_6(my_ivn8_io_Stationary_matrix_7_6),
    .io_Stationary_matrix_7_7(my_ivn8_io_Stationary_matrix_7_7),
    .io_o_vn_0(my_ivn8_io_o_vn_0),
    .io_o_vn_1(my_ivn8_io_o_vn_1),
    .io_o_vn_2(my_ivn8_io_o_vn_2),
    .io_o_vn_3(my_ivn8_io_o_vn_3),
    .io_o_vn2_0(my_ivn8_io_o_vn2_0),
    .io_o_vn2_1(my_ivn8_io_o_vn2_1),
    .io_o_vn2_2(my_ivn8_io_o_vn2_2),
    .io_o_vn2_3(my_ivn8_io_o_vn2_3),
    .io_validpin(my_ivn8_io_validpin)
  );
  assign io_ProcessValid = my_ivn1_io_ProcessValid; // @[ivntop.scala 74:21]
  assign io_o_vn_0_0 = i_vn_0_0; // @[ivntop.scala 16:12]
  assign io_o_vn_0_1 = i_vn_0_1; // @[ivntop.scala 16:12]
  assign io_o_vn_0_2 = i_vn_0_2; // @[ivntop.scala 16:12]
  assign io_o_vn_0_3 = i_vn_0_3; // @[ivntop.scala 16:12]
  assign io_o_vn_1_0 = i_vn_1_0; // @[ivntop.scala 16:12]
  assign io_o_vn_1_1 = i_vn_1_1; // @[ivntop.scala 16:12]
  assign io_o_vn_1_2 = i_vn_1_2; // @[ivntop.scala 16:12]
  assign io_o_vn_1_3 = i_vn_1_3; // @[ivntop.scala 16:12]
  assign io_o_vn_2_0 = i_vn_2_0; // @[ivntop.scala 16:12]
  assign io_o_vn_2_1 = i_vn_2_1; // @[ivntop.scala 16:12]
  assign io_o_vn_2_2 = i_vn_2_2; // @[ivntop.scala 16:12]
  assign io_o_vn_2_3 = i_vn_2_3; // @[ivntop.scala 16:12]
  assign io_o_vn_3_0 = i_vn_3_0; // @[ivntop.scala 16:12]
  assign io_o_vn_3_1 = i_vn_3_1; // @[ivntop.scala 16:12]
  assign io_o_vn_3_2 = i_vn_3_2; // @[ivntop.scala 16:12]
  assign io_o_vn_3_3 = i_vn_3_3; // @[ivntop.scala 16:12]
  assign io_o_vn_4_0 = i_vn_4_0; // @[ivntop.scala 16:12]
  assign io_o_vn_4_1 = i_vn_4_1; // @[ivntop.scala 16:12]
  assign io_o_vn_4_2 = i_vn_4_2; // @[ivntop.scala 16:12]
  assign io_o_vn_4_3 = i_vn_4_3; // @[ivntop.scala 16:12]
  assign io_o_vn_5_0 = i_vn_5_0; // @[ivntop.scala 16:12]
  assign io_o_vn_5_1 = i_vn_5_1; // @[ivntop.scala 16:12]
  assign io_o_vn_5_2 = i_vn_5_2; // @[ivntop.scala 16:12]
  assign io_o_vn_5_3 = i_vn_5_3; // @[ivntop.scala 16:12]
  assign io_o_vn_6_0 = i_vn_6_0; // @[ivntop.scala 16:12]
  assign io_o_vn_6_1 = i_vn_6_1; // @[ivntop.scala 16:12]
  assign io_o_vn_6_2 = i_vn_6_2; // @[ivntop.scala 16:12]
  assign io_o_vn_6_3 = i_vn_6_3; // @[ivntop.scala 16:12]
  assign io_o_vn_7_0 = i_vn_7_0; // @[ivntop.scala 16:12]
  assign io_o_vn_7_1 = i_vn_7_1; // @[ivntop.scala 16:12]
  assign io_o_vn_7_2 = i_vn_7_2; // @[ivntop.scala 16:12]
  assign io_o_vn_7_3 = i_vn_7_3; // @[ivntop.scala 16:12]
  assign io_o_vn_8_0 = i_vn_8_0; // @[ivntop.scala 16:12]
  assign io_o_vn_8_1 = i_vn_8_1; // @[ivntop.scala 16:12]
  assign io_o_vn_8_2 = i_vn_8_2; // @[ivntop.scala 16:12]
  assign io_o_vn_8_3 = i_vn_8_3; // @[ivntop.scala 16:12]
  assign io_o_vn_9_0 = i_vn_9_0; // @[ivntop.scala 16:12]
  assign io_o_vn_9_1 = i_vn_9_1; // @[ivntop.scala 16:12]
  assign io_o_vn_9_2 = i_vn_9_2; // @[ivntop.scala 16:12]
  assign io_o_vn_9_3 = i_vn_9_3; // @[ivntop.scala 16:12]
  assign io_o_vn_10_0 = i_vn_10_0; // @[ivntop.scala 16:12]
  assign io_o_vn_10_1 = i_vn_10_1; // @[ivntop.scala 16:12]
  assign io_o_vn_10_2 = i_vn_10_2; // @[ivntop.scala 16:12]
  assign io_o_vn_10_3 = i_vn_10_3; // @[ivntop.scala 16:12]
  assign io_o_vn_11_0 = i_vn_11_0; // @[ivntop.scala 16:12]
  assign io_o_vn_11_1 = i_vn_11_1; // @[ivntop.scala 16:12]
  assign io_o_vn_11_2 = i_vn_11_2; // @[ivntop.scala 16:12]
  assign io_o_vn_11_3 = i_vn_11_3; // @[ivntop.scala 16:12]
  assign io_o_vn_12_0 = i_vn_12_0; // @[ivntop.scala 16:12]
  assign io_o_vn_12_1 = i_vn_12_1; // @[ivntop.scala 16:12]
  assign io_o_vn_12_2 = i_vn_12_2; // @[ivntop.scala 16:12]
  assign io_o_vn_12_3 = i_vn_12_3; // @[ivntop.scala 16:12]
  assign io_o_vn_13_0 = i_vn_13_0; // @[ivntop.scala 16:12]
  assign io_o_vn_13_1 = i_vn_13_1; // @[ivntop.scala 16:12]
  assign io_o_vn_13_2 = i_vn_13_2; // @[ivntop.scala 16:12]
  assign io_o_vn_13_3 = i_vn_13_3; // @[ivntop.scala 16:12]
  assign io_o_vn_14_0 = i_vn_14_0; // @[ivntop.scala 16:12]
  assign io_o_vn_14_1 = i_vn_14_1; // @[ivntop.scala 16:12]
  assign io_o_vn_14_2 = i_vn_14_2; // @[ivntop.scala 16:12]
  assign io_o_vn_14_3 = i_vn_14_3; // @[ivntop.scala 16:12]
  assign io_o_vn_15_0 = i_vn_15_0; // @[ivntop.scala 16:12]
  assign io_o_vn_15_1 = i_vn_15_1; // @[ivntop.scala 16:12]
  assign io_o_vn_15_2 = i_vn_15_2; // @[ivntop.scala 16:12]
  assign io_o_vn_15_3 = i_vn_15_3; // @[ivntop.scala 16:12]
  assign my_stationary_clock = clock;
  assign my_stationary_reset = reset;
  assign my_stationary_io_Stationary_matrix_0_0 = io_Stationary_matrix_0_0; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_0_1 = io_Stationary_matrix_0_1; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_0_2 = io_Stationary_matrix_0_2; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_0_3 = io_Stationary_matrix_0_3; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_0_4 = io_Stationary_matrix_0_4; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_0_5 = io_Stationary_matrix_0_5; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_0_6 = io_Stationary_matrix_0_6; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_0_7 = io_Stationary_matrix_0_7; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_1_0 = io_Stationary_matrix_1_0; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_1_1 = io_Stationary_matrix_1_1; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_1_2 = io_Stationary_matrix_1_2; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_1_3 = io_Stationary_matrix_1_3; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_1_4 = io_Stationary_matrix_1_4; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_1_5 = io_Stationary_matrix_1_5; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_1_6 = io_Stationary_matrix_1_6; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_1_7 = io_Stationary_matrix_1_7; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_2_0 = io_Stationary_matrix_2_0; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_2_1 = io_Stationary_matrix_2_1; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_2_2 = io_Stationary_matrix_2_2; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_2_3 = io_Stationary_matrix_2_3; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_2_4 = io_Stationary_matrix_2_4; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_2_5 = io_Stationary_matrix_2_5; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_2_6 = io_Stationary_matrix_2_6; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_2_7 = io_Stationary_matrix_2_7; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_3_0 = io_Stationary_matrix_3_0; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_3_1 = io_Stationary_matrix_3_1; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_3_2 = io_Stationary_matrix_3_2; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_3_3 = io_Stationary_matrix_3_3; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_3_4 = io_Stationary_matrix_3_4; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_3_5 = io_Stationary_matrix_3_5; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_3_6 = io_Stationary_matrix_3_6; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_3_7 = io_Stationary_matrix_3_7; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_4_0 = io_Stationary_matrix_4_0; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_4_1 = io_Stationary_matrix_4_1; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_4_2 = io_Stationary_matrix_4_2; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_4_3 = io_Stationary_matrix_4_3; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_4_4 = io_Stationary_matrix_4_4; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_4_5 = io_Stationary_matrix_4_5; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_4_6 = io_Stationary_matrix_4_6; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_4_7 = io_Stationary_matrix_4_7; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_5_0 = io_Stationary_matrix_5_0; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_5_1 = io_Stationary_matrix_5_1; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_5_2 = io_Stationary_matrix_5_2; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_5_3 = io_Stationary_matrix_5_3; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_5_4 = io_Stationary_matrix_5_4; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_5_5 = io_Stationary_matrix_5_5; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_5_6 = io_Stationary_matrix_5_6; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_5_7 = io_Stationary_matrix_5_7; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_6_0 = io_Stationary_matrix_6_0; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_6_1 = io_Stationary_matrix_6_1; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_6_2 = io_Stationary_matrix_6_2; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_6_3 = io_Stationary_matrix_6_3; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_6_4 = io_Stationary_matrix_6_4; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_6_5 = io_Stationary_matrix_6_5; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_6_6 = io_Stationary_matrix_6_6; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_6_7 = io_Stationary_matrix_6_7; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_7_0 = io_Stationary_matrix_7_0; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_7_1 = io_Stationary_matrix_7_1; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_7_2 = io_Stationary_matrix_7_2; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_7_3 = io_Stationary_matrix_7_3; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_7_4 = io_Stationary_matrix_7_4; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_7_5 = io_Stationary_matrix_7_5; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_7_6 = io_Stationary_matrix_7_6; // @[ivntop.scala 30:40]
  assign my_stationary_io_Stationary_matrix_7_7 = io_Stationary_matrix_7_7; // @[ivntop.scala 30:40]
  assign my_ivn1_clock = clock;
  assign my_ivn1_reset = reset;
  assign my_ivn1_io_Stationary_matrix_0_0 = my_stationary_io_o_Stationary_matrix1_0_0; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_0_1 = my_stationary_io_o_Stationary_matrix1_0_1; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_0_2 = my_stationary_io_o_Stationary_matrix1_0_2; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_0_3 = my_stationary_io_o_Stationary_matrix1_0_3; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_0_4 = my_stationary_io_o_Stationary_matrix1_0_4; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_0_5 = my_stationary_io_o_Stationary_matrix1_0_5; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_0_6 = my_stationary_io_o_Stationary_matrix1_0_6; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_0_7 = my_stationary_io_o_Stationary_matrix1_0_7; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_1_0 = my_stationary_io_o_Stationary_matrix1_1_0; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_1_1 = my_stationary_io_o_Stationary_matrix1_1_1; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_1_2 = my_stationary_io_o_Stationary_matrix1_1_2; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_1_3 = my_stationary_io_o_Stationary_matrix1_1_3; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_1_4 = my_stationary_io_o_Stationary_matrix1_1_4; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_1_5 = my_stationary_io_o_Stationary_matrix1_1_5; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_1_6 = my_stationary_io_o_Stationary_matrix1_1_6; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_1_7 = my_stationary_io_o_Stationary_matrix1_1_7; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_2_0 = my_stationary_io_o_Stationary_matrix1_2_0; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_2_1 = my_stationary_io_o_Stationary_matrix1_2_1; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_2_2 = my_stationary_io_o_Stationary_matrix1_2_2; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_2_3 = my_stationary_io_o_Stationary_matrix1_2_3; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_2_4 = my_stationary_io_o_Stationary_matrix1_2_4; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_2_5 = my_stationary_io_o_Stationary_matrix1_2_5; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_2_6 = my_stationary_io_o_Stationary_matrix1_2_6; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_2_7 = my_stationary_io_o_Stationary_matrix1_2_7; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_3_0 = my_stationary_io_o_Stationary_matrix1_3_0; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_3_1 = my_stationary_io_o_Stationary_matrix1_3_1; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_3_2 = my_stationary_io_o_Stationary_matrix1_3_2; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_3_3 = my_stationary_io_o_Stationary_matrix1_3_3; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_3_4 = my_stationary_io_o_Stationary_matrix1_3_4; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_3_5 = my_stationary_io_o_Stationary_matrix1_3_5; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_3_6 = my_stationary_io_o_Stationary_matrix1_3_6; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_3_7 = my_stationary_io_o_Stationary_matrix1_3_7; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_4_0 = my_stationary_io_o_Stationary_matrix1_4_0; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_4_1 = my_stationary_io_o_Stationary_matrix1_4_1; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_4_2 = my_stationary_io_o_Stationary_matrix1_4_2; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_4_3 = my_stationary_io_o_Stationary_matrix1_4_3; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_4_4 = my_stationary_io_o_Stationary_matrix1_4_4; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_4_5 = my_stationary_io_o_Stationary_matrix1_4_5; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_4_6 = my_stationary_io_o_Stationary_matrix1_4_6; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_4_7 = my_stationary_io_o_Stationary_matrix1_4_7; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_5_0 = my_stationary_io_o_Stationary_matrix1_5_0; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_5_1 = my_stationary_io_o_Stationary_matrix1_5_1; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_5_2 = my_stationary_io_o_Stationary_matrix1_5_2; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_5_3 = my_stationary_io_o_Stationary_matrix1_5_3; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_5_4 = my_stationary_io_o_Stationary_matrix1_5_4; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_5_5 = my_stationary_io_o_Stationary_matrix1_5_5; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_5_6 = my_stationary_io_o_Stationary_matrix1_5_6; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_5_7 = my_stationary_io_o_Stationary_matrix1_5_7; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_6_0 = my_stationary_io_o_Stationary_matrix1_6_0; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_6_1 = my_stationary_io_o_Stationary_matrix1_6_1; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_6_2 = my_stationary_io_o_Stationary_matrix1_6_2; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_6_3 = my_stationary_io_o_Stationary_matrix1_6_3; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_6_4 = my_stationary_io_o_Stationary_matrix1_6_4; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_6_5 = my_stationary_io_o_Stationary_matrix1_6_5; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_6_6 = my_stationary_io_o_Stationary_matrix1_6_6; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_6_7 = my_stationary_io_o_Stationary_matrix1_6_7; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_7_0 = my_stationary_io_o_Stationary_matrix1_7_0; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_7_1 = my_stationary_io_o_Stationary_matrix1_7_1; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_7_2 = my_stationary_io_o_Stationary_matrix1_7_2; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_7_3 = my_stationary_io_o_Stationary_matrix1_7_3; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_7_4 = my_stationary_io_o_Stationary_matrix1_7_4; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_7_5 = my_stationary_io_o_Stationary_matrix1_7_5; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_7_6 = my_stationary_io_o_Stationary_matrix1_7_6; // @[ivntop.scala 70:34]
  assign my_ivn1_io_Stationary_matrix_7_7 = my_stationary_io_o_Stationary_matrix1_7_7; // @[ivntop.scala 70:34]
  assign my_ivn1_io_validpin = _T; // @[ivntop.scala 75:25]
  assign my_ivn2_clock = clock;
  assign my_ivn2_reset = reset;
  assign my_ivn2_io_Stationary_matrix_0_0 = my_stationary_io_o_Stationary_matrix2_0_0; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_0_1 = my_stationary_io_o_Stationary_matrix2_0_1; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_0_2 = my_stationary_io_o_Stationary_matrix2_0_2; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_0_3 = my_stationary_io_o_Stationary_matrix2_0_3; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_0_4 = my_stationary_io_o_Stationary_matrix2_0_4; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_0_5 = my_stationary_io_o_Stationary_matrix2_0_5; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_0_6 = my_stationary_io_o_Stationary_matrix2_0_6; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_0_7 = my_stationary_io_o_Stationary_matrix2_0_7; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_1_0 = my_stationary_io_o_Stationary_matrix2_1_0; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_1_1 = my_stationary_io_o_Stationary_matrix2_1_1; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_1_2 = my_stationary_io_o_Stationary_matrix2_1_2; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_1_3 = my_stationary_io_o_Stationary_matrix2_1_3; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_1_4 = my_stationary_io_o_Stationary_matrix2_1_4; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_1_5 = my_stationary_io_o_Stationary_matrix2_1_5; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_1_6 = my_stationary_io_o_Stationary_matrix2_1_6; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_1_7 = my_stationary_io_o_Stationary_matrix2_1_7; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_2_0 = my_stationary_io_o_Stationary_matrix2_2_0; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_2_1 = my_stationary_io_o_Stationary_matrix2_2_1; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_2_2 = my_stationary_io_o_Stationary_matrix2_2_2; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_2_3 = my_stationary_io_o_Stationary_matrix2_2_3; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_2_4 = my_stationary_io_o_Stationary_matrix2_2_4; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_2_5 = my_stationary_io_o_Stationary_matrix2_2_5; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_2_6 = my_stationary_io_o_Stationary_matrix2_2_6; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_2_7 = my_stationary_io_o_Stationary_matrix2_2_7; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_3_0 = my_stationary_io_o_Stationary_matrix2_3_0; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_3_1 = my_stationary_io_o_Stationary_matrix2_3_1; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_3_2 = my_stationary_io_o_Stationary_matrix2_3_2; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_3_3 = my_stationary_io_o_Stationary_matrix2_3_3; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_3_4 = my_stationary_io_o_Stationary_matrix2_3_4; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_3_5 = my_stationary_io_o_Stationary_matrix2_3_5; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_3_6 = my_stationary_io_o_Stationary_matrix2_3_6; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_3_7 = my_stationary_io_o_Stationary_matrix2_3_7; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_4_0 = my_stationary_io_o_Stationary_matrix2_4_0; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_4_1 = my_stationary_io_o_Stationary_matrix2_4_1; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_4_2 = my_stationary_io_o_Stationary_matrix2_4_2; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_4_3 = my_stationary_io_o_Stationary_matrix2_4_3; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_4_4 = my_stationary_io_o_Stationary_matrix2_4_4; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_4_5 = my_stationary_io_o_Stationary_matrix2_4_5; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_4_6 = my_stationary_io_o_Stationary_matrix2_4_6; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_4_7 = my_stationary_io_o_Stationary_matrix2_4_7; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_5_0 = my_stationary_io_o_Stationary_matrix2_5_0; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_5_1 = my_stationary_io_o_Stationary_matrix2_5_1; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_5_2 = my_stationary_io_o_Stationary_matrix2_5_2; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_5_3 = my_stationary_io_o_Stationary_matrix2_5_3; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_5_4 = my_stationary_io_o_Stationary_matrix2_5_4; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_5_5 = my_stationary_io_o_Stationary_matrix2_5_5; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_5_6 = my_stationary_io_o_Stationary_matrix2_5_6; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_5_7 = my_stationary_io_o_Stationary_matrix2_5_7; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_6_0 = my_stationary_io_o_Stationary_matrix2_6_0; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_6_1 = my_stationary_io_o_Stationary_matrix2_6_1; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_6_2 = my_stationary_io_o_Stationary_matrix2_6_2; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_6_3 = my_stationary_io_o_Stationary_matrix2_6_3; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_6_4 = my_stationary_io_o_Stationary_matrix2_6_4; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_6_5 = my_stationary_io_o_Stationary_matrix2_6_5; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_6_6 = my_stationary_io_o_Stationary_matrix2_6_6; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_6_7 = my_stationary_io_o_Stationary_matrix2_6_7; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_7_0 = my_stationary_io_o_Stationary_matrix2_7_0; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_7_1 = my_stationary_io_o_Stationary_matrix2_7_1; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_7_2 = my_stationary_io_o_Stationary_matrix2_7_2; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_7_3 = my_stationary_io_o_Stationary_matrix2_7_3; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_7_4 = my_stationary_io_o_Stationary_matrix2_7_4; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_7_5 = my_stationary_io_o_Stationary_matrix2_7_5; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_7_6 = my_stationary_io_o_Stationary_matrix2_7_6; // @[ivntop.scala 79:34]
  assign my_ivn2_io_Stationary_matrix_7_7 = my_stationary_io_o_Stationary_matrix2_7_7; // @[ivntop.scala 79:34]
  assign my_ivn2_io_validpin = counter >= 32'h14; // @[ivntop.scala 43:16]
  assign my_ivn3_clock = clock;
  assign my_ivn3_reset = reset;
  assign my_ivn3_io_Stationary_matrix_0_0 = my_stationary_io_o_Stationary_matrix3_0_0; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_0_1 = my_stationary_io_o_Stationary_matrix3_0_1; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_0_2 = my_stationary_io_o_Stationary_matrix3_0_2; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_0_3 = my_stationary_io_o_Stationary_matrix3_0_3; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_0_4 = my_stationary_io_o_Stationary_matrix3_0_4; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_0_5 = my_stationary_io_o_Stationary_matrix3_0_5; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_0_6 = my_stationary_io_o_Stationary_matrix3_0_6; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_0_7 = my_stationary_io_o_Stationary_matrix3_0_7; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_1_0 = my_stationary_io_o_Stationary_matrix3_1_0; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_1_1 = my_stationary_io_o_Stationary_matrix3_1_1; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_1_2 = my_stationary_io_o_Stationary_matrix3_1_2; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_1_3 = my_stationary_io_o_Stationary_matrix3_1_3; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_1_4 = my_stationary_io_o_Stationary_matrix3_1_4; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_1_5 = my_stationary_io_o_Stationary_matrix3_1_5; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_1_6 = my_stationary_io_o_Stationary_matrix3_1_6; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_1_7 = my_stationary_io_o_Stationary_matrix3_1_7; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_2_0 = my_stationary_io_o_Stationary_matrix3_2_0; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_2_1 = my_stationary_io_o_Stationary_matrix3_2_1; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_2_2 = my_stationary_io_o_Stationary_matrix3_2_2; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_2_3 = my_stationary_io_o_Stationary_matrix3_2_3; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_2_4 = my_stationary_io_o_Stationary_matrix3_2_4; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_2_5 = my_stationary_io_o_Stationary_matrix3_2_5; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_2_6 = my_stationary_io_o_Stationary_matrix3_2_6; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_2_7 = my_stationary_io_o_Stationary_matrix3_2_7; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_3_0 = my_stationary_io_o_Stationary_matrix3_3_0; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_3_1 = my_stationary_io_o_Stationary_matrix3_3_1; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_3_2 = my_stationary_io_o_Stationary_matrix3_3_2; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_3_3 = my_stationary_io_o_Stationary_matrix3_3_3; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_3_4 = my_stationary_io_o_Stationary_matrix3_3_4; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_3_5 = my_stationary_io_o_Stationary_matrix3_3_5; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_3_6 = my_stationary_io_o_Stationary_matrix3_3_6; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_3_7 = my_stationary_io_o_Stationary_matrix3_3_7; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_4_0 = my_stationary_io_o_Stationary_matrix3_4_0; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_4_1 = my_stationary_io_o_Stationary_matrix3_4_1; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_4_2 = my_stationary_io_o_Stationary_matrix3_4_2; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_4_3 = my_stationary_io_o_Stationary_matrix3_4_3; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_4_4 = my_stationary_io_o_Stationary_matrix3_4_4; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_4_5 = my_stationary_io_o_Stationary_matrix3_4_5; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_4_6 = my_stationary_io_o_Stationary_matrix3_4_6; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_4_7 = my_stationary_io_o_Stationary_matrix3_4_7; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_5_0 = my_stationary_io_o_Stationary_matrix3_5_0; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_5_1 = my_stationary_io_o_Stationary_matrix3_5_1; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_5_2 = my_stationary_io_o_Stationary_matrix3_5_2; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_5_3 = my_stationary_io_o_Stationary_matrix3_5_3; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_5_4 = my_stationary_io_o_Stationary_matrix3_5_4; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_5_5 = my_stationary_io_o_Stationary_matrix3_5_5; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_5_6 = my_stationary_io_o_Stationary_matrix3_5_6; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_5_7 = my_stationary_io_o_Stationary_matrix3_5_7; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_6_0 = my_stationary_io_o_Stationary_matrix3_6_0; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_6_1 = my_stationary_io_o_Stationary_matrix3_6_1; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_6_2 = my_stationary_io_o_Stationary_matrix3_6_2; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_6_3 = my_stationary_io_o_Stationary_matrix3_6_3; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_6_4 = my_stationary_io_o_Stationary_matrix3_6_4; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_6_5 = my_stationary_io_o_Stationary_matrix3_6_5; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_6_6 = my_stationary_io_o_Stationary_matrix3_6_6; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_6_7 = my_stationary_io_o_Stationary_matrix3_6_7; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_7_0 = my_stationary_io_o_Stationary_matrix3_7_0; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_7_1 = my_stationary_io_o_Stationary_matrix3_7_1; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_7_2 = my_stationary_io_o_Stationary_matrix3_7_2; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_7_3 = my_stationary_io_o_Stationary_matrix3_7_3; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_7_4 = my_stationary_io_o_Stationary_matrix3_7_4; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_7_5 = my_stationary_io_o_Stationary_matrix3_7_5; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_7_6 = my_stationary_io_o_Stationary_matrix3_7_6; // @[ivntop.scala 87:34]
  assign my_ivn3_io_Stationary_matrix_7_7 = my_stationary_io_o_Stationary_matrix3_7_7; // @[ivntop.scala 87:34]
  assign my_ivn3_io_validpin = counter >= 32'h1e; // @[ivntop.scala 46:16]
  assign my_ivn4_clock = clock;
  assign my_ivn4_reset = reset;
  assign my_ivn4_io_Stationary_matrix_0_0 = my_stationary_io_o_Stationary_matrix4_0_0; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_0_1 = my_stationary_io_o_Stationary_matrix4_0_1; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_0_2 = my_stationary_io_o_Stationary_matrix4_0_2; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_0_3 = my_stationary_io_o_Stationary_matrix4_0_3; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_0_4 = my_stationary_io_o_Stationary_matrix4_0_4; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_0_5 = my_stationary_io_o_Stationary_matrix4_0_5; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_0_6 = my_stationary_io_o_Stationary_matrix4_0_6; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_0_7 = my_stationary_io_o_Stationary_matrix4_0_7; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_1_0 = my_stationary_io_o_Stationary_matrix4_1_0; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_1_1 = my_stationary_io_o_Stationary_matrix4_1_1; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_1_2 = my_stationary_io_o_Stationary_matrix4_1_2; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_1_3 = my_stationary_io_o_Stationary_matrix4_1_3; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_1_4 = my_stationary_io_o_Stationary_matrix4_1_4; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_1_5 = my_stationary_io_o_Stationary_matrix4_1_5; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_1_6 = my_stationary_io_o_Stationary_matrix4_1_6; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_1_7 = my_stationary_io_o_Stationary_matrix4_1_7; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_2_0 = my_stationary_io_o_Stationary_matrix4_2_0; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_2_1 = my_stationary_io_o_Stationary_matrix4_2_1; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_2_2 = my_stationary_io_o_Stationary_matrix4_2_2; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_2_3 = my_stationary_io_o_Stationary_matrix4_2_3; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_2_4 = my_stationary_io_o_Stationary_matrix4_2_4; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_2_5 = my_stationary_io_o_Stationary_matrix4_2_5; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_2_6 = my_stationary_io_o_Stationary_matrix4_2_6; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_2_7 = my_stationary_io_o_Stationary_matrix4_2_7; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_3_0 = my_stationary_io_o_Stationary_matrix4_3_0; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_3_1 = my_stationary_io_o_Stationary_matrix4_3_1; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_3_2 = my_stationary_io_o_Stationary_matrix4_3_2; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_3_3 = my_stationary_io_o_Stationary_matrix4_3_3; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_3_4 = my_stationary_io_o_Stationary_matrix4_3_4; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_3_5 = my_stationary_io_o_Stationary_matrix4_3_5; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_3_6 = my_stationary_io_o_Stationary_matrix4_3_6; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_3_7 = my_stationary_io_o_Stationary_matrix4_3_7; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_4_0 = my_stationary_io_o_Stationary_matrix4_4_0; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_4_1 = my_stationary_io_o_Stationary_matrix4_4_1; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_4_2 = my_stationary_io_o_Stationary_matrix4_4_2; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_4_3 = my_stationary_io_o_Stationary_matrix4_4_3; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_4_4 = my_stationary_io_o_Stationary_matrix4_4_4; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_4_5 = my_stationary_io_o_Stationary_matrix4_4_5; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_4_6 = my_stationary_io_o_Stationary_matrix4_4_6; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_4_7 = my_stationary_io_o_Stationary_matrix4_4_7; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_5_0 = my_stationary_io_o_Stationary_matrix4_5_0; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_5_1 = my_stationary_io_o_Stationary_matrix4_5_1; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_5_2 = my_stationary_io_o_Stationary_matrix4_5_2; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_5_3 = my_stationary_io_o_Stationary_matrix4_5_3; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_5_4 = my_stationary_io_o_Stationary_matrix4_5_4; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_5_5 = my_stationary_io_o_Stationary_matrix4_5_5; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_5_6 = my_stationary_io_o_Stationary_matrix4_5_6; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_5_7 = my_stationary_io_o_Stationary_matrix4_5_7; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_6_0 = my_stationary_io_o_Stationary_matrix4_6_0; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_6_1 = my_stationary_io_o_Stationary_matrix4_6_1; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_6_2 = my_stationary_io_o_Stationary_matrix4_6_2; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_6_3 = my_stationary_io_o_Stationary_matrix4_6_3; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_6_4 = my_stationary_io_o_Stationary_matrix4_6_4; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_6_5 = my_stationary_io_o_Stationary_matrix4_6_5; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_6_6 = my_stationary_io_o_Stationary_matrix4_6_6; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_6_7 = my_stationary_io_o_Stationary_matrix4_6_7; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_7_0 = my_stationary_io_o_Stationary_matrix4_7_0; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_7_1 = my_stationary_io_o_Stationary_matrix4_7_1; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_7_2 = my_stationary_io_o_Stationary_matrix4_7_2; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_7_3 = my_stationary_io_o_Stationary_matrix4_7_3; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_7_4 = my_stationary_io_o_Stationary_matrix4_7_4; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_7_5 = my_stationary_io_o_Stationary_matrix4_7_5; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_7_6 = my_stationary_io_o_Stationary_matrix4_7_6; // @[ivntop.scala 94:34]
  assign my_ivn4_io_Stationary_matrix_7_7 = my_stationary_io_o_Stationary_matrix4_7_7; // @[ivntop.scala 94:34]
  assign my_ivn4_io_validpin = counter >= 32'h28; // @[ivntop.scala 49:16]
  assign my_ivn5_clock = clock;
  assign my_ivn5_reset = reset;
  assign my_ivn5_io_Stationary_matrix_0_0 = my_stationary_io_o_Stationary_matrix5_0_0; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_0_1 = my_stationary_io_o_Stationary_matrix5_0_1; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_0_2 = my_stationary_io_o_Stationary_matrix5_0_2; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_0_3 = my_stationary_io_o_Stationary_matrix5_0_3; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_0_4 = my_stationary_io_o_Stationary_matrix5_0_4; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_0_5 = my_stationary_io_o_Stationary_matrix5_0_5; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_0_6 = my_stationary_io_o_Stationary_matrix5_0_6; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_0_7 = my_stationary_io_o_Stationary_matrix5_0_7; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_1_0 = my_stationary_io_o_Stationary_matrix5_1_0; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_1_1 = my_stationary_io_o_Stationary_matrix5_1_1; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_1_2 = my_stationary_io_o_Stationary_matrix5_1_2; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_1_3 = my_stationary_io_o_Stationary_matrix5_1_3; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_1_4 = my_stationary_io_o_Stationary_matrix5_1_4; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_1_5 = my_stationary_io_o_Stationary_matrix5_1_5; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_1_6 = my_stationary_io_o_Stationary_matrix5_1_6; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_1_7 = my_stationary_io_o_Stationary_matrix5_1_7; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_2_0 = my_stationary_io_o_Stationary_matrix5_2_0; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_2_1 = my_stationary_io_o_Stationary_matrix5_2_1; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_2_2 = my_stationary_io_o_Stationary_matrix5_2_2; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_2_3 = my_stationary_io_o_Stationary_matrix5_2_3; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_2_4 = my_stationary_io_o_Stationary_matrix5_2_4; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_2_5 = my_stationary_io_o_Stationary_matrix5_2_5; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_2_6 = my_stationary_io_o_Stationary_matrix5_2_6; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_2_7 = my_stationary_io_o_Stationary_matrix5_2_7; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_3_0 = my_stationary_io_o_Stationary_matrix5_3_0; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_3_1 = my_stationary_io_o_Stationary_matrix5_3_1; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_3_2 = my_stationary_io_o_Stationary_matrix5_3_2; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_3_3 = my_stationary_io_o_Stationary_matrix5_3_3; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_3_4 = my_stationary_io_o_Stationary_matrix5_3_4; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_3_5 = my_stationary_io_o_Stationary_matrix5_3_5; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_3_6 = my_stationary_io_o_Stationary_matrix5_3_6; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_3_7 = my_stationary_io_o_Stationary_matrix5_3_7; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_4_0 = my_stationary_io_o_Stationary_matrix5_4_0; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_4_1 = my_stationary_io_o_Stationary_matrix5_4_1; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_4_2 = my_stationary_io_o_Stationary_matrix5_4_2; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_4_3 = my_stationary_io_o_Stationary_matrix5_4_3; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_4_4 = my_stationary_io_o_Stationary_matrix5_4_4; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_4_5 = my_stationary_io_o_Stationary_matrix5_4_5; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_4_6 = my_stationary_io_o_Stationary_matrix5_4_6; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_4_7 = my_stationary_io_o_Stationary_matrix5_4_7; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_5_0 = my_stationary_io_o_Stationary_matrix5_5_0; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_5_1 = my_stationary_io_o_Stationary_matrix5_5_1; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_5_2 = my_stationary_io_o_Stationary_matrix5_5_2; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_5_3 = my_stationary_io_o_Stationary_matrix5_5_3; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_5_4 = my_stationary_io_o_Stationary_matrix5_5_4; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_5_5 = my_stationary_io_o_Stationary_matrix5_5_5; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_5_6 = my_stationary_io_o_Stationary_matrix5_5_6; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_5_7 = my_stationary_io_o_Stationary_matrix5_5_7; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_6_0 = my_stationary_io_o_Stationary_matrix5_6_0; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_6_1 = my_stationary_io_o_Stationary_matrix5_6_1; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_6_2 = my_stationary_io_o_Stationary_matrix5_6_2; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_6_3 = my_stationary_io_o_Stationary_matrix5_6_3; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_6_4 = my_stationary_io_o_Stationary_matrix5_6_4; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_6_5 = my_stationary_io_o_Stationary_matrix5_6_5; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_6_6 = my_stationary_io_o_Stationary_matrix5_6_6; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_6_7 = my_stationary_io_o_Stationary_matrix5_6_7; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_7_0 = my_stationary_io_o_Stationary_matrix5_7_0; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_7_1 = my_stationary_io_o_Stationary_matrix5_7_1; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_7_2 = my_stationary_io_o_Stationary_matrix5_7_2; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_7_3 = my_stationary_io_o_Stationary_matrix5_7_3; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_7_4 = my_stationary_io_o_Stationary_matrix5_7_4; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_7_5 = my_stationary_io_o_Stationary_matrix5_7_5; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_7_6 = my_stationary_io_o_Stationary_matrix5_7_6; // @[ivntop.scala 101:34]
  assign my_ivn5_io_Stationary_matrix_7_7 = my_stationary_io_o_Stationary_matrix5_7_7; // @[ivntop.scala 101:34]
  assign my_ivn5_io_validpin = counter >= 32'h32; // @[ivntop.scala 52:16]
  assign my_ivn6_clock = clock;
  assign my_ivn6_reset = reset;
  assign my_ivn6_io_Stationary_matrix_0_0 = my_stationary_io_o_Stationary_matrix6_0_0; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_0_1 = my_stationary_io_o_Stationary_matrix6_0_1; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_0_2 = my_stationary_io_o_Stationary_matrix6_0_2; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_0_3 = my_stationary_io_o_Stationary_matrix6_0_3; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_0_4 = my_stationary_io_o_Stationary_matrix6_0_4; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_0_5 = my_stationary_io_o_Stationary_matrix6_0_5; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_0_6 = my_stationary_io_o_Stationary_matrix6_0_6; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_0_7 = my_stationary_io_o_Stationary_matrix6_0_7; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_1_0 = my_stationary_io_o_Stationary_matrix6_1_0; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_1_1 = my_stationary_io_o_Stationary_matrix6_1_1; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_1_2 = my_stationary_io_o_Stationary_matrix6_1_2; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_1_3 = my_stationary_io_o_Stationary_matrix6_1_3; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_1_4 = my_stationary_io_o_Stationary_matrix6_1_4; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_1_5 = my_stationary_io_o_Stationary_matrix6_1_5; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_1_6 = my_stationary_io_o_Stationary_matrix6_1_6; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_1_7 = my_stationary_io_o_Stationary_matrix6_1_7; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_2_0 = my_stationary_io_o_Stationary_matrix6_2_0; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_2_1 = my_stationary_io_o_Stationary_matrix6_2_1; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_2_2 = my_stationary_io_o_Stationary_matrix6_2_2; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_2_3 = my_stationary_io_o_Stationary_matrix6_2_3; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_2_4 = my_stationary_io_o_Stationary_matrix6_2_4; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_2_5 = my_stationary_io_o_Stationary_matrix6_2_5; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_2_6 = my_stationary_io_o_Stationary_matrix6_2_6; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_2_7 = my_stationary_io_o_Stationary_matrix6_2_7; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_3_0 = my_stationary_io_o_Stationary_matrix6_3_0; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_3_1 = my_stationary_io_o_Stationary_matrix6_3_1; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_3_2 = my_stationary_io_o_Stationary_matrix6_3_2; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_3_3 = my_stationary_io_o_Stationary_matrix6_3_3; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_3_4 = my_stationary_io_o_Stationary_matrix6_3_4; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_3_5 = my_stationary_io_o_Stationary_matrix6_3_5; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_3_6 = my_stationary_io_o_Stationary_matrix6_3_6; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_3_7 = my_stationary_io_o_Stationary_matrix6_3_7; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_4_0 = my_stationary_io_o_Stationary_matrix6_4_0; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_4_1 = my_stationary_io_o_Stationary_matrix6_4_1; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_4_2 = my_stationary_io_o_Stationary_matrix6_4_2; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_4_3 = my_stationary_io_o_Stationary_matrix6_4_3; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_4_4 = my_stationary_io_o_Stationary_matrix6_4_4; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_4_5 = my_stationary_io_o_Stationary_matrix6_4_5; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_4_6 = my_stationary_io_o_Stationary_matrix6_4_6; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_4_7 = my_stationary_io_o_Stationary_matrix6_4_7; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_5_0 = my_stationary_io_o_Stationary_matrix6_5_0; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_5_1 = my_stationary_io_o_Stationary_matrix6_5_1; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_5_2 = my_stationary_io_o_Stationary_matrix6_5_2; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_5_3 = my_stationary_io_o_Stationary_matrix6_5_3; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_5_4 = my_stationary_io_o_Stationary_matrix6_5_4; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_5_5 = my_stationary_io_o_Stationary_matrix6_5_5; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_5_6 = my_stationary_io_o_Stationary_matrix6_5_6; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_5_7 = my_stationary_io_o_Stationary_matrix6_5_7; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_6_0 = my_stationary_io_o_Stationary_matrix6_6_0; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_6_1 = my_stationary_io_o_Stationary_matrix6_6_1; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_6_2 = my_stationary_io_o_Stationary_matrix6_6_2; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_6_3 = my_stationary_io_o_Stationary_matrix6_6_3; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_6_4 = my_stationary_io_o_Stationary_matrix6_6_4; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_6_5 = my_stationary_io_o_Stationary_matrix6_6_5; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_6_6 = my_stationary_io_o_Stationary_matrix6_6_6; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_6_7 = my_stationary_io_o_Stationary_matrix6_6_7; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_7_0 = my_stationary_io_o_Stationary_matrix6_7_0; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_7_1 = my_stationary_io_o_Stationary_matrix6_7_1; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_7_2 = my_stationary_io_o_Stationary_matrix6_7_2; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_7_3 = my_stationary_io_o_Stationary_matrix6_7_3; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_7_4 = my_stationary_io_o_Stationary_matrix6_7_4; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_7_5 = my_stationary_io_o_Stationary_matrix6_7_5; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_7_6 = my_stationary_io_o_Stationary_matrix6_7_6; // @[ivntop.scala 108:34]
  assign my_ivn6_io_Stationary_matrix_7_7 = my_stationary_io_o_Stationary_matrix6_7_7; // @[ivntop.scala 108:34]
  assign my_ivn6_io_validpin = counter >= 32'h3c; // @[ivntop.scala 55:16]
  assign my_ivn7_clock = clock;
  assign my_ivn7_reset = reset;
  assign my_ivn7_io_Stationary_matrix_0_0 = my_stationary_io_o_Stationary_matrix7_0_0; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_0_1 = my_stationary_io_o_Stationary_matrix7_0_1; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_0_2 = my_stationary_io_o_Stationary_matrix7_0_2; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_0_3 = my_stationary_io_o_Stationary_matrix7_0_3; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_0_4 = my_stationary_io_o_Stationary_matrix7_0_4; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_0_5 = my_stationary_io_o_Stationary_matrix7_0_5; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_0_6 = my_stationary_io_o_Stationary_matrix7_0_6; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_0_7 = my_stationary_io_o_Stationary_matrix7_0_7; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_1_0 = my_stationary_io_o_Stationary_matrix7_1_0; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_1_1 = my_stationary_io_o_Stationary_matrix7_1_1; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_1_2 = my_stationary_io_o_Stationary_matrix7_1_2; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_1_3 = my_stationary_io_o_Stationary_matrix7_1_3; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_1_4 = my_stationary_io_o_Stationary_matrix7_1_4; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_1_5 = my_stationary_io_o_Stationary_matrix7_1_5; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_1_6 = my_stationary_io_o_Stationary_matrix7_1_6; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_1_7 = my_stationary_io_o_Stationary_matrix7_1_7; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_2_0 = my_stationary_io_o_Stationary_matrix7_2_0; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_2_1 = my_stationary_io_o_Stationary_matrix7_2_1; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_2_2 = my_stationary_io_o_Stationary_matrix7_2_2; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_2_3 = my_stationary_io_o_Stationary_matrix7_2_3; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_2_4 = my_stationary_io_o_Stationary_matrix7_2_4; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_2_5 = my_stationary_io_o_Stationary_matrix7_2_5; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_2_6 = my_stationary_io_o_Stationary_matrix7_2_6; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_2_7 = my_stationary_io_o_Stationary_matrix7_2_7; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_3_0 = my_stationary_io_o_Stationary_matrix7_3_0; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_3_1 = my_stationary_io_o_Stationary_matrix7_3_1; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_3_2 = my_stationary_io_o_Stationary_matrix7_3_2; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_3_3 = my_stationary_io_o_Stationary_matrix7_3_3; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_3_4 = my_stationary_io_o_Stationary_matrix7_3_4; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_3_5 = my_stationary_io_o_Stationary_matrix7_3_5; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_3_6 = my_stationary_io_o_Stationary_matrix7_3_6; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_3_7 = my_stationary_io_o_Stationary_matrix7_3_7; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_4_0 = my_stationary_io_o_Stationary_matrix7_4_0; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_4_1 = my_stationary_io_o_Stationary_matrix7_4_1; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_4_2 = my_stationary_io_o_Stationary_matrix7_4_2; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_4_3 = my_stationary_io_o_Stationary_matrix7_4_3; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_4_4 = my_stationary_io_o_Stationary_matrix7_4_4; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_4_5 = my_stationary_io_o_Stationary_matrix7_4_5; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_4_6 = my_stationary_io_o_Stationary_matrix7_4_6; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_4_7 = my_stationary_io_o_Stationary_matrix7_4_7; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_5_0 = my_stationary_io_o_Stationary_matrix7_5_0; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_5_1 = my_stationary_io_o_Stationary_matrix7_5_1; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_5_2 = my_stationary_io_o_Stationary_matrix7_5_2; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_5_3 = my_stationary_io_o_Stationary_matrix7_5_3; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_5_4 = my_stationary_io_o_Stationary_matrix7_5_4; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_5_5 = my_stationary_io_o_Stationary_matrix7_5_5; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_5_6 = my_stationary_io_o_Stationary_matrix7_5_6; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_5_7 = my_stationary_io_o_Stationary_matrix7_5_7; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_6_0 = my_stationary_io_o_Stationary_matrix7_6_0; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_6_1 = my_stationary_io_o_Stationary_matrix7_6_1; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_6_2 = my_stationary_io_o_Stationary_matrix7_6_2; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_6_3 = my_stationary_io_o_Stationary_matrix7_6_3; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_6_4 = my_stationary_io_o_Stationary_matrix7_6_4; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_6_5 = my_stationary_io_o_Stationary_matrix7_6_5; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_6_6 = my_stationary_io_o_Stationary_matrix7_6_6; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_6_7 = my_stationary_io_o_Stationary_matrix7_6_7; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_7_0 = my_stationary_io_o_Stationary_matrix7_7_0; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_7_1 = my_stationary_io_o_Stationary_matrix7_7_1; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_7_2 = my_stationary_io_o_Stationary_matrix7_7_2; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_7_3 = my_stationary_io_o_Stationary_matrix7_7_3; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_7_4 = my_stationary_io_o_Stationary_matrix7_7_4; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_7_5 = my_stationary_io_o_Stationary_matrix7_7_5; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_7_6 = my_stationary_io_o_Stationary_matrix7_7_6; // @[ivntop.scala 115:34]
  assign my_ivn7_io_Stationary_matrix_7_7 = my_stationary_io_o_Stationary_matrix7_7_7; // @[ivntop.scala 115:34]
  assign my_ivn7_io_validpin = counter >= 32'h46; // @[ivntop.scala 58:16]
  assign my_ivn8_clock = clock;
  assign my_ivn8_reset = reset;
  assign my_ivn8_io_Stationary_matrix_0_0 = my_stationary_io_o_Stationary_matrix8_0_0; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_0_1 = my_stationary_io_o_Stationary_matrix8_0_1; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_0_2 = my_stationary_io_o_Stationary_matrix8_0_2; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_0_3 = my_stationary_io_o_Stationary_matrix8_0_3; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_0_4 = my_stationary_io_o_Stationary_matrix8_0_4; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_0_5 = my_stationary_io_o_Stationary_matrix8_0_5; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_0_6 = my_stationary_io_o_Stationary_matrix8_0_6; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_0_7 = my_stationary_io_o_Stationary_matrix8_0_7; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_1_0 = my_stationary_io_o_Stationary_matrix8_1_0; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_1_1 = my_stationary_io_o_Stationary_matrix8_1_1; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_1_2 = my_stationary_io_o_Stationary_matrix8_1_2; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_1_3 = my_stationary_io_o_Stationary_matrix8_1_3; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_1_4 = my_stationary_io_o_Stationary_matrix8_1_4; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_1_5 = my_stationary_io_o_Stationary_matrix8_1_5; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_1_6 = my_stationary_io_o_Stationary_matrix8_1_6; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_1_7 = my_stationary_io_o_Stationary_matrix8_1_7; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_2_0 = my_stationary_io_o_Stationary_matrix8_2_0; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_2_1 = my_stationary_io_o_Stationary_matrix8_2_1; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_2_2 = my_stationary_io_o_Stationary_matrix8_2_2; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_2_3 = my_stationary_io_o_Stationary_matrix8_2_3; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_2_4 = my_stationary_io_o_Stationary_matrix8_2_4; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_2_5 = my_stationary_io_o_Stationary_matrix8_2_5; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_2_6 = my_stationary_io_o_Stationary_matrix8_2_6; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_2_7 = my_stationary_io_o_Stationary_matrix8_2_7; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_3_0 = my_stationary_io_o_Stationary_matrix8_3_0; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_3_1 = my_stationary_io_o_Stationary_matrix8_3_1; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_3_2 = my_stationary_io_o_Stationary_matrix8_3_2; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_3_3 = my_stationary_io_o_Stationary_matrix8_3_3; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_3_4 = my_stationary_io_o_Stationary_matrix8_3_4; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_3_5 = my_stationary_io_o_Stationary_matrix8_3_5; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_3_6 = my_stationary_io_o_Stationary_matrix8_3_6; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_3_7 = my_stationary_io_o_Stationary_matrix8_3_7; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_4_0 = my_stationary_io_o_Stationary_matrix8_4_0; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_4_1 = my_stationary_io_o_Stationary_matrix8_4_1; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_4_2 = my_stationary_io_o_Stationary_matrix8_4_2; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_4_3 = my_stationary_io_o_Stationary_matrix8_4_3; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_4_4 = my_stationary_io_o_Stationary_matrix8_4_4; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_4_5 = my_stationary_io_o_Stationary_matrix8_4_5; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_4_6 = my_stationary_io_o_Stationary_matrix8_4_6; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_4_7 = my_stationary_io_o_Stationary_matrix8_4_7; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_5_0 = my_stationary_io_o_Stationary_matrix8_5_0; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_5_1 = my_stationary_io_o_Stationary_matrix8_5_1; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_5_2 = my_stationary_io_o_Stationary_matrix8_5_2; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_5_3 = my_stationary_io_o_Stationary_matrix8_5_3; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_5_4 = my_stationary_io_o_Stationary_matrix8_5_4; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_5_5 = my_stationary_io_o_Stationary_matrix8_5_5; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_5_6 = my_stationary_io_o_Stationary_matrix8_5_6; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_5_7 = my_stationary_io_o_Stationary_matrix8_5_7; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_6_0 = my_stationary_io_o_Stationary_matrix8_6_0; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_6_1 = my_stationary_io_o_Stationary_matrix8_6_1; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_6_2 = my_stationary_io_o_Stationary_matrix8_6_2; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_6_3 = my_stationary_io_o_Stationary_matrix8_6_3; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_6_4 = my_stationary_io_o_Stationary_matrix8_6_4; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_6_5 = my_stationary_io_o_Stationary_matrix8_6_5; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_6_6 = my_stationary_io_o_Stationary_matrix8_6_6; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_6_7 = my_stationary_io_o_Stationary_matrix8_6_7; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_7_0 = my_stationary_io_o_Stationary_matrix8_7_0; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_7_1 = my_stationary_io_o_Stationary_matrix8_7_1; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_7_2 = my_stationary_io_o_Stationary_matrix8_7_2; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_7_3 = my_stationary_io_o_Stationary_matrix8_7_3; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_7_4 = my_stationary_io_o_Stationary_matrix8_7_4; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_7_5 = my_stationary_io_o_Stationary_matrix8_7_5; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_7_6 = my_stationary_io_o_Stationary_matrix8_7_6; // @[ivntop.scala 122:34]
  assign my_ivn8_io_Stationary_matrix_7_7 = my_stationary_io_o_Stationary_matrix8_7_7; // @[ivntop.scala 122:34]
  assign my_ivn8_io_validpin = counter >= 32'h50; // @[ivntop.scala 61:16]
  always @(posedge clock) begin
    i_vn_0_0 <= my_ivn1_io_o_vn_0; // @[ivntop.scala 135:13]
    i_vn_0_1 <= my_ivn1_io_o_vn_1; // @[ivntop.scala 135:13]
    i_vn_0_2 <= my_ivn1_io_o_vn_2; // @[ivntop.scala 135:13]
    i_vn_0_3 <= my_ivn1_io_o_vn_3; // @[ivntop.scala 135:13]
    i_vn_1_0 <= my_ivn1_io_o_vn2_0; // @[ivntop.scala 136:12]
    i_vn_1_1 <= my_ivn1_io_o_vn2_1; // @[ivntop.scala 136:12]
    i_vn_1_2 <= my_ivn1_io_o_vn2_2; // @[ivntop.scala 136:12]
    i_vn_1_3 <= my_ivn1_io_o_vn2_3; // @[ivntop.scala 136:12]
    i_vn_2_0 <= my_ivn2_io_o_vn_0; // @[ivntop.scala 137:13]
    i_vn_2_1 <= my_ivn2_io_o_vn_1; // @[ivntop.scala 137:13]
    i_vn_2_2 <= my_ivn2_io_o_vn_2; // @[ivntop.scala 137:13]
    i_vn_2_3 <= my_ivn2_io_o_vn_3; // @[ivntop.scala 137:13]
    i_vn_3_0 <= my_ivn2_io_o_vn2_0; // @[ivntop.scala 138:13]
    i_vn_3_1 <= my_ivn2_io_o_vn2_1; // @[ivntop.scala 138:13]
    i_vn_3_2 <= my_ivn2_io_o_vn2_2; // @[ivntop.scala 138:13]
    i_vn_3_3 <= my_ivn2_io_o_vn2_3; // @[ivntop.scala 138:13]
    i_vn_4_0 <= my_ivn3_io_o_vn_0; // @[ivntop.scala 139:13]
    i_vn_4_1 <= my_ivn3_io_o_vn_1; // @[ivntop.scala 139:13]
    i_vn_4_2 <= my_ivn3_io_o_vn_2; // @[ivntop.scala 139:13]
    i_vn_4_3 <= my_ivn3_io_o_vn_3; // @[ivntop.scala 139:13]
    i_vn_5_0 <= my_ivn3_io_o_vn2_0; // @[ivntop.scala 140:13]
    i_vn_5_1 <= my_ivn3_io_o_vn2_1; // @[ivntop.scala 140:13]
    i_vn_5_2 <= my_ivn3_io_o_vn2_2; // @[ivntop.scala 140:13]
    i_vn_5_3 <= my_ivn3_io_o_vn2_3; // @[ivntop.scala 140:13]
    i_vn_6_0 <= my_ivn4_io_o_vn_0; // @[ivntop.scala 141:13]
    i_vn_6_1 <= my_ivn4_io_o_vn_1; // @[ivntop.scala 141:13]
    i_vn_6_2 <= my_ivn4_io_o_vn_2; // @[ivntop.scala 141:13]
    i_vn_6_3 <= my_ivn4_io_o_vn_3; // @[ivntop.scala 141:13]
    i_vn_7_0 <= my_ivn4_io_o_vn2_0; // @[ivntop.scala 142:13]
    i_vn_7_1 <= my_ivn4_io_o_vn2_1; // @[ivntop.scala 142:13]
    i_vn_7_2 <= my_ivn4_io_o_vn2_2; // @[ivntop.scala 142:13]
    i_vn_7_3 <= my_ivn4_io_o_vn2_3; // @[ivntop.scala 142:13]
    i_vn_8_0 <= my_ivn5_io_o_vn_0; // @[ivntop.scala 143:13]
    i_vn_8_1 <= my_ivn5_io_o_vn_1; // @[ivntop.scala 143:13]
    i_vn_8_2 <= my_ivn5_io_o_vn_2; // @[ivntop.scala 143:13]
    i_vn_8_3 <= my_ivn5_io_o_vn_3; // @[ivntop.scala 143:13]
    i_vn_9_0 <= my_ivn5_io_o_vn2_0; // @[ivntop.scala 144:13]
    i_vn_9_1 <= my_ivn5_io_o_vn2_1; // @[ivntop.scala 144:13]
    i_vn_9_2 <= my_ivn5_io_o_vn2_2; // @[ivntop.scala 144:13]
    i_vn_9_3 <= my_ivn5_io_o_vn2_3; // @[ivntop.scala 144:13]
    i_vn_10_0 <= my_ivn6_io_o_vn_0; // @[ivntop.scala 145:14]
    i_vn_10_1 <= my_ivn6_io_o_vn_1; // @[ivntop.scala 145:14]
    i_vn_10_2 <= my_ivn6_io_o_vn_2; // @[ivntop.scala 145:14]
    i_vn_10_3 <= my_ivn6_io_o_vn_3; // @[ivntop.scala 145:14]
    i_vn_11_0 <= my_ivn6_io_o_vn2_0; // @[ivntop.scala 146:13]
    i_vn_11_1 <= my_ivn6_io_o_vn2_1; // @[ivntop.scala 146:13]
    i_vn_11_2 <= my_ivn6_io_o_vn2_2; // @[ivntop.scala 146:13]
    i_vn_11_3 <= my_ivn6_io_o_vn2_3; // @[ivntop.scala 146:13]
    i_vn_12_0 <= my_ivn7_io_o_vn_0; // @[ivntop.scala 147:14]
    i_vn_12_1 <= my_ivn7_io_o_vn_1; // @[ivntop.scala 147:14]
    i_vn_12_2 <= my_ivn7_io_o_vn_2; // @[ivntop.scala 147:14]
    i_vn_12_3 <= my_ivn7_io_o_vn_3; // @[ivntop.scala 147:14]
    i_vn_13_0 <= my_ivn7_io_o_vn2_0; // @[ivntop.scala 148:14]
    i_vn_13_1 <= my_ivn7_io_o_vn2_1; // @[ivntop.scala 148:14]
    i_vn_13_2 <= my_ivn7_io_o_vn2_2; // @[ivntop.scala 148:14]
    i_vn_13_3 <= my_ivn7_io_o_vn2_3; // @[ivntop.scala 148:14]
    i_vn_14_0 <= my_ivn8_io_o_vn_0; // @[ivntop.scala 149:14]
    i_vn_14_1 <= my_ivn8_io_o_vn_1; // @[ivntop.scala 149:14]
    i_vn_14_2 <= my_ivn8_io_o_vn_2; // @[ivntop.scala 149:14]
    i_vn_14_3 <= my_ivn8_io_o_vn_3; // @[ivntop.scala 149:14]
    i_vn_15_0 <= my_ivn8_io_o_vn2_0; // @[ivntop.scala 150:14]
    i_vn_15_1 <= my_ivn8_io_o_vn2_1; // @[ivntop.scala 150:14]
    i_vn_15_2 <= my_ivn8_io_o_vn2_2; // @[ivntop.scala 150:14]
    i_vn_15_3 <= my_ivn8_io_o_vn2_3; // @[ivntop.scala 150:14]
    if (reset) begin // @[ivntop.scala 27:26]
      counter <= 32'h0; // @[ivntop.scala 27:26]
    end else begin
      counter <= _counter_T_1; // @[ivntop.scala 156:11]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  i_vn_0_0 = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  i_vn_0_1 = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  i_vn_0_2 = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  i_vn_0_3 = _RAND_3[4:0];
  _RAND_4 = {1{`RANDOM}};
  i_vn_1_0 = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  i_vn_1_1 = _RAND_5[4:0];
  _RAND_6 = {1{`RANDOM}};
  i_vn_1_2 = _RAND_6[4:0];
  _RAND_7 = {1{`RANDOM}};
  i_vn_1_3 = _RAND_7[4:0];
  _RAND_8 = {1{`RANDOM}};
  i_vn_2_0 = _RAND_8[4:0];
  _RAND_9 = {1{`RANDOM}};
  i_vn_2_1 = _RAND_9[4:0];
  _RAND_10 = {1{`RANDOM}};
  i_vn_2_2 = _RAND_10[4:0];
  _RAND_11 = {1{`RANDOM}};
  i_vn_2_3 = _RAND_11[4:0];
  _RAND_12 = {1{`RANDOM}};
  i_vn_3_0 = _RAND_12[4:0];
  _RAND_13 = {1{`RANDOM}};
  i_vn_3_1 = _RAND_13[4:0];
  _RAND_14 = {1{`RANDOM}};
  i_vn_3_2 = _RAND_14[4:0];
  _RAND_15 = {1{`RANDOM}};
  i_vn_3_3 = _RAND_15[4:0];
  _RAND_16 = {1{`RANDOM}};
  i_vn_4_0 = _RAND_16[4:0];
  _RAND_17 = {1{`RANDOM}};
  i_vn_4_1 = _RAND_17[4:0];
  _RAND_18 = {1{`RANDOM}};
  i_vn_4_2 = _RAND_18[4:0];
  _RAND_19 = {1{`RANDOM}};
  i_vn_4_3 = _RAND_19[4:0];
  _RAND_20 = {1{`RANDOM}};
  i_vn_5_0 = _RAND_20[4:0];
  _RAND_21 = {1{`RANDOM}};
  i_vn_5_1 = _RAND_21[4:0];
  _RAND_22 = {1{`RANDOM}};
  i_vn_5_2 = _RAND_22[4:0];
  _RAND_23 = {1{`RANDOM}};
  i_vn_5_3 = _RAND_23[4:0];
  _RAND_24 = {1{`RANDOM}};
  i_vn_6_0 = _RAND_24[4:0];
  _RAND_25 = {1{`RANDOM}};
  i_vn_6_1 = _RAND_25[4:0];
  _RAND_26 = {1{`RANDOM}};
  i_vn_6_2 = _RAND_26[4:0];
  _RAND_27 = {1{`RANDOM}};
  i_vn_6_3 = _RAND_27[4:0];
  _RAND_28 = {1{`RANDOM}};
  i_vn_7_0 = _RAND_28[4:0];
  _RAND_29 = {1{`RANDOM}};
  i_vn_7_1 = _RAND_29[4:0];
  _RAND_30 = {1{`RANDOM}};
  i_vn_7_2 = _RAND_30[4:0];
  _RAND_31 = {1{`RANDOM}};
  i_vn_7_3 = _RAND_31[4:0];
  _RAND_32 = {1{`RANDOM}};
  i_vn_8_0 = _RAND_32[4:0];
  _RAND_33 = {1{`RANDOM}};
  i_vn_8_1 = _RAND_33[4:0];
  _RAND_34 = {1{`RANDOM}};
  i_vn_8_2 = _RAND_34[4:0];
  _RAND_35 = {1{`RANDOM}};
  i_vn_8_3 = _RAND_35[4:0];
  _RAND_36 = {1{`RANDOM}};
  i_vn_9_0 = _RAND_36[4:0];
  _RAND_37 = {1{`RANDOM}};
  i_vn_9_1 = _RAND_37[4:0];
  _RAND_38 = {1{`RANDOM}};
  i_vn_9_2 = _RAND_38[4:0];
  _RAND_39 = {1{`RANDOM}};
  i_vn_9_3 = _RAND_39[4:0];
  _RAND_40 = {1{`RANDOM}};
  i_vn_10_0 = _RAND_40[4:0];
  _RAND_41 = {1{`RANDOM}};
  i_vn_10_1 = _RAND_41[4:0];
  _RAND_42 = {1{`RANDOM}};
  i_vn_10_2 = _RAND_42[4:0];
  _RAND_43 = {1{`RANDOM}};
  i_vn_10_3 = _RAND_43[4:0];
  _RAND_44 = {1{`RANDOM}};
  i_vn_11_0 = _RAND_44[4:0];
  _RAND_45 = {1{`RANDOM}};
  i_vn_11_1 = _RAND_45[4:0];
  _RAND_46 = {1{`RANDOM}};
  i_vn_11_2 = _RAND_46[4:0];
  _RAND_47 = {1{`RANDOM}};
  i_vn_11_3 = _RAND_47[4:0];
  _RAND_48 = {1{`RANDOM}};
  i_vn_12_0 = _RAND_48[4:0];
  _RAND_49 = {1{`RANDOM}};
  i_vn_12_1 = _RAND_49[4:0];
  _RAND_50 = {1{`RANDOM}};
  i_vn_12_2 = _RAND_50[4:0];
  _RAND_51 = {1{`RANDOM}};
  i_vn_12_3 = _RAND_51[4:0];
  _RAND_52 = {1{`RANDOM}};
  i_vn_13_0 = _RAND_52[4:0];
  _RAND_53 = {1{`RANDOM}};
  i_vn_13_1 = _RAND_53[4:0];
  _RAND_54 = {1{`RANDOM}};
  i_vn_13_2 = _RAND_54[4:0];
  _RAND_55 = {1{`RANDOM}};
  i_vn_13_3 = _RAND_55[4:0];
  _RAND_56 = {1{`RANDOM}};
  i_vn_14_0 = _RAND_56[4:0];
  _RAND_57 = {1{`RANDOM}};
  i_vn_14_1 = _RAND_57[4:0];
  _RAND_58 = {1{`RANDOM}};
  i_vn_14_2 = _RAND_58[4:0];
  _RAND_59 = {1{`RANDOM}};
  i_vn_14_3 = _RAND_59[4:0];
  _RAND_60 = {1{`RANDOM}};
  i_vn_15_0 = _RAND_60[4:0];
  _RAND_61 = {1{`RANDOM}};
  i_vn_15_1 = _RAND_61[4:0];
  _RAND_62 = {1{`RANDOM}};
  i_vn_15_2 = _RAND_62[4:0];
  _RAND_63 = {1{`RANDOM}};
  i_vn_15_3 = _RAND_63[4:0];
  _RAND_64 = {1{`RANDOM}};
  counter = _RAND_64[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MuxesWrapper(
  input         io_valid,
  input  [31:0] io_src_0,
  input  [31:0] io_src_1,
  input  [31:0] io_src_2,
  input  [31:0] io_src_3,
  input  [31:0] io_muxes_0,
  input  [31:0] io_muxes_1,
  input  [31:0] io_muxes_2,
  input  [31:0] io_muxes_3,
  output [31:0] io_Osrc_0,
  output [31:0] io_Osrc_1,
  output [31:0] io_Osrc_2,
  output [31:0] io_Osrc_3,
  output [31:0] io_Omuxes_0_0,
  output [31:0] io_Omuxes_0_1,
  output [31:0] io_Omuxes_0_2,
  output [31:0] io_Omuxes_0_3,
  output [31:0] io_Omuxes_1_0,
  output [31:0] io_Omuxes_1_1,
  output [31:0] io_Omuxes_1_2,
  output [31:0] io_Omuxes_2_0,
  output [31:0] io_Omuxes_2_1,
  output [31:0] io_Omuxes_3_0
);
  wire  _T = io_src_0 != io_src_1; // @[MuxesWrapper.scala 24:25]
  wire [31:0] _GEN_108 = {{31'd0}, io_src_0 != io_src_1}; // @[MuxesWrapper.scala 24:39]
  wire [31:0] _GEN_109 = {{31'd0}, _GEN_108 != io_src_2}; // @[MuxesWrapper.scala 24:53]
  wire [31:0] _GEN_0 = _GEN_109 != io_src_3 ? io_src_0 : 32'h0; // @[MuxesWrapper.scala 24:67 25:17]
  wire [31:0] _GEN_1 = _GEN_109 != io_src_3 ? io_src_1 : 32'h0; // @[MuxesWrapper.scala 24:67 25:17]
  wire [31:0] _GEN_2 = _GEN_109 != io_src_3 ? io_src_2 : 32'h0; // @[MuxesWrapper.scala 24:67 25:17]
  wire [31:0] _GEN_3 = _GEN_109 != io_src_3 ? io_src_3 : 32'h0; // @[MuxesWrapper.scala 24:67 25:17]
  wire [31:0] _GEN_4 = _GEN_109 != io_src_3 ? io_muxes_0 : 32'h0; // @[MuxesWrapper.scala 24:67 26:23]
  wire [31:0] _GEN_5 = _GEN_109 != io_src_3 ? io_muxes_1 : 32'h0; // @[MuxesWrapper.scala 24:67 27:23]
  wire [31:0] _GEN_6 = _GEN_109 != io_src_3 ? io_muxes_2 : 32'h0; // @[MuxesWrapper.scala 24:67 28:23]
  wire [31:0] _GEN_7 = _GEN_109 != io_src_3 ? io_muxes_3 : 32'h0; // @[MuxesWrapper.scala 24:67 29:23]
  wire  _T_4 = io_src_1 != io_src_2; // @[MuxesWrapper.scala 31:56]
  wire  _T_6 = io_src_2 == io_src_3; // @[MuxesWrapper.scala 31:85]
  wire [31:0] _GEN_8 = _T & io_src_1 != io_src_2 & io_src_2 == io_src_3 ? 32'h0 : _GEN_3; // @[MuxesWrapper.scala 31:100 32:20]
  wire [31:0] _GEN_9 = _T & io_src_1 != io_src_2 & io_src_2 == io_src_3 ? io_src_2 : _GEN_2; // @[MuxesWrapper.scala 31:100 33:20]
  wire [31:0] _GEN_10 = _T & io_src_1 != io_src_2 & io_src_2 == io_src_3 ? io_src_1 : _GEN_1; // @[MuxesWrapper.scala 31:100 34:20]
  wire [31:0] _GEN_11 = _T & io_src_1 != io_src_2 & io_src_2 == io_src_3 ? io_src_0 : _GEN_0; // @[MuxesWrapper.scala 31:100 35:20]
  wire [31:0] _GEN_12 = _T & io_src_1 != io_src_2 & io_src_2 == io_src_3 ? io_muxes_0 : _GEN_4; // @[MuxesWrapper.scala 31:100 36:23]
  wire [31:0] _GEN_13 = _T & io_src_1 != io_src_2 & io_src_2 == io_src_3 ? io_muxes_1 : _GEN_5; // @[MuxesWrapper.scala 31:100 37:23]
  wire [31:0] _GEN_14 = _T & io_src_1 != io_src_2 & io_src_2 == io_src_3 ? io_muxes_2 : _GEN_6; // @[MuxesWrapper.scala 31:100 38:23]
  wire [31:0] _GEN_15 = _T & io_src_1 != io_src_2 & io_src_2 == io_src_3 ? io_muxes_3 : 32'h0; // @[MuxesWrapper.scala 31:100 39:23]
  wire [31:0] _GEN_16 = _T & io_src_1 != io_src_2 & io_src_2 == io_src_3 ? 32'h0 : _GEN_7; // @[MuxesWrapper.scala 31:100 40:23]
  wire  _T_8 = io_src_0 == io_src_1; // @[MuxesWrapper.scala 44:30]
  wire  _T_10 = io_src_0 == io_src_1 & _T_4; // @[MuxesWrapper.scala 44:45]
  wire [31:0] _GEN_17 = io_src_0 == io_src_1 & _T_4 & _T_6 ? io_src_2 : _GEN_9; // @[MuxesWrapper.scala 44:104 45:20]
  wire [31:0] _GEN_18 = io_src_0 == io_src_1 & _T_4 & _T_6 ? io_src_0 : _GEN_11; // @[MuxesWrapper.scala 44:104 46:20]
  wire [31:0] _GEN_19 = io_src_0 == io_src_1 & _T_4 & _T_6 ? 32'h0 : _GEN_10; // @[MuxesWrapper.scala 44:104 47:20]
  wire [31:0] _GEN_20 = io_src_0 == io_src_1 & _T_4 & _T_6 ? 32'h0 : _GEN_8; // @[MuxesWrapper.scala 44:104 48:20]
  wire [31:0] _GEN_21 = io_src_0 == io_src_1 & _T_4 & _T_6 ? io_muxes_0 : _GEN_12; // @[MuxesWrapper.scala 44:104 49:23]
  wire [31:0] _GEN_22 = io_src_0 == io_src_1 & _T_4 & _T_6 ? io_muxes_1 : 32'h0; // @[MuxesWrapper.scala 44:104 50:23]
  wire [31:0] _GEN_23 = io_src_0 == io_src_1 & _T_4 & _T_6 ? io_muxes_2 : _GEN_14; // @[MuxesWrapper.scala 44:104 51:23]
  wire [31:0] _GEN_24 = io_src_0 == io_src_1 & _T_4 & _T_6 ? io_muxes_3 : _GEN_15; // @[MuxesWrapper.scala 44:104 52:23]
  wire  _T_16 = io_src_2 != io_src_3; // @[MuxesWrapper.scala 55:85]
  wire [31:0] _GEN_25 = _T_10 & io_src_2 != io_src_3 ? io_src_3 : _GEN_20; // @[MuxesWrapper.scala 55:100 56:20]
  wire [31:0] _GEN_26 = _T_10 & io_src_2 != io_src_3 ? io_src_2 : _GEN_17; // @[MuxesWrapper.scala 55:100 57:20]
  wire [31:0] _GEN_27 = _T_10 & io_src_2 != io_src_3 ? 32'h0 : _GEN_19; // @[MuxesWrapper.scala 55:100 58:20]
  wire [31:0] _GEN_28 = _T_10 & io_src_2 != io_src_3 ? io_src_0 : _GEN_18; // @[MuxesWrapper.scala 55:100 59:20]
  wire [31:0] _GEN_29 = _T_10 & io_src_2 != io_src_3 ? io_muxes_0 : _GEN_21; // @[MuxesWrapper.scala 55:100 60:23]
  wire [31:0] _GEN_30 = _T_10 & io_src_2 != io_src_3 ? io_muxes_1 : _GEN_22; // @[MuxesWrapper.scala 55:100 61:23]
  wire [31:0] _GEN_31 = _T_10 & io_src_2 != io_src_3 ? 32'h0 : _GEN_13; // @[MuxesWrapper.scala 55:100 62:23]
  wire [31:0] _GEN_32 = _T_10 & io_src_2 != io_src_3 ? io_muxes_2 : _GEN_23; // @[MuxesWrapper.scala 55:100 63:23]
  wire [31:0] _GEN_33 = _T_10 & io_src_2 != io_src_3 ? 32'h0 : _GEN_16; // @[MuxesWrapper.scala 55:100 64:23]
  wire  _T_19 = io_src_1 == io_src_2; // @[MuxesWrapper.scala 75:60]
  wire  _T_20 = _T & io_src_1 == io_src_2; // @[MuxesWrapper.scala 75:45]
  wire [31:0] _GEN_34 = _T & io_src_1 == io_src_2 & _T_16 ? 32'h0 : _GEN_26; // @[MuxesWrapper.scala 75:104 76:20]
  wire [31:0] _GEN_35 = _T & io_src_1 == io_src_2 & _T_16 ? io_src_3 : _GEN_25; // @[MuxesWrapper.scala 75:104 77:20]
  wire [31:0] _GEN_36 = _T & io_src_1 == io_src_2 & _T_16 ? io_src_1 : _GEN_27; // @[MuxesWrapper.scala 75:104 78:20]
  wire [31:0] _GEN_37 = _T & io_src_1 == io_src_2 & _T_16 ? io_src_0 : _GEN_28; // @[MuxesWrapper.scala 75:104 79:20]
  wire [31:0] _GEN_38 = _T & io_src_1 == io_src_2 & _T_16 ? io_muxes_0 : _GEN_29; // @[MuxesWrapper.scala 75:104 80:23]
  wire [31:0] _GEN_39 = _T & io_src_1 == io_src_2 & _T_16 ? io_muxes_1 : _GEN_31; // @[MuxesWrapper.scala 75:104 81:23]
  wire [31:0] _GEN_40 = _T & io_src_1 == io_src_2 & _T_16 ? io_muxes_2 : 32'h0; // @[MuxesWrapper.scala 75:104 82:23]
  wire [31:0] _GEN_41 = _T & io_src_1 == io_src_2 & _T_16 ? 32'h0 : _GEN_32; // @[MuxesWrapper.scala 75:104 83:23]
  wire [31:0] _GEN_42 = _T & io_src_1 == io_src_2 & _T_16 ? io_muxes_3 : _GEN_33; // @[MuxesWrapper.scala 75:104 84:23]
  wire [31:0] _GEN_43 = _T_20 & _T_6 ? 32'h0 : _GEN_34; // @[MuxesWrapper.scala 94:100 95:20]
  wire [31:0] _GEN_44 = _T_20 & _T_6 ? 32'h0 : _GEN_35; // @[MuxesWrapper.scala 94:100 96:20]
  wire [31:0] _GEN_45 = _T_20 & _T_6 ? io_src_1 : _GEN_36; // @[MuxesWrapper.scala 94:100 97:20]
  wire [31:0] _GEN_46 = _T_20 & _T_6 ? io_src_0 : _GEN_37; // @[MuxesWrapper.scala 94:100 98:20]
  wire [31:0] _GEN_47 = _T_20 & _T_6 ? io_muxes_0 : _GEN_38; // @[MuxesWrapper.scala 94:100 99:23]
  wire [31:0] _GEN_48 = _T_20 & _T_6 ? io_muxes_1 : _GEN_39; // @[MuxesWrapper.scala 94:100 100:23]
  wire [31:0] _GEN_49 = _T_20 & _T_6 ? io_muxes_2 : _GEN_40; // @[MuxesWrapper.scala 94:100 101:23]
  wire [31:0] _GEN_50 = _T_20 & _T_6 ? io_muxes_3 : 32'h0; // @[MuxesWrapper.scala 94:100 102:23]
  wire [31:0] _GEN_51 = _T_20 & _T_6 ? 32'h0 : _GEN_41; // @[MuxesWrapper.scala 94:100 103:23]
  wire [31:0] _GEN_52 = _T_20 & _T_6 ? 32'h0 : _GEN_42; // @[MuxesWrapper.scala 94:100 104:23]
  wire  _T_30 = _T_8 & _T_19; // @[MuxesWrapper.scala 114:41]
  wire [31:0] _GEN_53 = _T_8 & _T_19 & _T_16 ? 32'h0 : _GEN_43; // @[MuxesWrapper.scala 114:100 115:20]
  wire [31:0] _GEN_54 = _T_8 & _T_19 & _T_16 ? io_src_3 : _GEN_44; // @[MuxesWrapper.scala 114:100 116:20]
  wire [31:0] _GEN_55 = _T_8 & _T_19 & _T_16 ? 32'h0 : _GEN_45; // @[MuxesWrapper.scala 114:100 117:20]
  wire [31:0] _GEN_56 = _T_8 & _T_19 & _T_16 ? io_src_0 : _GEN_46; // @[MuxesWrapper.scala 114:100 118:20]
  wire [31:0] _GEN_57 = _T_8 & _T_19 & _T_16 ? io_muxes_0 : _GEN_47; // @[MuxesWrapper.scala 114:100 119:23]
  wire [31:0] _GEN_58 = _T_8 & _T_19 & _T_16 ? io_muxes_1 : _GEN_30; // @[MuxesWrapper.scala 114:100 120:23]
  wire [31:0] _GEN_59 = _T_8 & _T_19 & _T_16 ? io_muxes_2 : 32'h0; // @[MuxesWrapper.scala 114:100 121:23]
  wire [31:0] _GEN_60 = _T_8 & _T_19 & _T_16 ? 32'h0 : _GEN_48; // @[MuxesWrapper.scala 114:100 122:23]
  wire [31:0] _GEN_61 = _T_8 & _T_19 & _T_16 ? 32'h0 : _GEN_51; // @[MuxesWrapper.scala 114:100 123:23]
  wire [31:0] _GEN_62 = _T_8 & _T_19 & _T_16 ? io_muxes_3 : _GEN_52; // @[MuxesWrapper.scala 114:100 124:23]
  wire [31:0] _GEN_63 = _T_30 & _T_6 ? 32'h0 : _GEN_53; // @[MuxesWrapper.scala 136:100 137:20]
  wire [31:0] _GEN_64 = _T_30 & _T_6 ? 32'h0 : _GEN_54; // @[MuxesWrapper.scala 136:100 138:20]
  wire [31:0] _GEN_65 = _T_30 & _T_6 ? 32'h0 : _GEN_55; // @[MuxesWrapper.scala 136:100 139:20]
  wire [31:0] _GEN_66 = _T_30 & _T_6 ? io_src_0 : _GEN_56; // @[MuxesWrapper.scala 136:100 140:20]
  wire [31:0] _GEN_67 = _T_30 & _T_6 ? io_muxes_0 : _GEN_57; // @[MuxesWrapper.scala 136:100 141:23]
  wire [31:0] _GEN_68 = _T_30 & _T_6 ? io_muxes_1 : _GEN_58; // @[MuxesWrapper.scala 136:100 142:23]
  wire [31:0] _GEN_69 = _T_30 & _T_6 ? io_muxes_2 : _GEN_59; // @[MuxesWrapper.scala 136:100 143:23]
  wire [31:0] _GEN_70 = _T_30 & _T_6 ? io_muxes_3 : 32'h0; // @[MuxesWrapper.scala 136:100 144:23]
  wire [31:0] _GEN_71 = _T_30 & _T_6 ? 32'h0 : _GEN_60; // @[MuxesWrapper.scala 136:100 145:23]
  wire [31:0] _GEN_72 = _T_30 & _T_6 ? 32'h0 : _GEN_61; // @[MuxesWrapper.scala 136:100 146:23]
  wire [31:0] _GEN_73 = _T_30 & _T_6 ? 32'h0 : _GEN_62; // @[MuxesWrapper.scala 136:100 147:23]
  wire [31:0] mat_0_0 = io_valid ? _GEN_67 : 32'h0; // @[MuxesWrapper.scala 21:20]
  wire [31:0] mat_0_1 = io_valid ? _GEN_68 : 32'h0; // @[MuxesWrapper.scala 21:20]
  wire [31:0] mat_0_2 = io_valid ? _GEN_69 : 32'h0; // @[MuxesWrapper.scala 21:20]
  wire [31:0] mat_0_3 = io_valid ? _GEN_70 : 32'h0; // @[MuxesWrapper.scala 21:20]
  wire [31:0] mat_1_0 = io_valid ? _GEN_71 : 32'h0; // @[MuxesWrapper.scala 21:20]
  wire [31:0] mat_1_1 = io_valid ? _GEN_49 : 32'h0; // @[MuxesWrapper.scala 21:20]
  wire [31:0] mat_1_2 = io_valid ? _GEN_50 : 32'h0; // @[MuxesWrapper.scala 21:20]
  wire [31:0] mat_2_0 = io_valid ? _GEN_72 : 32'h0; // @[MuxesWrapper.scala 21:20]
  wire [31:0] mat_2_1 = io_valid ? _GEN_24 : 32'h0; // @[MuxesWrapper.scala 21:20]
  wire [31:0] mat_3_0 = io_valid ? _GEN_73 : 32'h0; // @[MuxesWrapper.scala 21:20]
  wire [31:0] src_0 = io_valid ? _GEN_66 : 32'h0; // @[MuxesWrapper.scala 21:20]
  wire [31:0] src_1 = io_valid ? _GEN_65 : 32'h0; // @[MuxesWrapper.scala 21:20]
  wire [31:0] src_2 = io_valid ? _GEN_63 : 32'h0; // @[MuxesWrapper.scala 21:20]
  wire [31:0] src_3 = io_valid ? _GEN_64 : 32'h0; // @[MuxesWrapper.scala 21:20]
  assign io_Osrc_0 = io_valid ? src_0 : 32'h0; // @[MuxesWrapper.scala 163:17 21:20 23:17]
  assign io_Osrc_1 = io_valid ? src_1 : 32'h0; // @[MuxesWrapper.scala 163:17 21:20 23:17]
  assign io_Osrc_2 = io_valid ? src_2 : 32'h0; // @[MuxesWrapper.scala 163:17 21:20 23:17]
  assign io_Osrc_3 = io_valid ? src_3 : 32'h0; // @[MuxesWrapper.scala 163:17 21:20 23:17]
  assign io_Omuxes_0_0 = io_valid ? mat_0_0 : 32'h0; // @[MuxesWrapper.scala 162:19 21:20 22:19]
  assign io_Omuxes_0_1 = io_valid ? mat_0_1 : 32'h0; // @[MuxesWrapper.scala 162:19 21:20 22:19]
  assign io_Omuxes_0_2 = io_valid ? mat_0_2 : 32'h0; // @[MuxesWrapper.scala 162:19 21:20 22:19]
  assign io_Omuxes_0_3 = io_valid ? mat_0_3 : 32'h0; // @[MuxesWrapper.scala 162:19 21:20 22:19]
  assign io_Omuxes_1_0 = io_valid ? mat_1_0 : 32'h0; // @[MuxesWrapper.scala 162:19 21:20 22:19]
  assign io_Omuxes_1_1 = io_valid ? mat_1_1 : 32'h0; // @[MuxesWrapper.scala 162:19 21:20 22:19]
  assign io_Omuxes_1_2 = io_valid ? mat_1_2 : 32'h0; // @[MuxesWrapper.scala 162:19 21:20 22:19]
  assign io_Omuxes_2_0 = io_valid ? mat_2_0 : 32'h0; // @[MuxesWrapper.scala 162:19 21:20 22:19]
  assign io_Omuxes_2_1 = io_valid ? mat_2_1 : 32'h0; // @[MuxesWrapper.scala 162:19 21:20 22:19]
  assign io_Omuxes_3_0 = io_valid ? mat_3_0 : 32'h0; // @[MuxesWrapper.scala 162:19 21:20 22:19]
endmodule
module fancontrol4(
  input        clock,
  input        reset,
  input  [4:0] io_i_vn_0,
  input  [4:0] io_i_vn_1,
  input  [4:0] io_i_vn_2,
  input  [4:0] io_i_vn_3,
  input        io_i_data_valid,
  output       io_o_reduction_add_0,
  output       io_o_reduction_add_1,
  output       io_o_reduction_add_2,
  output [2:0] io_o_reduction_cmd_0,
  output [2:0] io_o_reduction_cmd_1,
  output [2:0] io_o_reduction_cmd_2,
  output       io_o_reduction_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
`endif // RANDOMIZE_REG_INIT
  reg  r_reduction_add_0; // @[FanCtrl.scala 19:34]
  reg  r_reduction_add_1; // @[FanCtrl.scala 19:34]
  reg  r_reduction_add_2; // @[FanCtrl.scala 19:34]
  reg [2:0] r_reduction_cmd_0; // @[FanCtrl.scala 20:34]
  reg [2:0] r_reduction_cmd_1; // @[FanCtrl.scala 20:34]
  reg [2:0] r_reduction_cmd_2; // @[FanCtrl.scala 20:34]
  reg  r_add_lvl_0Reg_6; // @[FanCtrl.scala 23:33]
  reg  r_add_lvl_0Reg_7; // @[FanCtrl.scala 23:33]
  reg  r_add_lvl_1Reg_4; // @[FanCtrl.scala 24:33]
  reg [2:0] r_cmd_lvl_0Reg_6; // @[FanCtrl.scala 27:33]
  reg [2:0] r_cmd_lvl_0Reg_7; // @[FanCtrl.scala 27:33]
  reg [2:0] r_cmd_lvl_1Reg_4; // @[FanCtrl.scala 28:33]
  reg [4:0] w_vn_0; // @[FanCtrl.scala 34:23]
  reg [4:0] w_vn_1; // @[FanCtrl.scala 34:23]
  reg [4:0] w_vn_2; // @[FanCtrl.scala 34:23]
  reg [4:0] w_vn_3; // @[FanCtrl.scala 34:23]
  reg  r_valid_0; // @[FanCtrl.scala 35:26]
  reg  r_valid_1; // @[FanCtrl.scala 35:26]
  reg  r_valid_2; // @[FanCtrl.scala 35:26]
  reg  r_valid_3; // @[FanCtrl.scala 35:26]
  wire [2:0] _T_2 = 2'h2 * 1'h0; // @[FanCtrl.scala 42:25]
  wire [3:0] _T_3 = {{1'd0}, _T_2}; // @[FanCtrl.scala 42:31]
  wire [2:0] _T_8 = _T_2 + 3'h1; // @[FanCtrl.scala 42:58]
  wire [4:0] _GEN_1 = 2'h1 == _T_3[1:0] ? w_vn_1 : w_vn_0; // @[FanCtrl.scala 42:{39,39}]
  wire [4:0] _GEN_2 = 2'h2 == _T_3[1:0] ? w_vn_2 : _GEN_1; // @[FanCtrl.scala 42:{39,39}]
  wire [4:0] _GEN_3 = 2'h3 == _T_3[1:0] ? w_vn_3 : _GEN_2; // @[FanCtrl.scala 42:{39,39}]
  wire [4:0] _GEN_5 = 2'h1 == _T_8[1:0] ? w_vn_1 : w_vn_0; // @[FanCtrl.scala 42:{39,39}]
  wire [4:0] _GEN_6 = 2'h2 == _T_8[1:0] ? w_vn_2 : _GEN_5; // @[FanCtrl.scala 42:{39,39}]
  wire [4:0] _GEN_7 = 2'h3 == _T_8[1:0] ? w_vn_3 : _GEN_6; // @[FanCtrl.scala 42:{39,39}]
  wire  _T_10 = _GEN_3 == _GEN_7; // @[FanCtrl.scala 42:39]
  wire [2:0] _T_21 = _T_2 + 3'h2; // @[FanCtrl.scala 49:32]
  wire [4:0] _GEN_22 = 2'h1 == _T_21[1:0] ? w_vn_1 : w_vn_0; // @[FanCtrl.scala 48:{41,41}]
  wire [4:0] _GEN_23 = 2'h2 == _T_21[1:0] ? w_vn_2 : _GEN_22; // @[FanCtrl.scala 48:{41,41}]
  wire [4:0] _GEN_24 = 2'h3 == _T_21[1:0] ? w_vn_3 : _GEN_23; // @[FanCtrl.scala 48:{41,41}]
  wire  _T_23 = _GEN_7 != _GEN_24; // @[FanCtrl.scala 48:41]
  wire  _T_32 = _GEN_3 != _GEN_7; // @[FanCtrl.scala 50:41]
  wire  _T_33 = _T_23 & _T_32; // @[FanCtrl.scala 49:41]
  wire  _T_42 = _GEN_7 == _GEN_24; // @[FanCtrl.scala 55:48]
  wire  _T_52 = _T_42 & _T_32; // @[FanCtrl.scala 56:46]
  wire [1:0] _GEN_49 = _T_52 ? 2'h3 : 2'h0; // @[FanCtrl.scala 58:48 60:40 63:38]
  wire  _GEN_54 = r_valid_1 & _T_10; // @[FanCtrl.scala 41:34]
  wire [2:0] _T_113 = 2'h2 * 1'h1; // @[FanCtrl.scala 42:25]
  wire [3:0] _T_114 = {{1'd0}, _T_113}; // @[FanCtrl.scala 42:31]
  wire [2:0] _T_119 = _T_113 + 3'h1; // @[FanCtrl.scala 42:58]
  wire [4:0] _GEN_124 = 2'h1 == _T_114[1:0] ? w_vn_1 : w_vn_0; // @[FanCtrl.scala 42:{39,39}]
  wire [4:0] _GEN_125 = 2'h2 == _T_114[1:0] ? w_vn_2 : _GEN_124; // @[FanCtrl.scala 42:{39,39}]
  wire [4:0] _GEN_126 = 2'h3 == _T_114[1:0] ? w_vn_3 : _GEN_125; // @[FanCtrl.scala 42:{39,39}]
  wire [4:0] _GEN_128 = 2'h1 == _T_119[1:0] ? w_vn_1 : w_vn_0; // @[FanCtrl.scala 42:{39,39}]
  wire [4:0] _GEN_129 = 2'h2 == _T_119[1:0] ? w_vn_2 : _GEN_128; // @[FanCtrl.scala 42:{39,39}]
  wire [4:0] _GEN_130 = 2'h3 == _T_119[1:0] ? w_vn_3 : _GEN_129; // @[FanCtrl.scala 42:{39,39}]
  wire  _T_121 = _GEN_126 == _GEN_130; // @[FanCtrl.scala 42:39]
  wire  _T_143 = _GEN_126 != _GEN_130; // @[FanCtrl.scala 50:41]
  wire  _GEN_178 = r_valid_1 & _T_121; // @[FanCtrl.scala 41:34]
  wire [2:0] _T_188 = _T_113 - 3'h1; // @[FanCtrl.scala 88:58]
  wire [4:0] _GEN_206 = 2'h1 == _T_188[1:0] ? w_vn_1 : w_vn_0; // @[FanCtrl.scala 88:{39,39}]
  wire [4:0] _GEN_207 = 2'h2 == _T_188[1:0] ? w_vn_2 : _GEN_206; // @[FanCtrl.scala 88:{39,39}]
  wire [4:0] _GEN_208 = 2'h3 == _T_188[1:0] ? w_vn_3 : _GEN_207; // @[FanCtrl.scala 88:{39,39}]
  wire  _T_200 = _GEN_126 != _GEN_208 & _T_143; // @[FanCtrl.scala 88:67]
  wire  _T_219 = _GEN_126 == _GEN_208 & _T_143; // @[FanCtrl.scala 93:73]
  wire [3:0] _T_228 = 3'h4 * 1'h0; // @[FanCtrl.scala 117:23]
  wire [3:0] _T_230 = _T_228 + 4'h1; // @[FanCtrl.scala 117:29]
  wire [3:0] _T_234 = _T_228 + 4'h2; // @[FanCtrl.scala 117:56]
  wire [4:0] _GEN_254 = 2'h1 == _T_230[1:0] ? w_vn_1 : w_vn_0; // @[FanCtrl.scala 117:{37,37}]
  wire [4:0] _GEN_255 = 2'h2 == _T_230[1:0] ? w_vn_2 : _GEN_254; // @[FanCtrl.scala 117:{37,37}]
  wire [4:0] _GEN_256 = 2'h3 == _T_230[1:0] ? w_vn_3 : _GEN_255; // @[FanCtrl.scala 117:{37,37}]
  wire [4:0] _GEN_258 = 2'h1 == _T_234[1:0] ? w_vn_1 : w_vn_0; // @[FanCtrl.scala 117:{37,37}]
  wire [4:0] _GEN_259 = 2'h2 == _T_234[1:0] ? w_vn_2 : _GEN_258; // @[FanCtrl.scala 117:{37,37}]
  wire [4:0] _GEN_260 = 2'h3 == _T_234[1:0] ? w_vn_3 : _GEN_259; // @[FanCtrl.scala 117:{37,37}]
  wire  _T_236 = _GEN_256 == _GEN_260; // @[FanCtrl.scala 117:37]
  wire [4:0] _T_242 = {{1'd0}, _T_228}; // @[FanCtrl.scala 123:30]
  wire [4:0] _GEN_271 = 2'h1 == _T_242[1:0] ? w_vn_1 : w_vn_0; // @[FanCtrl.scala 123:{38,38}]
  wire [4:0] _GEN_272 = 2'h2 == _T_242[1:0] ? w_vn_2 : _GEN_271; // @[FanCtrl.scala 123:{38,38}]
  wire [4:0] _GEN_273 = 2'h3 == _T_242[1:0] ? w_vn_3 : _GEN_272; // @[FanCtrl.scala 123:{38,38}]
  wire  _T_249 = _GEN_273 == _GEN_256; // @[FanCtrl.scala 123:38]
  wire [3:0] _T_256 = _T_228 + 4'h3; // @[FanCtrl.scala 124:55]
  wire [4:0] _GEN_283 = 2'h1 == _T_256[1:0] ? w_vn_1 : w_vn_0; // @[FanCtrl.scala 124:{36,36}]
  wire [4:0] _GEN_284 = 2'h2 == _T_256[1:0] ? w_vn_2 : _GEN_283; // @[FanCtrl.scala 124:{36,36}]
  wire [4:0] _GEN_285 = 2'h3 == _T_256[1:0] ? w_vn_3 : _GEN_284; // @[FanCtrl.scala 124:{36,36}]
  wire  _T_258 = _GEN_260 == _GEN_285; // @[FanCtrl.scala 124:36]
  wire  _T_259 = _GEN_273 == _GEN_256 & _T_258; // @[FanCtrl.scala 123:65]
  wire [3:0] _T_262 = _T_228 + 4'h4; // @[FanCtrl.scala 125:29]
  wire [4:0] _GEN_287 = 2'h1 == _T_262[1:0] ? w_vn_1 : w_vn_0; // @[FanCtrl.scala 125:{37,37}]
  wire [4:0] _GEN_288 = 2'h2 == _T_262[1:0] ? w_vn_2 : _GEN_287; // @[FanCtrl.scala 125:{37,37}]
  wire [4:0] _GEN_289 = 2'h3 == _T_262[1:0] ? w_vn_3 : _GEN_288; // @[FanCtrl.scala 125:{37,37}]
  wire  _T_268 = _GEN_289 != _GEN_285; // @[FanCtrl.scala 125:37]
  wire  _T_269 = _T_259 & _T_268; // @[FanCtrl.scala 124:64]
  wire  _T_278 = _GEN_256 != _GEN_260; // @[FanCtrl.scala 126:37]
  wire  _T_279 = _T_269 & _T_278; // @[FanCtrl.scala 125:64]
  wire  _T_300 = _T_258 & _T_268; // @[FanCtrl.scala 130:71]
  wire  _T_310 = _T_300 & _T_278; // @[FanCtrl.scala 131:71]
  wire  _T_331 = _T_249 & _T_278; // @[FanCtrl.scala 136:71]
  wire [2:0] _GEN_356 = _T_331 ? 3'h3 : 3'h0; // @[FanCtrl.scala 137:72]
  wire  _GEN_371 = r_valid_1 & _T_236; // @[FanCtrl.scala 116:32]
  assign io_o_reduction_add_0 = r_add_lvl_0Reg_6; // @[FanCtrl.scala 227:{35,35}]
  assign io_o_reduction_add_1 = r_add_lvl_0Reg_7; // @[FanCtrl.scala 227:{35,35}]
  assign io_o_reduction_add_2 = r_add_lvl_1Reg_4; // @[FanCtrl.scala 227:{35,35}]
  assign io_o_reduction_cmd_0 = r_cmd_lvl_0Reg_6; // @[FanCtrl.scala 236:{34,34}]
  assign io_o_reduction_cmd_1 = r_cmd_lvl_0Reg_7; // @[FanCtrl.scala 236:{34,34}]
  assign io_o_reduction_cmd_2 = r_cmd_lvl_1Reg_4; // @[FanCtrl.scala 236:{34,34}]
  assign io_o_reduction_valid = r_valid_3; // @[FanCtrl.scala 226:26]
  always @(posedge clock) begin
    if (reset) begin // @[FanCtrl.scala 19:34]
      r_reduction_add_0 <= 1'h0; // @[FanCtrl.scala 19:34]
    end else begin
      r_reduction_add_0 <= _GEN_54;
    end
    if (reset) begin // @[FanCtrl.scala 19:34]
      r_reduction_add_1 <= 1'h0; // @[FanCtrl.scala 19:34]
    end else begin
      r_reduction_add_1 <= _GEN_178;
    end
    if (reset) begin // @[FanCtrl.scala 19:34]
      r_reduction_add_2 <= 1'h0; // @[FanCtrl.scala 19:34]
    end else begin
      r_reduction_add_2 <= _GEN_371;
    end
    if (reset) begin // @[FanCtrl.scala 20:34]
      r_reduction_cmd_0 <= 3'h0; // @[FanCtrl.scala 20:34]
    end else if (r_valid_1) begin // @[FanCtrl.scala 41:34]
      if (_T_33) begin // @[FanCtrl.scala 51:42]
        r_reduction_cmd_0 <= 3'h5; // @[FanCtrl.scala 53:37]
      end else begin
        r_reduction_cmd_0 <= {{1'd0}, _GEN_49};
      end
    end else begin
      r_reduction_cmd_0 <= 3'h0; // @[FanCtrl.scala 68:33]
    end
    if (reset) begin // @[FanCtrl.scala 20:34]
      r_reduction_cmd_1 <= 3'h0; // @[FanCtrl.scala 20:34]
    end else if (r_valid_1) begin // @[FanCtrl.scala 81:34]
      if (_T_200) begin // @[FanCtrl.scala 89:66]
        r_reduction_cmd_1 <= 3'h5; // @[FanCtrl.scala 91:36]
      end else if (_T_219) begin // @[FanCtrl.scala 94:66]
        r_reduction_cmd_1 <= 3'h4; // @[FanCtrl.scala 96:35]
      end else begin
        r_reduction_cmd_1 <= 3'h0; // @[FanCtrl.scala 99:35]
      end
    end else begin
      r_reduction_cmd_1 <= 3'h0; // @[FanCtrl.scala 103:33]
    end
    if (reset) begin // @[FanCtrl.scala 20:34]
      r_reduction_cmd_2 <= 3'h0; // @[FanCtrl.scala 20:34]
    end else if (r_valid_1) begin // @[FanCtrl.scala 116:32]
      if (_T_279) begin // @[FanCtrl.scala 126:66]
        r_reduction_cmd_2 <= 3'h5;
      end else if (_T_310) begin // @[FanCtrl.scala 132:72]
        r_reduction_cmd_2 <= 3'h4;
      end else begin
        r_reduction_cmd_2 <= _GEN_356;
      end
    end else begin
      r_reduction_cmd_2 <= 3'h0;
    end
    if (reset) begin // @[FanCtrl.scala 23:33]
      r_add_lvl_0Reg_6 <= 1'h0; // @[FanCtrl.scala 23:33]
    end else begin
      r_add_lvl_0Reg_6 <= r_reduction_add_0; // @[FanCtrl.scala 157:20]
    end
    if (reset) begin // @[FanCtrl.scala 23:33]
      r_add_lvl_0Reg_7 <= 1'h0; // @[FanCtrl.scala 23:33]
    end else begin
      r_add_lvl_0Reg_7 <= r_reduction_add_1; // @[FanCtrl.scala 157:20]
    end
    if (reset) begin // @[FanCtrl.scala 24:33]
      r_add_lvl_1Reg_4 <= 1'h0; // @[FanCtrl.scala 24:33]
    end else begin
      r_add_lvl_1Reg_4 <= r_reduction_add_2; // @[FanCtrl.scala 168:20]
    end
    if (reset) begin // @[FanCtrl.scala 27:33]
      r_cmd_lvl_0Reg_6 <= 3'h0; // @[FanCtrl.scala 27:33]
    end else begin
      r_cmd_lvl_0Reg_6 <= r_reduction_cmd_0; // @[FanCtrl.scala 185:20]
    end
    if (reset) begin // @[FanCtrl.scala 27:33]
      r_cmd_lvl_0Reg_7 <= 3'h0; // @[FanCtrl.scala 27:33]
    end else begin
      r_cmd_lvl_0Reg_7 <= r_reduction_cmd_1; // @[FanCtrl.scala 185:20]
    end
    if (reset) begin // @[FanCtrl.scala 28:33]
      r_cmd_lvl_1Reg_4 <= 3'h0; // @[FanCtrl.scala 28:33]
    end else begin
      r_cmd_lvl_1Reg_4 <= r_reduction_cmd_2; // @[FanCtrl.scala 199:20]
    end
    if (reset) begin // @[FanCtrl.scala 34:23]
      w_vn_0 <= 5'h0; // @[FanCtrl.scala 34:23]
    end else begin
      w_vn_0 <= io_i_vn_0; // @[FanCtrl.scala 37:10]
    end
    if (reset) begin // @[FanCtrl.scala 34:23]
      w_vn_1 <= 5'h0; // @[FanCtrl.scala 34:23]
    end else begin
      w_vn_1 <= io_i_vn_1; // @[FanCtrl.scala 37:10]
    end
    if (reset) begin // @[FanCtrl.scala 34:23]
      w_vn_2 <= 5'h0; // @[FanCtrl.scala 34:23]
    end else begin
      w_vn_2 <= io_i_vn_2; // @[FanCtrl.scala 37:10]
    end
    if (reset) begin // @[FanCtrl.scala 34:23]
      w_vn_3 <= 5'h0; // @[FanCtrl.scala 34:23]
    end else begin
      w_vn_3 <= io_i_vn_3; // @[FanCtrl.scala 37:10]
    end
    if (reset) begin // @[FanCtrl.scala 35:26]
      r_valid_0 <= 1'h0; // @[FanCtrl.scala 35:26]
    end else begin
      r_valid_0 <= io_i_data_valid;
    end
    if (reset) begin // @[FanCtrl.scala 35:26]
      r_valid_1 <= 1'h0; // @[FanCtrl.scala 35:26]
    end else begin
      r_valid_1 <= r_valid_0; // @[FanCtrl.scala 222:24]
    end
    if (reset) begin // @[FanCtrl.scala 35:26]
      r_valid_2 <= 1'h0; // @[FanCtrl.scala 35:26]
    end else begin
      r_valid_2 <= r_valid_1; // @[FanCtrl.scala 222:24]
    end
    if (reset) begin // @[FanCtrl.scala 35:26]
      r_valid_3 <= 1'h0; // @[FanCtrl.scala 35:26]
    end else begin
      r_valid_3 <= r_valid_2; // @[FanCtrl.scala 222:24]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_reduction_add_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  r_reduction_add_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  r_reduction_add_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  r_reduction_cmd_0 = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  r_reduction_cmd_1 = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  r_reduction_cmd_2 = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  r_add_lvl_0Reg_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  r_add_lvl_0Reg_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  r_add_lvl_1Reg_4 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  r_cmd_lvl_0Reg_6 = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  r_cmd_lvl_0Reg_7 = _RAND_10[2:0];
  _RAND_11 = {1{`RANDOM}};
  r_cmd_lvl_1Reg_4 = _RAND_11[2:0];
  _RAND_12 = {1{`RANDOM}};
  w_vn_0 = _RAND_12[4:0];
  _RAND_13 = {1{`RANDOM}};
  w_vn_1 = _RAND_13[4:0];
  _RAND_14 = {1{`RANDOM}};
  w_vn_2 = _RAND_14[4:0];
  _RAND_15 = {1{`RANDOM}};
  w_vn_3 = _RAND_15[4:0];
  _RAND_16 = {1{`RANDOM}};
  r_valid_0 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  r_valid_1 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  r_valid_2 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  r_valid_3 = _RAND_19[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Benes3(
  input  [15:0] io_i_data_bus2_0,
  input  [15:0] io_i_data_bus2_1,
  input  [15:0] io_i_data_bus2_2,
  input  [15:0] io_i_data_bus2_3,
  input  [15:0] io_i_data_bus1_0,
  input  [15:0] io_i_data_bus1_1,
  input  [15:0] io_i_data_bus1_2,
  input  [15:0] io_i_data_bus1_3,
  input  [3:0]  io_i_mux_bus_0_0,
  input  [3:0]  io_i_mux_bus_0_1,
  input  [3:0]  io_i_mux_bus_0_2,
  input  [3:0]  io_i_mux_bus_0_3,
  input  [3:0]  io_i_mux_bus_1_0,
  input  [3:0]  io_i_mux_bus_1_1,
  input  [3:0]  io_i_mux_bus_1_2,
  input  [3:0]  io_i_mux_bus_2_0,
  input  [3:0]  io_i_mux_bus_2_1,
  input  [3:0]  io_i_mux_bus_3_0,
  output [15:0] io_o_dist_bus1_0,
  output [15:0] io_o_dist_bus1_1,
  output [15:0] io_o_dist_bus1_2,
  output [15:0] io_o_dist_bus1_3,
  output [15:0] io_o_dist_bus2_0,
  output [15:0] io_o_dist_bus2_1,
  output [15:0] io_o_dist_bus2_2,
  output [15:0] io_o_dist_bus2_3
);
  wire  _T_1 = |io_i_mux_bus_0_0; // @[Benes3.scala 64:35]
  wire  _T_2 = ~(|io_i_mux_bus_0_0); // @[Benes3.scala 64:39]
  wire [1:0] _GEN_4 = 2'h0 % 2'h2; // @[Benes3.scala 25:52]
  wire  parsedindexvalue_first_stage = io_i_mux_bus_0_0[0] & (~_GEN_4[0] | 1'h0 - 1'h1); // @[Benes3.scala 25:26]
  wire  parsedindexvalue_boolArray__0 = io_i_mux_bus_0_0[1]; // @[Benes3.scala 29:92]
  wire  parsedindexvalue_boolArray__1 = io_i_mux_bus_0_0[2]; // @[Benes3.scala 29:92]
  wire [2:0] _GEN_9 = {{2'd0}, parsedindexvalue_first_stage}; // @[Benes3.scala 34:40]
  wire [2:0] _GEN_14 = _GEN_9 % 3'h4; // @[Benes3.scala 34:40]
  wire  parsedindexvalue_calculation = _GEN_14[0]; // @[Benes3.scala 34:40]
  wire  _parsedindexvalue_nextIndex_T = ~parsedindexvalue_calculation; // @[Benes3.scala 36:27]
  wire  _parsedindexvalue_nextIndex_T_1 = ~parsedindexvalue_boolArray__0; // @[Benes3.scala 36:53]
  wire  _parsedindexvalue_nextIndex_T_2 = ~parsedindexvalue_calculation & ~parsedindexvalue_boolArray__0; // @[Benes3.scala 36:36]
  wire  _parsedindexvalue_nextIndex_T_5 = parsedindexvalue_calculation & _parsedindexvalue_nextIndex_T_1; // @[Benes3.scala 37:36]
  wire [1:0] _GEN_440 = {{1'd0}, parsedindexvalue_calculation}; // @[Benes3.scala 38:27]
  wire  _parsedindexvalue_nextIndex_T_6 = _GEN_440 == 2'h2; // @[Benes3.scala 38:27]
  wire  _parsedindexvalue_nextIndex_T_8 = _GEN_440 == 2'h2 & _parsedindexvalue_nextIndex_T_1; // @[Benes3.scala 38:36]
  wire  _parsedindexvalue_nextIndex_T_9 = _GEN_440 == 2'h3; // @[Benes3.scala 39:27]
  wire  _parsedindexvalue_nextIndex_T_11 = _GEN_440 == 2'h3 & _parsedindexvalue_nextIndex_T_1; // @[Benes3.scala 39:36]
  wire  _parsedindexvalue_nextIndex_T_14 = _parsedindexvalue_nextIndex_T & parsedindexvalue_boolArray__0; // @[Benes3.scala 40:36]
  wire [1:0] _GEN_442 = {{1'd0}, parsedindexvalue_first_stage}; // @[Benes3.scala 40:76]
  wire [1:0] _parsedindexvalue_nextIndex_T_16 = _GEN_442 + 2'h2; // @[Benes3.scala 40:76]
  wire  _parsedindexvalue_nextIndex_T_19 = parsedindexvalue_calculation & parsedindexvalue_boolArray__0; // @[Benes3.scala 41:36]
  wire  _parsedindexvalue_nextIndex_T_24 = _parsedindexvalue_nextIndex_T_6 & parsedindexvalue_boolArray__0; // @[Benes3.scala 42:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_26 = _GEN_442 - 2'h2; // @[Benes3.scala 42:76]
  wire  _parsedindexvalue_nextIndex_T_29 = _parsedindexvalue_nextIndex_T_9 & parsedindexvalue_boolArray__0; // @[Benes3.scala 43:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_32 = _parsedindexvalue_nextIndex_T_29 ? _parsedindexvalue_nextIndex_T_26 : {{
    1'd0}, parsedindexvalue_first_stage}; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_33 = _parsedindexvalue_nextIndex_T_24 ? _parsedindexvalue_nextIndex_T_26 :
    _parsedindexvalue_nextIndex_T_32; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_34 = _parsedindexvalue_nextIndex_T_19 ? _parsedindexvalue_nextIndex_T_16 :
    _parsedindexvalue_nextIndex_T_33; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_35 = _parsedindexvalue_nextIndex_T_14 ? _parsedindexvalue_nextIndex_T_16 :
    _parsedindexvalue_nextIndex_T_34; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_36 = _parsedindexvalue_nextIndex_T_11 ? {{1'd0}, parsedindexvalue_first_stage
    } : _parsedindexvalue_nextIndex_T_35; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_37 = _parsedindexvalue_nextIndex_T_8 ? {{1'd0}, parsedindexvalue_first_stage}
     : _parsedindexvalue_nextIndex_T_36; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_38 = _parsedindexvalue_nextIndex_T_5 ? {{1'd0}, parsedindexvalue_first_stage}
     : _parsedindexvalue_nextIndex_T_37; // @[Mux.scala 101:16]
  wire [1:0] parsedindexvalue_nextIndex = _parsedindexvalue_nextIndex_T_2 ? {{1'd0}, parsedindexvalue_first_stage} :
    _parsedindexvalue_nextIndex_T_38; // @[Mux.scala 101:16]
  wire [2:0] _GEN_19 = {{1'd0}, parsedindexvalue_nextIndex}; // @[Benes3.scala 34:40]
  wire [2:0] _GEN_24 = _GEN_19 % 3'h4; // @[Benes3.scala 34:40]
  wire [1:0] parsedindexvalue_calculation_1 = _GEN_24[1:0]; // @[Benes3.scala 34:40]
  wire  _parsedindexvalue_nextIndex_T_39 = parsedindexvalue_calculation_1 == 2'h0; // @[Benes3.scala 36:27]
  wire  _parsedindexvalue_nextIndex_T_40 = ~parsedindexvalue_boolArray__1; // @[Benes3.scala 36:53]
  wire  _parsedindexvalue_nextIndex_T_41 = parsedindexvalue_calculation_1 == 2'h0 & ~parsedindexvalue_boolArray__1; // @[Benes3.scala 36:36]
  wire  _parsedindexvalue_nextIndex_T_42 = parsedindexvalue_calculation_1 == 2'h1; // @[Benes3.scala 37:27]
  wire  _parsedindexvalue_nextIndex_T_44 = parsedindexvalue_calculation_1 == 2'h1 & _parsedindexvalue_nextIndex_T_40; // @[Benes3.scala 37:36]
  wire  _parsedindexvalue_nextIndex_T_45 = parsedindexvalue_calculation_1 == 2'h2; // @[Benes3.scala 38:27]
  wire  _parsedindexvalue_nextIndex_T_47 = parsedindexvalue_calculation_1 == 2'h2 & _parsedindexvalue_nextIndex_T_40; // @[Benes3.scala 38:36]
  wire  _parsedindexvalue_nextIndex_T_48 = parsedindexvalue_calculation_1 == 2'h3; // @[Benes3.scala 39:27]
  wire  _parsedindexvalue_nextIndex_T_50 = parsedindexvalue_calculation_1 == 2'h3 & _parsedindexvalue_nextIndex_T_40; // @[Benes3.scala 39:36]
  wire  _parsedindexvalue_nextIndex_T_53 = _parsedindexvalue_nextIndex_T_39 & parsedindexvalue_boolArray__1; // @[Benes3.scala 40:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_55 = parsedindexvalue_nextIndex + 2'h2; // @[Benes3.scala 40:76]
  wire  _parsedindexvalue_nextIndex_T_58 = _parsedindexvalue_nextIndex_T_42 & parsedindexvalue_boolArray__1; // @[Benes3.scala 41:36]
  wire  _parsedindexvalue_nextIndex_T_63 = _parsedindexvalue_nextIndex_T_45 & parsedindexvalue_boolArray__1; // @[Benes3.scala 42:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_65 = parsedindexvalue_nextIndex - 2'h2; // @[Benes3.scala 42:76]
  wire  _parsedindexvalue_nextIndex_T_68 = _parsedindexvalue_nextIndex_T_48 & parsedindexvalue_boolArray__1; // @[Benes3.scala 43:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_71 = _parsedindexvalue_nextIndex_T_68 ? _parsedindexvalue_nextIndex_T_65 :
    parsedindexvalue_nextIndex; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_72 = _parsedindexvalue_nextIndex_T_63 ? _parsedindexvalue_nextIndex_T_65 :
    _parsedindexvalue_nextIndex_T_71; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_73 = _parsedindexvalue_nextIndex_T_58 ? _parsedindexvalue_nextIndex_T_55 :
    _parsedindexvalue_nextIndex_T_72; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_74 = _parsedindexvalue_nextIndex_T_53 ? _parsedindexvalue_nextIndex_T_55 :
    _parsedindexvalue_nextIndex_T_73; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_75 = _parsedindexvalue_nextIndex_T_50 ? parsedindexvalue_nextIndex :
    _parsedindexvalue_nextIndex_T_74; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_76 = _parsedindexvalue_nextIndex_T_47 ? parsedindexvalue_nextIndex :
    _parsedindexvalue_nextIndex_T_75; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_77 = _parsedindexvalue_nextIndex_T_44 ? parsedindexvalue_nextIndex :
    _parsedindexvalue_nextIndex_T_76; // @[Mux.scala 101:16]
  wire [1:0] parsedindexvalue_nextIndex_1 = _parsedindexvalue_nextIndex_T_41 ? parsedindexvalue_nextIndex :
    _parsedindexvalue_nextIndex_T_77; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_third_stage_T_1 = parsedindexvalue_nextIndex_1 % 2'h2; // @[Benes3.scala 49:61]
  wire [1:0] _parsedindexvalue_third_stage_T_4 = parsedindexvalue_nextIndex_1 + 2'h1; // @[Benes3.scala 49:89]
  wire [1:0] _parsedindexvalue_third_stage_T_6 = parsedindexvalue_nextIndex_1 - 2'h1; // @[Benes3.scala 49:109]
  wire [1:0] _parsedindexvalue_third_stage_T_7 = _parsedindexvalue_third_stage_T_1 == 2'h0 ?
    _parsedindexvalue_third_stage_T_4 : _parsedindexvalue_third_stage_T_6; // @[Benes3.scala 49:47]
  wire [1:0] parsedindexvalue = io_i_mux_bus_0_0[3] ? _parsedindexvalue_third_stage_T_7 : parsedindexvalue_nextIndex_1; // @[Benes3.scala 49:24]
  wire [2:0] _T_3 = {{1'd0}, parsedindexvalue};
  wire [15:0] _GEN_0 = 3'h0 == _T_3 ? io_i_data_bus2_0 : 16'h0; // @[Benes3.scala 67:{47,47}]
  wire [15:0] _GEN_1 = 3'h1 == _T_3 ? io_i_data_bus2_0 : 16'h0; // @[Benes3.scala 67:{47,47}]
  wire [15:0] _GEN_2 = 3'h2 == _T_3 ? io_i_data_bus2_0 : 16'h0; // @[Benes3.scala 67:{47,47}]
  wire [15:0] _GEN_3 = 3'h3 == _T_3 ? io_i_data_bus2_0 : 16'h0; // @[Benes3.scala 67:{47,47}]
  wire [15:0] _GEN_5 = ~(|io_i_mux_bus_0_0) ? _GEN_0 : 16'h0; // @[Benes3.scala 64:49]
  wire [15:0] _GEN_6 = ~(|io_i_mux_bus_0_0) ? _GEN_1 : 16'h0; // @[Benes3.scala 64:49]
  wire [15:0] _GEN_7 = ~(|io_i_mux_bus_0_0) ? _GEN_2 : 16'h0; // @[Benes3.scala 64:49]
  wire [15:0] _GEN_8 = ~(|io_i_mux_bus_0_0) ? _GEN_3 : 16'h0; // @[Benes3.scala 64:49]
  wire [15:0] _GEN_10 = 3'h0 == _T_3 ? io_i_data_bus2_0 : _GEN_5; // @[Benes3.scala 77:{47,47}]
  wire [15:0] _GEN_11 = 3'h1 == _T_3 ? io_i_data_bus2_0 : _GEN_6; // @[Benes3.scala 77:{47,47}]
  wire [15:0] _GEN_12 = 3'h2 == _T_3 ? io_i_data_bus2_0 : _GEN_7; // @[Benes3.scala 77:{47,47}]
  wire [15:0] _GEN_13 = 3'h3 == _T_3 ? io_i_data_bus2_0 : _GEN_8; // @[Benes3.scala 77:{47,47}]
  wire [15:0] _GEN_15 = _T_1 ? _GEN_10 : _GEN_5; // @[Benes3.scala 74:48]
  wire [15:0] _GEN_16 = _T_1 ? _GEN_11 : _GEN_6; // @[Benes3.scala 74:48]
  wire [15:0] _GEN_17 = _T_1 ? _GEN_12 : _GEN_7; // @[Benes3.scala 74:48]
  wire [15:0] _GEN_18 = _T_1 ? _GEN_13 : _GEN_8; // @[Benes3.scala 74:48]
  wire  _T_11 = |io_i_mux_bus_0_1; // @[Benes3.scala 92:71]
  wire  _T_13 = _T_1 & |io_i_mux_bus_0_1; // @[Benes3.scala 92:48]
  wire [15:0] _GEN_20 = 3'h0 == _T_3 ? io_i_data_bus2_0 : _GEN_15; // @[Benes3.scala 95:{48,48}]
  wire [15:0] _GEN_21 = 3'h1 == _T_3 ? io_i_data_bus2_0 : _GEN_16; // @[Benes3.scala 95:{48,48}]
  wire [15:0] _GEN_22 = 3'h2 == _T_3 ? io_i_data_bus2_0 : _GEN_17; // @[Benes3.scala 95:{48,48}]
  wire [15:0] _GEN_23 = 3'h3 == _T_3 ? io_i_data_bus2_0 : _GEN_18; // @[Benes3.scala 95:{48,48}]
  wire  parsedindexvalue2_first_stage = io_i_mux_bus_0_1[0] & (~_GEN_4[0] | 1'h0 - 1'h1); // @[Benes3.scala 25:26]
  wire  parsedindexvalue2_boolArray__0 = io_i_mux_bus_0_1[1]; // @[Benes3.scala 29:92]
  wire  parsedindexvalue2_boolArray__1 = io_i_mux_bus_0_1[2]; // @[Benes3.scala 29:92]
  wire [2:0] _GEN_29 = {{2'd0}, parsedindexvalue2_first_stage}; // @[Benes3.scala 34:40]
  wire [2:0] _GEN_34 = _GEN_29 % 3'h4; // @[Benes3.scala 34:40]
  wire  parsedindexvalue2_calculation = _GEN_34[0]; // @[Benes3.scala 34:40]
  wire  _parsedindexvalue2_nextIndex_T = ~parsedindexvalue2_calculation; // @[Benes3.scala 36:27]
  wire  _parsedindexvalue2_nextIndex_T_1 = ~parsedindexvalue2_boolArray__0; // @[Benes3.scala 36:53]
  wire  _parsedindexvalue2_nextIndex_T_2 = ~parsedindexvalue2_calculation & ~parsedindexvalue2_boolArray__0; // @[Benes3.scala 36:36]
  wire  _parsedindexvalue2_nextIndex_T_5 = parsedindexvalue2_calculation & _parsedindexvalue2_nextIndex_T_1; // @[Benes3.scala 37:36]
  wire [1:0] _GEN_464 = {{1'd0}, parsedindexvalue2_calculation}; // @[Benes3.scala 38:27]
  wire  _parsedindexvalue2_nextIndex_T_6 = _GEN_464 == 2'h2; // @[Benes3.scala 38:27]
  wire  _parsedindexvalue2_nextIndex_T_8 = _GEN_464 == 2'h2 & _parsedindexvalue2_nextIndex_T_1; // @[Benes3.scala 38:36]
  wire  _parsedindexvalue2_nextIndex_T_9 = _GEN_464 == 2'h3; // @[Benes3.scala 39:27]
  wire  _parsedindexvalue2_nextIndex_T_11 = _GEN_464 == 2'h3 & _parsedindexvalue2_nextIndex_T_1; // @[Benes3.scala 39:36]
  wire  _parsedindexvalue2_nextIndex_T_14 = _parsedindexvalue2_nextIndex_T & parsedindexvalue2_boolArray__0; // @[Benes3.scala 40:36]
  wire [1:0] _GEN_466 = {{1'd0}, parsedindexvalue2_first_stage}; // @[Benes3.scala 40:76]
  wire [1:0] _parsedindexvalue2_nextIndex_T_16 = _GEN_466 + 2'h2; // @[Benes3.scala 40:76]
  wire  _parsedindexvalue2_nextIndex_T_19 = parsedindexvalue2_calculation & parsedindexvalue2_boolArray__0; // @[Benes3.scala 41:36]
  wire  _parsedindexvalue2_nextIndex_T_24 = _parsedindexvalue2_nextIndex_T_6 & parsedindexvalue2_boolArray__0; // @[Benes3.scala 42:36]
  wire [1:0] _parsedindexvalue2_nextIndex_T_26 = _GEN_466 - 2'h2; // @[Benes3.scala 42:76]
  wire  _parsedindexvalue2_nextIndex_T_29 = _parsedindexvalue2_nextIndex_T_9 & parsedindexvalue2_boolArray__0; // @[Benes3.scala 43:36]
  wire [1:0] _parsedindexvalue2_nextIndex_T_32 = _parsedindexvalue2_nextIndex_T_29 ? _parsedindexvalue2_nextIndex_T_26
     : {{1'd0}, parsedindexvalue2_first_stage}; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue2_nextIndex_T_33 = _parsedindexvalue2_nextIndex_T_24 ? _parsedindexvalue2_nextIndex_T_26
     : _parsedindexvalue2_nextIndex_T_32; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue2_nextIndex_T_34 = _parsedindexvalue2_nextIndex_T_19 ? _parsedindexvalue2_nextIndex_T_16
     : _parsedindexvalue2_nextIndex_T_33; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue2_nextIndex_T_35 = _parsedindexvalue2_nextIndex_T_14 ? _parsedindexvalue2_nextIndex_T_16
     : _parsedindexvalue2_nextIndex_T_34; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue2_nextIndex_T_36 = _parsedindexvalue2_nextIndex_T_11 ? {{1'd0},
    parsedindexvalue2_first_stage} : _parsedindexvalue2_nextIndex_T_35; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue2_nextIndex_T_37 = _parsedindexvalue2_nextIndex_T_8 ? {{1'd0},
    parsedindexvalue2_first_stage} : _parsedindexvalue2_nextIndex_T_36; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue2_nextIndex_T_38 = _parsedindexvalue2_nextIndex_T_5 ? {{1'd0},
    parsedindexvalue2_first_stage} : _parsedindexvalue2_nextIndex_T_37; // @[Mux.scala 101:16]
  wire [1:0] parsedindexvalue2_nextIndex = _parsedindexvalue2_nextIndex_T_2 ? {{1'd0}, parsedindexvalue2_first_stage} :
    _parsedindexvalue2_nextIndex_T_38; // @[Mux.scala 101:16]
  wire [2:0] _GEN_39 = {{1'd0}, parsedindexvalue2_nextIndex}; // @[Benes3.scala 34:40]
  wire [2:0] _GEN_44 = _GEN_39 % 3'h4; // @[Benes3.scala 34:40]
  wire [1:0] parsedindexvalue2_calculation_1 = _GEN_44[1:0]; // @[Benes3.scala 34:40]
  wire  _parsedindexvalue2_nextIndex_T_39 = parsedindexvalue2_calculation_1 == 2'h0; // @[Benes3.scala 36:27]
  wire  _parsedindexvalue2_nextIndex_T_40 = ~parsedindexvalue2_boolArray__1; // @[Benes3.scala 36:53]
  wire  _parsedindexvalue2_nextIndex_T_41 = parsedindexvalue2_calculation_1 == 2'h0 & ~parsedindexvalue2_boolArray__1; // @[Benes3.scala 36:36]
  wire  _parsedindexvalue2_nextIndex_T_42 = parsedindexvalue2_calculation_1 == 2'h1; // @[Benes3.scala 37:27]
  wire  _parsedindexvalue2_nextIndex_T_44 = parsedindexvalue2_calculation_1 == 2'h1 & _parsedindexvalue2_nextIndex_T_40; // @[Benes3.scala 37:36]
  wire  _parsedindexvalue2_nextIndex_T_45 = parsedindexvalue2_calculation_1 == 2'h2; // @[Benes3.scala 38:27]
  wire  _parsedindexvalue2_nextIndex_T_47 = parsedindexvalue2_calculation_1 == 2'h2 & _parsedindexvalue2_nextIndex_T_40; // @[Benes3.scala 38:36]
  wire  _parsedindexvalue2_nextIndex_T_48 = parsedindexvalue2_calculation_1 == 2'h3; // @[Benes3.scala 39:27]
  wire  _parsedindexvalue2_nextIndex_T_50 = parsedindexvalue2_calculation_1 == 2'h3 & _parsedindexvalue2_nextIndex_T_40; // @[Benes3.scala 39:36]
  wire  _parsedindexvalue2_nextIndex_T_53 = _parsedindexvalue2_nextIndex_T_39 & parsedindexvalue2_boolArray__1; // @[Benes3.scala 40:36]
  wire [1:0] _parsedindexvalue2_nextIndex_T_55 = parsedindexvalue2_nextIndex + 2'h2; // @[Benes3.scala 40:76]
  wire  _parsedindexvalue2_nextIndex_T_58 = _parsedindexvalue2_nextIndex_T_42 & parsedindexvalue2_boolArray__1; // @[Benes3.scala 41:36]
  wire  _parsedindexvalue2_nextIndex_T_63 = _parsedindexvalue2_nextIndex_T_45 & parsedindexvalue2_boolArray__1; // @[Benes3.scala 42:36]
  wire [1:0] _parsedindexvalue2_nextIndex_T_65 = parsedindexvalue2_nextIndex - 2'h2; // @[Benes3.scala 42:76]
  wire  _parsedindexvalue2_nextIndex_T_68 = _parsedindexvalue2_nextIndex_T_48 & parsedindexvalue2_boolArray__1; // @[Benes3.scala 43:36]
  wire [1:0] _parsedindexvalue2_nextIndex_T_71 = _parsedindexvalue2_nextIndex_T_68 ? _parsedindexvalue2_nextIndex_T_65
     : parsedindexvalue2_nextIndex; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue2_nextIndex_T_72 = _parsedindexvalue2_nextIndex_T_63 ? _parsedindexvalue2_nextIndex_T_65
     : _parsedindexvalue2_nextIndex_T_71; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue2_nextIndex_T_73 = _parsedindexvalue2_nextIndex_T_58 ? _parsedindexvalue2_nextIndex_T_55
     : _parsedindexvalue2_nextIndex_T_72; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue2_nextIndex_T_74 = _parsedindexvalue2_nextIndex_T_53 ? _parsedindexvalue2_nextIndex_T_55
     : _parsedindexvalue2_nextIndex_T_73; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue2_nextIndex_T_75 = _parsedindexvalue2_nextIndex_T_50 ? parsedindexvalue2_nextIndex :
    _parsedindexvalue2_nextIndex_T_74; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue2_nextIndex_T_76 = _parsedindexvalue2_nextIndex_T_47 ? parsedindexvalue2_nextIndex :
    _parsedindexvalue2_nextIndex_T_75; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue2_nextIndex_T_77 = _parsedindexvalue2_nextIndex_T_44 ? parsedindexvalue2_nextIndex :
    _parsedindexvalue2_nextIndex_T_76; // @[Mux.scala 101:16]
  wire [1:0] parsedindexvalue2_nextIndex_1 = _parsedindexvalue2_nextIndex_T_41 ? parsedindexvalue2_nextIndex :
    _parsedindexvalue2_nextIndex_T_77; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue2_third_stage_T_1 = parsedindexvalue2_nextIndex_1 % 2'h2; // @[Benes3.scala 49:61]
  wire [1:0] _parsedindexvalue2_third_stage_T_4 = parsedindexvalue2_nextIndex_1 + 2'h1; // @[Benes3.scala 49:89]
  wire [1:0] _parsedindexvalue2_third_stage_T_6 = parsedindexvalue2_nextIndex_1 - 2'h1; // @[Benes3.scala 49:109]
  wire [1:0] _parsedindexvalue2_third_stage_T_7 = _parsedindexvalue2_third_stage_T_1 == 2'h0 ?
    _parsedindexvalue2_third_stage_T_4 : _parsedindexvalue2_third_stage_T_6; // @[Benes3.scala 49:47]
  wire [1:0] parsedindexvalue2 = io_i_mux_bus_0_1[3] ? _parsedindexvalue2_third_stage_T_7 :
    parsedindexvalue2_nextIndex_1; // @[Benes3.scala 49:24]
  wire [2:0] _T_16 = {{1'd0}, parsedindexvalue2};
  wire [15:0] _GEN_25 = 3'h0 == _T_16 ? io_i_data_bus2_0 : _GEN_20; // @[Benes3.scala 100:{44,44}]
  wire [15:0] _GEN_26 = 3'h1 == _T_16 ? io_i_data_bus2_0 : _GEN_21; // @[Benes3.scala 100:{44,44}]
  wire [15:0] _GEN_27 = 3'h2 == _T_16 ? io_i_data_bus2_0 : _GEN_22; // @[Benes3.scala 100:{44,44}]
  wire [15:0] _GEN_28 = 3'h3 == _T_16 ? io_i_data_bus2_0 : _GEN_23; // @[Benes3.scala 100:{44,44}]
  wire [15:0] _GEN_30 = _T_1 & |io_i_mux_bus_0_1 ? _GEN_25 : _GEN_15; // @[Benes3.scala 92:84]
  wire [15:0] _GEN_31 = _T_1 & |io_i_mux_bus_0_1 ? _GEN_26 : _GEN_16; // @[Benes3.scala 92:84]
  wire [15:0] _GEN_32 = _T_1 & |io_i_mux_bus_0_1 ? _GEN_27 : _GEN_17; // @[Benes3.scala 92:84]
  wire [15:0] _GEN_33 = _T_1 & |io_i_mux_bus_0_1 ? _GEN_28 : _GEN_18; // @[Benes3.scala 92:84]
  wire  _T_23 = |io_i_mux_bus_0_2; // @[Benes3.scala 114:107]
  wire  _T_25 = _T_13 & |io_i_mux_bus_0_2; // @[Benes3.scala 114:84]
  wire [15:0] _GEN_35 = 3'h0 == _T_3 ? io_i_data_bus2_0 : _GEN_30; // @[Benes3.scala 117:{48,48}]
  wire [15:0] _GEN_36 = 3'h1 == _T_3 ? io_i_data_bus2_0 : _GEN_31; // @[Benes3.scala 117:{48,48}]
  wire [15:0] _GEN_37 = 3'h2 == _T_3 ? io_i_data_bus2_0 : _GEN_32; // @[Benes3.scala 117:{48,48}]
  wire [15:0] _GEN_38 = 3'h3 == _T_3 ? io_i_data_bus2_0 : _GEN_33; // @[Benes3.scala 117:{48,48}]
  wire [15:0] _GEN_40 = 3'h0 == _T_16 ? io_i_data_bus2_0 : _GEN_35; // @[Benes3.scala 122:{44,44}]
  wire [15:0] _GEN_41 = 3'h1 == _T_16 ? io_i_data_bus2_0 : _GEN_36; // @[Benes3.scala 122:{44,44}]
  wire [15:0] _GEN_42 = 3'h2 == _T_16 ? io_i_data_bus2_0 : _GEN_37; // @[Benes3.scala 122:{44,44}]
  wire [15:0] _GEN_43 = 3'h3 == _T_16 ? io_i_data_bus2_0 : _GEN_38; // @[Benes3.scala 122:{44,44}]
  wire  parsedindexvalue3_first_stage = io_i_mux_bus_0_2[0] & (~_GEN_4[0] | 1'h0 - 1'h1); // @[Benes3.scala 25:26]
  wire  parsedindexvalue3_boolArray__0 = io_i_mux_bus_0_2[1]; // @[Benes3.scala 29:92]
  wire  parsedindexvalue3_boolArray__1 = io_i_mux_bus_0_2[2]; // @[Benes3.scala 29:92]
  wire [2:0] _GEN_49 = {{2'd0}, parsedindexvalue3_first_stage}; // @[Benes3.scala 34:40]
  wire [2:0] _GEN_54 = _GEN_49 % 3'h4; // @[Benes3.scala 34:40]
  wire  parsedindexvalue3_calculation = _GEN_54[0]; // @[Benes3.scala 34:40]
  wire  _parsedindexvalue3_nextIndex_T = ~parsedindexvalue3_calculation; // @[Benes3.scala 36:27]
  wire  _parsedindexvalue3_nextIndex_T_1 = ~parsedindexvalue3_boolArray__0; // @[Benes3.scala 36:53]
  wire  _parsedindexvalue3_nextIndex_T_2 = ~parsedindexvalue3_calculation & ~parsedindexvalue3_boolArray__0; // @[Benes3.scala 36:36]
  wire  _parsedindexvalue3_nextIndex_T_5 = parsedindexvalue3_calculation & _parsedindexvalue3_nextIndex_T_1; // @[Benes3.scala 37:36]
  wire [1:0] _GEN_488 = {{1'd0}, parsedindexvalue3_calculation}; // @[Benes3.scala 38:27]
  wire  _parsedindexvalue3_nextIndex_T_6 = _GEN_488 == 2'h2; // @[Benes3.scala 38:27]
  wire  _parsedindexvalue3_nextIndex_T_8 = _GEN_488 == 2'h2 & _parsedindexvalue3_nextIndex_T_1; // @[Benes3.scala 38:36]
  wire  _parsedindexvalue3_nextIndex_T_9 = _GEN_488 == 2'h3; // @[Benes3.scala 39:27]
  wire  _parsedindexvalue3_nextIndex_T_11 = _GEN_488 == 2'h3 & _parsedindexvalue3_nextIndex_T_1; // @[Benes3.scala 39:36]
  wire  _parsedindexvalue3_nextIndex_T_14 = _parsedindexvalue3_nextIndex_T & parsedindexvalue3_boolArray__0; // @[Benes3.scala 40:36]
  wire [1:0] _GEN_490 = {{1'd0}, parsedindexvalue3_first_stage}; // @[Benes3.scala 40:76]
  wire [1:0] _parsedindexvalue3_nextIndex_T_16 = _GEN_490 + 2'h2; // @[Benes3.scala 40:76]
  wire  _parsedindexvalue3_nextIndex_T_19 = parsedindexvalue3_calculation & parsedindexvalue3_boolArray__0; // @[Benes3.scala 41:36]
  wire  _parsedindexvalue3_nextIndex_T_24 = _parsedindexvalue3_nextIndex_T_6 & parsedindexvalue3_boolArray__0; // @[Benes3.scala 42:36]
  wire [1:0] _parsedindexvalue3_nextIndex_T_26 = _GEN_490 - 2'h2; // @[Benes3.scala 42:76]
  wire  _parsedindexvalue3_nextIndex_T_29 = _parsedindexvalue3_nextIndex_T_9 & parsedindexvalue3_boolArray__0; // @[Benes3.scala 43:36]
  wire [1:0] _parsedindexvalue3_nextIndex_T_32 = _parsedindexvalue3_nextIndex_T_29 ? _parsedindexvalue3_nextIndex_T_26
     : {{1'd0}, parsedindexvalue3_first_stage}; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue3_nextIndex_T_33 = _parsedindexvalue3_nextIndex_T_24 ? _parsedindexvalue3_nextIndex_T_26
     : _parsedindexvalue3_nextIndex_T_32; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue3_nextIndex_T_34 = _parsedindexvalue3_nextIndex_T_19 ? _parsedindexvalue3_nextIndex_T_16
     : _parsedindexvalue3_nextIndex_T_33; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue3_nextIndex_T_35 = _parsedindexvalue3_nextIndex_T_14 ? _parsedindexvalue3_nextIndex_T_16
     : _parsedindexvalue3_nextIndex_T_34; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue3_nextIndex_T_36 = _parsedindexvalue3_nextIndex_T_11 ? {{1'd0},
    parsedindexvalue3_first_stage} : _parsedindexvalue3_nextIndex_T_35; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue3_nextIndex_T_37 = _parsedindexvalue3_nextIndex_T_8 ? {{1'd0},
    parsedindexvalue3_first_stage} : _parsedindexvalue3_nextIndex_T_36; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue3_nextIndex_T_38 = _parsedindexvalue3_nextIndex_T_5 ? {{1'd0},
    parsedindexvalue3_first_stage} : _parsedindexvalue3_nextIndex_T_37; // @[Mux.scala 101:16]
  wire [1:0] parsedindexvalue3_nextIndex = _parsedindexvalue3_nextIndex_T_2 ? {{1'd0}, parsedindexvalue3_first_stage} :
    _parsedindexvalue3_nextIndex_T_38; // @[Mux.scala 101:16]
  wire [2:0] _GEN_59 = {{1'd0}, parsedindexvalue3_nextIndex}; // @[Benes3.scala 34:40]
  wire [2:0] _GEN_64 = _GEN_59 % 3'h4; // @[Benes3.scala 34:40]
  wire [1:0] parsedindexvalue3_calculation_1 = _GEN_64[1:0]; // @[Benes3.scala 34:40]
  wire  _parsedindexvalue3_nextIndex_T_39 = parsedindexvalue3_calculation_1 == 2'h0; // @[Benes3.scala 36:27]
  wire  _parsedindexvalue3_nextIndex_T_40 = ~parsedindexvalue3_boolArray__1; // @[Benes3.scala 36:53]
  wire  _parsedindexvalue3_nextIndex_T_41 = parsedindexvalue3_calculation_1 == 2'h0 & ~parsedindexvalue3_boolArray__1; // @[Benes3.scala 36:36]
  wire  _parsedindexvalue3_nextIndex_T_42 = parsedindexvalue3_calculation_1 == 2'h1; // @[Benes3.scala 37:27]
  wire  _parsedindexvalue3_nextIndex_T_44 = parsedindexvalue3_calculation_1 == 2'h1 & _parsedindexvalue3_nextIndex_T_40; // @[Benes3.scala 37:36]
  wire  _parsedindexvalue3_nextIndex_T_45 = parsedindexvalue3_calculation_1 == 2'h2; // @[Benes3.scala 38:27]
  wire  _parsedindexvalue3_nextIndex_T_47 = parsedindexvalue3_calculation_1 == 2'h2 & _parsedindexvalue3_nextIndex_T_40; // @[Benes3.scala 38:36]
  wire  _parsedindexvalue3_nextIndex_T_48 = parsedindexvalue3_calculation_1 == 2'h3; // @[Benes3.scala 39:27]
  wire  _parsedindexvalue3_nextIndex_T_50 = parsedindexvalue3_calculation_1 == 2'h3 & _parsedindexvalue3_nextIndex_T_40; // @[Benes3.scala 39:36]
  wire  _parsedindexvalue3_nextIndex_T_53 = _parsedindexvalue3_nextIndex_T_39 & parsedindexvalue3_boolArray__1; // @[Benes3.scala 40:36]
  wire [1:0] _parsedindexvalue3_nextIndex_T_55 = parsedindexvalue3_nextIndex + 2'h2; // @[Benes3.scala 40:76]
  wire  _parsedindexvalue3_nextIndex_T_58 = _parsedindexvalue3_nextIndex_T_42 & parsedindexvalue3_boolArray__1; // @[Benes3.scala 41:36]
  wire  _parsedindexvalue3_nextIndex_T_63 = _parsedindexvalue3_nextIndex_T_45 & parsedindexvalue3_boolArray__1; // @[Benes3.scala 42:36]
  wire [1:0] _parsedindexvalue3_nextIndex_T_65 = parsedindexvalue3_nextIndex - 2'h2; // @[Benes3.scala 42:76]
  wire  _parsedindexvalue3_nextIndex_T_68 = _parsedindexvalue3_nextIndex_T_48 & parsedindexvalue3_boolArray__1; // @[Benes3.scala 43:36]
  wire [1:0] _parsedindexvalue3_nextIndex_T_71 = _parsedindexvalue3_nextIndex_T_68 ? _parsedindexvalue3_nextIndex_T_65
     : parsedindexvalue3_nextIndex; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue3_nextIndex_T_72 = _parsedindexvalue3_nextIndex_T_63 ? _parsedindexvalue3_nextIndex_T_65
     : _parsedindexvalue3_nextIndex_T_71; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue3_nextIndex_T_73 = _parsedindexvalue3_nextIndex_T_58 ? _parsedindexvalue3_nextIndex_T_55
     : _parsedindexvalue3_nextIndex_T_72; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue3_nextIndex_T_74 = _parsedindexvalue3_nextIndex_T_53 ? _parsedindexvalue3_nextIndex_T_55
     : _parsedindexvalue3_nextIndex_T_73; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue3_nextIndex_T_75 = _parsedindexvalue3_nextIndex_T_50 ? parsedindexvalue3_nextIndex :
    _parsedindexvalue3_nextIndex_T_74; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue3_nextIndex_T_76 = _parsedindexvalue3_nextIndex_T_47 ? parsedindexvalue3_nextIndex :
    _parsedindexvalue3_nextIndex_T_75; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue3_nextIndex_T_77 = _parsedindexvalue3_nextIndex_T_44 ? parsedindexvalue3_nextIndex :
    _parsedindexvalue3_nextIndex_T_76; // @[Mux.scala 101:16]
  wire [1:0] parsedindexvalue3_nextIndex_1 = _parsedindexvalue3_nextIndex_T_41 ? parsedindexvalue3_nextIndex :
    _parsedindexvalue3_nextIndex_T_77; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue3_third_stage_T_1 = parsedindexvalue3_nextIndex_1 % 2'h2; // @[Benes3.scala 49:61]
  wire [1:0] _parsedindexvalue3_third_stage_T_4 = parsedindexvalue3_nextIndex_1 + 2'h1; // @[Benes3.scala 49:89]
  wire [1:0] _parsedindexvalue3_third_stage_T_6 = parsedindexvalue3_nextIndex_1 - 2'h1; // @[Benes3.scala 49:109]
  wire [1:0] _parsedindexvalue3_third_stage_T_7 = _parsedindexvalue3_third_stage_T_1 == 2'h0 ?
    _parsedindexvalue3_third_stage_T_4 : _parsedindexvalue3_third_stage_T_6; // @[Benes3.scala 49:47]
  wire [1:0] parsedindexvalue3 = io_i_mux_bus_0_2[3] ? _parsedindexvalue3_third_stage_T_7 :
    parsedindexvalue3_nextIndex_1; // @[Benes3.scala 49:24]
  wire [2:0] _T_30 = {{1'd0}, parsedindexvalue3};
  wire [15:0] _GEN_45 = 3'h0 == _T_30 ? io_i_data_bus2_0 : _GEN_40; // @[Benes3.scala 126:{44,44}]
  wire [15:0] _GEN_46 = 3'h1 == _T_30 ? io_i_data_bus2_0 : _GEN_41; // @[Benes3.scala 126:{44,44}]
  wire [15:0] _GEN_47 = 3'h2 == _T_30 ? io_i_data_bus2_0 : _GEN_42; // @[Benes3.scala 126:{44,44}]
  wire [15:0] _GEN_48 = 3'h3 == _T_30 ? io_i_data_bus2_0 : _GEN_43; // @[Benes3.scala 126:{44,44}]
  wire [15:0] _GEN_50 = _T_13 & |io_i_mux_bus_0_2 ? _GEN_45 : _GEN_30; // @[Benes3.scala 114:120]
  wire [15:0] _GEN_51 = _T_13 & |io_i_mux_bus_0_2 ? _GEN_46 : _GEN_31; // @[Benes3.scala 114:120]
  wire [15:0] _GEN_52 = _T_13 & |io_i_mux_bus_0_2 ? _GEN_47 : _GEN_32; // @[Benes3.scala 114:120]
  wire [15:0] _GEN_53 = _T_13 & |io_i_mux_bus_0_2 ? _GEN_48 : _GEN_33; // @[Benes3.scala 114:120]
  wire  _T_40 = |io_i_mux_bus_0_3; // @[Benes3.scala 139:143]
  wire [15:0] _GEN_55 = 3'h0 == _T_3 ? io_i_data_bus2_0 : _GEN_50; // @[Benes3.scala 142:{48,48}]
  wire [15:0] _GEN_56 = 3'h1 == _T_3 ? io_i_data_bus2_0 : _GEN_51; // @[Benes3.scala 142:{48,48}]
  wire [15:0] _GEN_57 = 3'h2 == _T_3 ? io_i_data_bus2_0 : _GEN_52; // @[Benes3.scala 142:{48,48}]
  wire [15:0] _GEN_58 = 3'h3 == _T_3 ? io_i_data_bus2_0 : _GEN_53; // @[Benes3.scala 142:{48,48}]
  wire [15:0] _GEN_60 = 3'h0 == _T_16 ? io_i_data_bus2_0 : _GEN_55; // @[Benes3.scala 147:{44,44}]
  wire [15:0] _GEN_61 = 3'h1 == _T_16 ? io_i_data_bus2_0 : _GEN_56; // @[Benes3.scala 147:{44,44}]
  wire [15:0] _GEN_62 = 3'h2 == _T_16 ? io_i_data_bus2_0 : _GEN_57; // @[Benes3.scala 147:{44,44}]
  wire [15:0] _GEN_63 = 3'h3 == _T_16 ? io_i_data_bus2_0 : _GEN_58; // @[Benes3.scala 147:{44,44}]
  wire [15:0] _GEN_65 = 3'h0 == _T_30 ? io_i_data_bus2_0 : _GEN_60; // @[Benes3.scala 151:{44,44}]
  wire [15:0] _GEN_66 = 3'h1 == _T_30 ? io_i_data_bus2_0 : _GEN_61; // @[Benes3.scala 151:{44,44}]
  wire [15:0] _GEN_67 = 3'h2 == _T_30 ? io_i_data_bus2_0 : _GEN_62; // @[Benes3.scala 151:{44,44}]
  wire [15:0] _GEN_68 = 3'h3 == _T_30 ? io_i_data_bus2_0 : _GEN_63; // @[Benes3.scala 151:{44,44}]
  wire  parsedindexvalue4_first_stage = io_i_mux_bus_0_3[0] & (~_GEN_4[0] | 1'h0 - 1'h1); // @[Benes3.scala 25:26]
  wire  parsedindexvalue4_boolArray__0 = io_i_mux_bus_0_3[1]; // @[Benes3.scala 29:92]
  wire  parsedindexvalue4_boolArray__1 = io_i_mux_bus_0_3[2]; // @[Benes3.scala 29:92]
  wire [2:0] _GEN_69 = {{2'd0}, parsedindexvalue4_first_stage}; // @[Benes3.scala 34:40]
  wire [2:0] _GEN_74 = _GEN_69 % 3'h4; // @[Benes3.scala 34:40]
  wire  parsedindexvalue4_calculation = _GEN_74[0]; // @[Benes3.scala 34:40]
  wire  _parsedindexvalue4_nextIndex_T = ~parsedindexvalue4_calculation; // @[Benes3.scala 36:27]
  wire  _parsedindexvalue4_nextIndex_T_1 = ~parsedindexvalue4_boolArray__0; // @[Benes3.scala 36:53]
  wire  _parsedindexvalue4_nextIndex_T_2 = ~parsedindexvalue4_calculation & ~parsedindexvalue4_boolArray__0; // @[Benes3.scala 36:36]
  wire  _parsedindexvalue4_nextIndex_T_5 = parsedindexvalue4_calculation & _parsedindexvalue4_nextIndex_T_1; // @[Benes3.scala 37:36]
  wire [1:0] _GEN_520 = {{1'd0}, parsedindexvalue4_calculation}; // @[Benes3.scala 38:27]
  wire  _parsedindexvalue4_nextIndex_T_6 = _GEN_520 == 2'h2; // @[Benes3.scala 38:27]
  wire  _parsedindexvalue4_nextIndex_T_8 = _GEN_520 == 2'h2 & _parsedindexvalue4_nextIndex_T_1; // @[Benes3.scala 38:36]
  wire  _parsedindexvalue4_nextIndex_T_9 = _GEN_520 == 2'h3; // @[Benes3.scala 39:27]
  wire  _parsedindexvalue4_nextIndex_T_11 = _GEN_520 == 2'h3 & _parsedindexvalue4_nextIndex_T_1; // @[Benes3.scala 39:36]
  wire  _parsedindexvalue4_nextIndex_T_14 = _parsedindexvalue4_nextIndex_T & parsedindexvalue4_boolArray__0; // @[Benes3.scala 40:36]
  wire [1:0] _GEN_522 = {{1'd0}, parsedindexvalue4_first_stage}; // @[Benes3.scala 40:76]
  wire [1:0] _parsedindexvalue4_nextIndex_T_16 = _GEN_522 + 2'h2; // @[Benes3.scala 40:76]
  wire  _parsedindexvalue4_nextIndex_T_19 = parsedindexvalue4_calculation & parsedindexvalue4_boolArray__0; // @[Benes3.scala 41:36]
  wire  _parsedindexvalue4_nextIndex_T_24 = _parsedindexvalue4_nextIndex_T_6 & parsedindexvalue4_boolArray__0; // @[Benes3.scala 42:36]
  wire [1:0] _parsedindexvalue4_nextIndex_T_26 = _GEN_522 - 2'h2; // @[Benes3.scala 42:76]
  wire  _parsedindexvalue4_nextIndex_T_29 = _parsedindexvalue4_nextIndex_T_9 & parsedindexvalue4_boolArray__0; // @[Benes3.scala 43:36]
  wire [1:0] _parsedindexvalue4_nextIndex_T_32 = _parsedindexvalue4_nextIndex_T_29 ? _parsedindexvalue4_nextIndex_T_26
     : {{1'd0}, parsedindexvalue4_first_stage}; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue4_nextIndex_T_33 = _parsedindexvalue4_nextIndex_T_24 ? _parsedindexvalue4_nextIndex_T_26
     : _parsedindexvalue4_nextIndex_T_32; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue4_nextIndex_T_34 = _parsedindexvalue4_nextIndex_T_19 ? _parsedindexvalue4_nextIndex_T_16
     : _parsedindexvalue4_nextIndex_T_33; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue4_nextIndex_T_35 = _parsedindexvalue4_nextIndex_T_14 ? _parsedindexvalue4_nextIndex_T_16
     : _parsedindexvalue4_nextIndex_T_34; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue4_nextIndex_T_36 = _parsedindexvalue4_nextIndex_T_11 ? {{1'd0},
    parsedindexvalue4_first_stage} : _parsedindexvalue4_nextIndex_T_35; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue4_nextIndex_T_37 = _parsedindexvalue4_nextIndex_T_8 ? {{1'd0},
    parsedindexvalue4_first_stage} : _parsedindexvalue4_nextIndex_T_36; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue4_nextIndex_T_38 = _parsedindexvalue4_nextIndex_T_5 ? {{1'd0},
    parsedindexvalue4_first_stage} : _parsedindexvalue4_nextIndex_T_37; // @[Mux.scala 101:16]
  wire [1:0] parsedindexvalue4_nextIndex = _parsedindexvalue4_nextIndex_T_2 ? {{1'd0}, parsedindexvalue4_first_stage} :
    _parsedindexvalue4_nextIndex_T_38; // @[Mux.scala 101:16]
  wire [2:0] _GEN_79 = {{1'd0}, parsedindexvalue4_nextIndex}; // @[Benes3.scala 34:40]
  wire [2:0] _GEN_84 = _GEN_79 % 3'h4; // @[Benes3.scala 34:40]
  wire [1:0] parsedindexvalue4_calculation_1 = _GEN_84[1:0]; // @[Benes3.scala 34:40]
  wire  _parsedindexvalue4_nextIndex_T_39 = parsedindexvalue4_calculation_1 == 2'h0; // @[Benes3.scala 36:27]
  wire  _parsedindexvalue4_nextIndex_T_40 = ~parsedindexvalue4_boolArray__1; // @[Benes3.scala 36:53]
  wire  _parsedindexvalue4_nextIndex_T_41 = parsedindexvalue4_calculation_1 == 2'h0 & ~parsedindexvalue4_boolArray__1; // @[Benes3.scala 36:36]
  wire  _parsedindexvalue4_nextIndex_T_42 = parsedindexvalue4_calculation_1 == 2'h1; // @[Benes3.scala 37:27]
  wire  _parsedindexvalue4_nextIndex_T_44 = parsedindexvalue4_calculation_1 == 2'h1 & _parsedindexvalue4_nextIndex_T_40; // @[Benes3.scala 37:36]
  wire  _parsedindexvalue4_nextIndex_T_45 = parsedindexvalue4_calculation_1 == 2'h2; // @[Benes3.scala 38:27]
  wire  _parsedindexvalue4_nextIndex_T_47 = parsedindexvalue4_calculation_1 == 2'h2 & _parsedindexvalue4_nextIndex_T_40; // @[Benes3.scala 38:36]
  wire  _parsedindexvalue4_nextIndex_T_48 = parsedindexvalue4_calculation_1 == 2'h3; // @[Benes3.scala 39:27]
  wire  _parsedindexvalue4_nextIndex_T_50 = parsedindexvalue4_calculation_1 == 2'h3 & _parsedindexvalue4_nextIndex_T_40; // @[Benes3.scala 39:36]
  wire  _parsedindexvalue4_nextIndex_T_53 = _parsedindexvalue4_nextIndex_T_39 & parsedindexvalue4_boolArray__1; // @[Benes3.scala 40:36]
  wire [1:0] _parsedindexvalue4_nextIndex_T_55 = parsedindexvalue4_nextIndex + 2'h2; // @[Benes3.scala 40:76]
  wire  _parsedindexvalue4_nextIndex_T_58 = _parsedindexvalue4_nextIndex_T_42 & parsedindexvalue4_boolArray__1; // @[Benes3.scala 41:36]
  wire  _parsedindexvalue4_nextIndex_T_63 = _parsedindexvalue4_nextIndex_T_45 & parsedindexvalue4_boolArray__1; // @[Benes3.scala 42:36]
  wire [1:0] _parsedindexvalue4_nextIndex_T_65 = parsedindexvalue4_nextIndex - 2'h2; // @[Benes3.scala 42:76]
  wire  _parsedindexvalue4_nextIndex_T_68 = _parsedindexvalue4_nextIndex_T_48 & parsedindexvalue4_boolArray__1; // @[Benes3.scala 43:36]
  wire [1:0] _parsedindexvalue4_nextIndex_T_71 = _parsedindexvalue4_nextIndex_T_68 ? _parsedindexvalue4_nextIndex_T_65
     : parsedindexvalue4_nextIndex; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue4_nextIndex_T_72 = _parsedindexvalue4_nextIndex_T_63 ? _parsedindexvalue4_nextIndex_T_65
     : _parsedindexvalue4_nextIndex_T_71; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue4_nextIndex_T_73 = _parsedindexvalue4_nextIndex_T_58 ? _parsedindexvalue4_nextIndex_T_55
     : _parsedindexvalue4_nextIndex_T_72; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue4_nextIndex_T_74 = _parsedindexvalue4_nextIndex_T_53 ? _parsedindexvalue4_nextIndex_T_55
     : _parsedindexvalue4_nextIndex_T_73; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue4_nextIndex_T_75 = _parsedindexvalue4_nextIndex_T_50 ? parsedindexvalue4_nextIndex :
    _parsedindexvalue4_nextIndex_T_74; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue4_nextIndex_T_76 = _parsedindexvalue4_nextIndex_T_47 ? parsedindexvalue4_nextIndex :
    _parsedindexvalue4_nextIndex_T_75; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue4_nextIndex_T_77 = _parsedindexvalue4_nextIndex_T_44 ? parsedindexvalue4_nextIndex :
    _parsedindexvalue4_nextIndex_T_76; // @[Mux.scala 101:16]
  wire [1:0] parsedindexvalue4_nextIndex_1 = _parsedindexvalue4_nextIndex_T_41 ? parsedindexvalue4_nextIndex :
    _parsedindexvalue4_nextIndex_T_77; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue4_third_stage_T_1 = parsedindexvalue4_nextIndex_1 % 2'h2; // @[Benes3.scala 49:61]
  wire [1:0] _parsedindexvalue4_third_stage_T_4 = parsedindexvalue4_nextIndex_1 + 2'h1; // @[Benes3.scala 49:89]
  wire [1:0] _parsedindexvalue4_third_stage_T_6 = parsedindexvalue4_nextIndex_1 - 2'h1; // @[Benes3.scala 49:109]
  wire [1:0] _parsedindexvalue4_third_stage_T_7 = _parsedindexvalue4_third_stage_T_1 == 2'h0 ?
    _parsedindexvalue4_third_stage_T_4 : _parsedindexvalue4_third_stage_T_6; // @[Benes3.scala 49:47]
  wire [1:0] parsedindexvalue4 = io_i_mux_bus_0_3[3] ? _parsedindexvalue4_third_stage_T_7 :
    parsedindexvalue4_nextIndex_1; // @[Benes3.scala 49:24]
  wire [2:0] _T_49 = {{1'd0}, parsedindexvalue4};
  wire [15:0] _GEN_70 = 3'h0 == _T_49 ? io_i_data_bus2_0 : _GEN_65; // @[Benes3.scala 155:{44,44}]
  wire [15:0] _GEN_71 = 3'h1 == _T_49 ? io_i_data_bus2_0 : _GEN_66; // @[Benes3.scala 155:{44,44}]
  wire [15:0] _GEN_72 = 3'h2 == _T_49 ? io_i_data_bus2_0 : _GEN_67; // @[Benes3.scala 155:{44,44}]
  wire [15:0] _GEN_73 = 3'h3 == _T_49 ? io_i_data_bus2_0 : _GEN_68; // @[Benes3.scala 155:{44,44}]
  wire [15:0] _GEN_75 = _T_25 & |io_i_mux_bus_0_3 ? _GEN_70 : _GEN_50; // @[Benes3.scala 139:156]
  wire [15:0] _GEN_76 = _T_25 & |io_i_mux_bus_0_3 ? _GEN_71 : _GEN_51; // @[Benes3.scala 139:156]
  wire [15:0] _GEN_77 = _T_25 & |io_i_mux_bus_0_3 ? _GEN_72 : _GEN_52; // @[Benes3.scala 139:156]
  wire [15:0] _GEN_78 = _T_25 & |io_i_mux_bus_0_3 ? _GEN_73 : _GEN_53; // @[Benes3.scala 139:156]
  wire [15:0] _GEN_80 = 3'h0 == _T_3 ? io_i_data_bus2_0 : _GEN_75; // @[Benes3.scala 164:{48,48}]
  wire [15:0] _GEN_81 = 3'h1 == _T_3 ? io_i_data_bus2_0 : _GEN_76; // @[Benes3.scala 164:{48,48}]
  wire [15:0] _GEN_82 = 3'h2 == _T_3 ? io_i_data_bus2_0 : _GEN_77; // @[Benes3.scala 164:{48,48}]
  wire [15:0] _GEN_83 = 3'h3 == _T_3 ? io_i_data_bus2_0 : _GEN_78; // @[Benes3.scala 164:{48,48}]
  wire [15:0] _GEN_85 = 3'h0 == _T_16 ? io_i_data_bus2_0 : _GEN_80; // @[Benes3.scala 169:{44,44}]
  wire [15:0] _GEN_86 = 3'h1 == _T_16 ? io_i_data_bus2_0 : _GEN_81; // @[Benes3.scala 169:{44,44}]
  wire [15:0] _GEN_87 = 3'h2 == _T_16 ? io_i_data_bus2_0 : _GEN_82; // @[Benes3.scala 169:{44,44}]
  wire [15:0] _GEN_88 = 3'h3 == _T_16 ? io_i_data_bus2_0 : _GEN_83; // @[Benes3.scala 169:{44,44}]
  wire [15:0] _GEN_90 = 3'h0 == _T_30 ? io_i_data_bus2_0 : _GEN_85; // @[Benes3.scala 173:{44,44}]
  wire [15:0] _GEN_91 = 3'h1 == _T_30 ? io_i_data_bus2_0 : _GEN_86; // @[Benes3.scala 173:{44,44}]
  wire [15:0] _GEN_92 = 3'h2 == _T_30 ? io_i_data_bus2_0 : _GEN_87; // @[Benes3.scala 173:{44,44}]
  wire [15:0] _GEN_93 = 3'h3 == _T_30 ? io_i_data_bus2_0 : _GEN_88; // @[Benes3.scala 173:{44,44}]
  wire [15:0] _GEN_95 = 3'h0 == _T_49 ? io_i_data_bus2_0 : _GEN_90; // @[Benes3.scala 177:{44,44}]
  wire [15:0] _GEN_96 = 3'h1 == _T_49 ? io_i_data_bus2_0 : _GEN_91; // @[Benes3.scala 177:{44,44}]
  wire [15:0] _GEN_97 = 3'h2 == _T_49 ? io_i_data_bus2_0 : _GEN_92; // @[Benes3.scala 177:{44,44}]
  wire [15:0] _GEN_98 = 3'h3 == _T_49 ? io_i_data_bus2_0 : _GEN_93; // @[Benes3.scala 177:{44,44}]
  wire [15:0] _GEN_100 = _T_2 & _T_11 & _T_23 & _T_40 ? _GEN_95 : _GEN_75; // @[Benes3.scala 161:160]
  wire [15:0] _GEN_101 = _T_2 & _T_11 & _T_23 & _T_40 ? _GEN_96 : _GEN_76; // @[Benes3.scala 161:160]
  wire [15:0] _GEN_102 = _T_2 & _T_11 & _T_23 & _T_40 ? _GEN_97 : _GEN_77; // @[Benes3.scala 161:160]
  wire [15:0] _GEN_103 = _T_2 & _T_11 & _T_23 & _T_40 ? _GEN_98 : _GEN_78; // @[Benes3.scala 161:160]
  wire [15:0] _GEN_105 = io_i_data_bus2_0 != 16'h0 ? _GEN_100 : 16'h0; // @[Benes3.scala 62:39]
  wire [15:0] _GEN_106 = io_i_data_bus2_0 != 16'h0 ? _GEN_101 : 16'h0; // @[Benes3.scala 62:39]
  wire [15:0] _GEN_107 = io_i_data_bus2_0 != 16'h0 ? _GEN_102 : 16'h0; // @[Benes3.scala 62:39]
  wire [15:0] _GEN_108 = io_i_data_bus2_0 != 16'h0 ? _GEN_103 : 16'h0; // @[Benes3.scala 62:39]
  wire  _T_71 = |io_i_mux_bus_1_0; // @[Benes3.scala 64:35]
  wire  parsedindexvalue_first_stage_2 = io_i_mux_bus_1_0[0] ? 1'h0 : 1'h1; // @[Benes3.scala 25:26]
  wire  parsedindexvalue_boolArray_2_0 = io_i_mux_bus_1_0[1]; // @[Benes3.scala 29:92]
  wire  parsedindexvalue_boolArray_2_1 = io_i_mux_bus_1_0[2]; // @[Benes3.scala 29:92]
  wire [2:0] _GEN_89 = {{2'd0}, parsedindexvalue_first_stage_2}; // @[Benes3.scala 34:40]
  wire [2:0] _GEN_94 = _GEN_89 % 3'h4; // @[Benes3.scala 34:40]
  wire  parsedindexvalue_calculation_4 = _GEN_94[0]; // @[Benes3.scala 34:40]
  wire  _parsedindexvalue_nextIndex_T_156 = ~parsedindexvalue_calculation_4; // @[Benes3.scala 36:27]
  wire  _parsedindexvalue_nextIndex_T_157 = ~parsedindexvalue_boolArray_2_0; // @[Benes3.scala 36:53]
  wire  _parsedindexvalue_nextIndex_T_158 = ~parsedindexvalue_calculation_4 & ~parsedindexvalue_boolArray_2_0; // @[Benes3.scala 36:36]
  wire  _parsedindexvalue_nextIndex_T_161 = parsedindexvalue_calculation_4 & _parsedindexvalue_nextIndex_T_157; // @[Benes3.scala 37:36]
  wire [1:0] _GEN_560 = {{1'd0}, parsedindexvalue_calculation_4}; // @[Benes3.scala 38:27]
  wire  _parsedindexvalue_nextIndex_T_162 = _GEN_560 == 2'h2; // @[Benes3.scala 38:27]
  wire  _parsedindexvalue_nextIndex_T_164 = _GEN_560 == 2'h2 & _parsedindexvalue_nextIndex_T_157; // @[Benes3.scala 38:36]
  wire  _parsedindexvalue_nextIndex_T_165 = _GEN_560 == 2'h3; // @[Benes3.scala 39:27]
  wire  _parsedindexvalue_nextIndex_T_167 = _GEN_560 == 2'h3 & _parsedindexvalue_nextIndex_T_157; // @[Benes3.scala 39:36]
  wire  _parsedindexvalue_nextIndex_T_170 = _parsedindexvalue_nextIndex_T_156 & parsedindexvalue_boolArray_2_0; // @[Benes3.scala 40:36]
  wire [1:0] _GEN_562 = {{1'd0}, parsedindexvalue_first_stage_2}; // @[Benes3.scala 40:76]
  wire [1:0] _parsedindexvalue_nextIndex_T_172 = _GEN_562 + 2'h2; // @[Benes3.scala 40:76]
  wire  _parsedindexvalue_nextIndex_T_175 = parsedindexvalue_calculation_4 & parsedindexvalue_boolArray_2_0; // @[Benes3.scala 41:36]
  wire  _parsedindexvalue_nextIndex_T_180 = _parsedindexvalue_nextIndex_T_162 & parsedindexvalue_boolArray_2_0; // @[Benes3.scala 42:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_182 = _GEN_562 - 2'h2; // @[Benes3.scala 42:76]
  wire  _parsedindexvalue_nextIndex_T_185 = _parsedindexvalue_nextIndex_T_165 & parsedindexvalue_boolArray_2_0; // @[Benes3.scala 43:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_188 = _parsedindexvalue_nextIndex_T_185 ? _parsedindexvalue_nextIndex_T_182
     : {{1'd0}, parsedindexvalue_first_stage_2}; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_189 = _parsedindexvalue_nextIndex_T_180 ? _parsedindexvalue_nextIndex_T_182
     : _parsedindexvalue_nextIndex_T_188; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_190 = _parsedindexvalue_nextIndex_T_175 ? _parsedindexvalue_nextIndex_T_172
     : _parsedindexvalue_nextIndex_T_189; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_191 = _parsedindexvalue_nextIndex_T_170 ? _parsedindexvalue_nextIndex_T_172
     : _parsedindexvalue_nextIndex_T_190; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_192 = _parsedindexvalue_nextIndex_T_167 ? {{1'd0},
    parsedindexvalue_first_stage_2} : _parsedindexvalue_nextIndex_T_191; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_193 = _parsedindexvalue_nextIndex_T_164 ? {{1'd0},
    parsedindexvalue_first_stage_2} : _parsedindexvalue_nextIndex_T_192; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_194 = _parsedindexvalue_nextIndex_T_161 ? {{1'd0},
    parsedindexvalue_first_stage_2} : _parsedindexvalue_nextIndex_T_193; // @[Mux.scala 101:16]
  wire [1:0] parsedindexvalue_nextIndex_4 = _parsedindexvalue_nextIndex_T_158 ? {{1'd0}, parsedindexvalue_first_stage_2}
     : _parsedindexvalue_nextIndex_T_194; // @[Mux.scala 101:16]
  wire [2:0] _GEN_99 = {{1'd0}, parsedindexvalue_nextIndex_4}; // @[Benes3.scala 34:40]
  wire [2:0] _GEN_104 = _GEN_99 % 3'h4; // @[Benes3.scala 34:40]
  wire [1:0] parsedindexvalue_calculation_5 = _GEN_104[1:0]; // @[Benes3.scala 34:40]
  wire  _parsedindexvalue_nextIndex_T_195 = parsedindexvalue_calculation_5 == 2'h0; // @[Benes3.scala 36:27]
  wire  _parsedindexvalue_nextIndex_T_196 = ~parsedindexvalue_boolArray_2_1; // @[Benes3.scala 36:53]
  wire  _parsedindexvalue_nextIndex_T_197 = parsedindexvalue_calculation_5 == 2'h0 & ~parsedindexvalue_boolArray_2_1; // @[Benes3.scala 36:36]
  wire  _parsedindexvalue_nextIndex_T_198 = parsedindexvalue_calculation_5 == 2'h1; // @[Benes3.scala 37:27]
  wire  _parsedindexvalue_nextIndex_T_200 = parsedindexvalue_calculation_5 == 2'h1 & _parsedindexvalue_nextIndex_T_196; // @[Benes3.scala 37:36]
  wire  _parsedindexvalue_nextIndex_T_201 = parsedindexvalue_calculation_5 == 2'h2; // @[Benes3.scala 38:27]
  wire  _parsedindexvalue_nextIndex_T_203 = parsedindexvalue_calculation_5 == 2'h2 & _parsedindexvalue_nextIndex_T_196; // @[Benes3.scala 38:36]
  wire  _parsedindexvalue_nextIndex_T_204 = parsedindexvalue_calculation_5 == 2'h3; // @[Benes3.scala 39:27]
  wire  _parsedindexvalue_nextIndex_T_206 = parsedindexvalue_calculation_5 == 2'h3 & _parsedindexvalue_nextIndex_T_196; // @[Benes3.scala 39:36]
  wire  _parsedindexvalue_nextIndex_T_209 = _parsedindexvalue_nextIndex_T_195 & parsedindexvalue_boolArray_2_1; // @[Benes3.scala 40:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_211 = parsedindexvalue_nextIndex_4 + 2'h2; // @[Benes3.scala 40:76]
  wire  _parsedindexvalue_nextIndex_T_214 = _parsedindexvalue_nextIndex_T_198 & parsedindexvalue_boolArray_2_1; // @[Benes3.scala 41:36]
  wire  _parsedindexvalue_nextIndex_T_219 = _parsedindexvalue_nextIndex_T_201 & parsedindexvalue_boolArray_2_1; // @[Benes3.scala 42:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_221 = parsedindexvalue_nextIndex_4 - 2'h2; // @[Benes3.scala 42:76]
  wire  _parsedindexvalue_nextIndex_T_224 = _parsedindexvalue_nextIndex_T_204 & parsedindexvalue_boolArray_2_1; // @[Benes3.scala 43:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_227 = _parsedindexvalue_nextIndex_T_224 ? _parsedindexvalue_nextIndex_T_221
     : parsedindexvalue_nextIndex_4; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_228 = _parsedindexvalue_nextIndex_T_219 ? _parsedindexvalue_nextIndex_T_221
     : _parsedindexvalue_nextIndex_T_227; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_229 = _parsedindexvalue_nextIndex_T_214 ? _parsedindexvalue_nextIndex_T_211
     : _parsedindexvalue_nextIndex_T_228; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_230 = _parsedindexvalue_nextIndex_T_209 ? _parsedindexvalue_nextIndex_T_211
     : _parsedindexvalue_nextIndex_T_229; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_231 = _parsedindexvalue_nextIndex_T_206 ? parsedindexvalue_nextIndex_4 :
    _parsedindexvalue_nextIndex_T_230; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_232 = _parsedindexvalue_nextIndex_T_203 ? parsedindexvalue_nextIndex_4 :
    _parsedindexvalue_nextIndex_T_231; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_233 = _parsedindexvalue_nextIndex_T_200 ? parsedindexvalue_nextIndex_4 :
    _parsedindexvalue_nextIndex_T_232; // @[Mux.scala 101:16]
  wire [1:0] parsedindexvalue_nextIndex_5 = _parsedindexvalue_nextIndex_T_197 ? parsedindexvalue_nextIndex_4 :
    _parsedindexvalue_nextIndex_T_233; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_third_stage_T_17 = parsedindexvalue_nextIndex_5 % 2'h2; // @[Benes3.scala 49:61]
  wire [1:0] _parsedindexvalue_third_stage_T_20 = parsedindexvalue_nextIndex_5 + 2'h1; // @[Benes3.scala 49:89]
  wire [1:0] _parsedindexvalue_third_stage_T_22 = parsedindexvalue_nextIndex_5 - 2'h1; // @[Benes3.scala 49:109]
  wire [1:0] _parsedindexvalue_third_stage_T_23 = _parsedindexvalue_third_stage_T_17 == 2'h0 ?
    _parsedindexvalue_third_stage_T_20 : _parsedindexvalue_third_stage_T_22; // @[Benes3.scala 49:47]
  wire [1:0] parsedindexvalue_2 = io_i_mux_bus_1_0[3] ? _parsedindexvalue_third_stage_T_23 :
    parsedindexvalue_nextIndex_5; // @[Benes3.scala 49:24]
  wire [2:0] _T_73 = {{1'd0}, parsedindexvalue_2};
  wire [15:0] _GEN_110 = 3'h0 == _T_73 ? io_i_data_bus2_1 : _GEN_105; // @[Benes3.scala 67:{47,47}]
  wire [15:0] _GEN_111 = 3'h1 == _T_73 ? io_i_data_bus2_1 : _GEN_106; // @[Benes3.scala 67:{47,47}]
  wire [15:0] _GEN_112 = 3'h2 == _T_73 ? io_i_data_bus2_1 : _GEN_107; // @[Benes3.scala 67:{47,47}]
  wire [15:0] _GEN_113 = 3'h3 == _T_73 ? io_i_data_bus2_1 : _GEN_108; // @[Benes3.scala 67:{47,47}]
  wire [15:0] _GEN_115 = ~(|io_i_mux_bus_1_0) ? _GEN_110 : _GEN_105; // @[Benes3.scala 64:49]
  wire [15:0] _GEN_116 = ~(|io_i_mux_bus_1_0) ? _GEN_111 : _GEN_106; // @[Benes3.scala 64:49]
  wire [15:0] _GEN_117 = ~(|io_i_mux_bus_1_0) ? _GEN_112 : _GEN_107; // @[Benes3.scala 64:49]
  wire [15:0] _GEN_118 = ~(|io_i_mux_bus_1_0) ? _GEN_113 : _GEN_108; // @[Benes3.scala 64:49]
  wire [15:0] _GEN_120 = 3'h0 == _T_73 ? io_i_data_bus2_1 : _GEN_115; // @[Benes3.scala 77:{47,47}]
  wire [15:0] _GEN_121 = 3'h1 == _T_73 ? io_i_data_bus2_1 : _GEN_116; // @[Benes3.scala 77:{47,47}]
  wire [15:0] _GEN_122 = 3'h2 == _T_73 ? io_i_data_bus2_1 : _GEN_117; // @[Benes3.scala 77:{47,47}]
  wire [15:0] _GEN_123 = 3'h3 == _T_73 ? io_i_data_bus2_1 : _GEN_118; // @[Benes3.scala 77:{47,47}]
  wire [15:0] _GEN_125 = _T_71 ? _GEN_120 : _GEN_115; // @[Benes3.scala 74:48]
  wire [15:0] _GEN_126 = _T_71 ? _GEN_121 : _GEN_116; // @[Benes3.scala 74:48]
  wire [15:0] _GEN_127 = _T_71 ? _GEN_122 : _GEN_117; // @[Benes3.scala 74:48]
  wire [15:0] _GEN_128 = _T_71 ? _GEN_123 : _GEN_118; // @[Benes3.scala 74:48]
  wire  _T_83 = _T_71 & |io_i_mux_bus_1_1; // @[Benes3.scala 92:48]
  wire [15:0] _GEN_130 = 3'h0 == _T_73 ? io_i_data_bus2_1 : _GEN_125; // @[Benes3.scala 95:{48,48}]
  wire [15:0] _GEN_131 = 3'h1 == _T_73 ? io_i_data_bus2_1 : _GEN_126; // @[Benes3.scala 95:{48,48}]
  wire [15:0] _GEN_132 = 3'h2 == _T_73 ? io_i_data_bus2_1 : _GEN_127; // @[Benes3.scala 95:{48,48}]
  wire [15:0] _GEN_133 = 3'h3 == _T_73 ? io_i_data_bus2_1 : _GEN_128; // @[Benes3.scala 95:{48,48}]
  wire  parsedindexvalue2_first_stage_4 = io_i_mux_bus_1_1[0] ? 1'h0 : 1'h1; // @[Benes3.scala 25:26]
  wire  parsedindexvalue2_boolArray_4_0 = io_i_mux_bus_1_1[1]; // @[Benes3.scala 29:92]
  wire  parsedindexvalue2_boolArray_4_1 = io_i_mux_bus_1_1[2]; // @[Benes3.scala 29:92]
  wire [2:0] _GEN_109 = {{2'd0}, parsedindexvalue2_first_stage_4}; // @[Benes3.scala 34:40]
  wire [2:0] _GEN_114 = _GEN_109 % 3'h4; // @[Benes3.scala 34:40]
  wire  parsedindexvalue2_calculation_8 = _GEN_114[0]; // @[Benes3.scala 34:40]
  wire  _parsedindexvalue2_nextIndex_T_312 = ~parsedindexvalue2_calculation_8; // @[Benes3.scala 36:27]
  wire  _parsedindexvalue2_nextIndex_T_313 = ~parsedindexvalue2_boolArray_4_0; // @[Benes3.scala 36:53]
  wire  _parsedindexvalue2_nextIndex_T_314 = ~parsedindexvalue2_calculation_8 & ~parsedindexvalue2_boolArray_4_0; // @[Benes3.scala 36:36]
  wire  _parsedindexvalue2_nextIndex_T_317 = parsedindexvalue2_calculation_8 & _parsedindexvalue2_nextIndex_T_313; // @[Benes3.scala 37:36]
  wire [1:0] _GEN_584 = {{1'd0}, parsedindexvalue2_calculation_8}; // @[Benes3.scala 38:27]
  wire  _parsedindexvalue2_nextIndex_T_318 = _GEN_584 == 2'h2; // @[Benes3.scala 38:27]
  wire  _parsedindexvalue2_nextIndex_T_320 = _GEN_584 == 2'h2 & _parsedindexvalue2_nextIndex_T_313; // @[Benes3.scala 38:36]
  wire  _parsedindexvalue2_nextIndex_T_321 = _GEN_584 == 2'h3; // @[Benes3.scala 39:27]
  wire  _parsedindexvalue2_nextIndex_T_323 = _GEN_584 == 2'h3 & _parsedindexvalue2_nextIndex_T_313; // @[Benes3.scala 39:36]
  wire  _parsedindexvalue2_nextIndex_T_326 = _parsedindexvalue2_nextIndex_T_312 & parsedindexvalue2_boolArray_4_0; // @[Benes3.scala 40:36]
  wire [1:0] _GEN_586 = {{1'd0}, parsedindexvalue2_first_stage_4}; // @[Benes3.scala 40:76]
  wire [1:0] _parsedindexvalue2_nextIndex_T_328 = _GEN_586 + 2'h2; // @[Benes3.scala 40:76]
  wire  _parsedindexvalue2_nextIndex_T_331 = parsedindexvalue2_calculation_8 & parsedindexvalue2_boolArray_4_0; // @[Benes3.scala 41:36]
  wire  _parsedindexvalue2_nextIndex_T_336 = _parsedindexvalue2_nextIndex_T_318 & parsedindexvalue2_boolArray_4_0; // @[Benes3.scala 42:36]
  wire [1:0] _parsedindexvalue2_nextIndex_T_338 = _GEN_586 - 2'h2; // @[Benes3.scala 42:76]
  wire  _parsedindexvalue2_nextIndex_T_341 = _parsedindexvalue2_nextIndex_T_321 & parsedindexvalue2_boolArray_4_0; // @[Benes3.scala 43:36]
  wire [1:0] _parsedindexvalue2_nextIndex_T_344 = _parsedindexvalue2_nextIndex_T_341 ?
    _parsedindexvalue2_nextIndex_T_338 : {{1'd0}, parsedindexvalue2_first_stage_4}; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue2_nextIndex_T_345 = _parsedindexvalue2_nextIndex_T_336 ?
    _parsedindexvalue2_nextIndex_T_338 : _parsedindexvalue2_nextIndex_T_344; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue2_nextIndex_T_346 = _parsedindexvalue2_nextIndex_T_331 ?
    _parsedindexvalue2_nextIndex_T_328 : _parsedindexvalue2_nextIndex_T_345; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue2_nextIndex_T_347 = _parsedindexvalue2_nextIndex_T_326 ?
    _parsedindexvalue2_nextIndex_T_328 : _parsedindexvalue2_nextIndex_T_346; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue2_nextIndex_T_348 = _parsedindexvalue2_nextIndex_T_323 ? {{1'd0},
    parsedindexvalue2_first_stage_4} : _parsedindexvalue2_nextIndex_T_347; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue2_nextIndex_T_349 = _parsedindexvalue2_nextIndex_T_320 ? {{1'd0},
    parsedindexvalue2_first_stage_4} : _parsedindexvalue2_nextIndex_T_348; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue2_nextIndex_T_350 = _parsedindexvalue2_nextIndex_T_317 ? {{1'd0},
    parsedindexvalue2_first_stage_4} : _parsedindexvalue2_nextIndex_T_349; // @[Mux.scala 101:16]
  wire [1:0] parsedindexvalue2_nextIndex_8 = _parsedindexvalue2_nextIndex_T_314 ? {{1'd0},
    parsedindexvalue2_first_stage_4} : _parsedindexvalue2_nextIndex_T_350; // @[Mux.scala 101:16]
  wire [2:0] _GEN_119 = {{1'd0}, parsedindexvalue2_nextIndex_8}; // @[Benes3.scala 34:40]
  wire [2:0] _GEN_124 = _GEN_119 % 3'h4; // @[Benes3.scala 34:40]
  wire [1:0] parsedindexvalue2_calculation_9 = _GEN_124[1:0]; // @[Benes3.scala 34:40]
  wire  _parsedindexvalue2_nextIndex_T_351 = parsedindexvalue2_calculation_9 == 2'h0; // @[Benes3.scala 36:27]
  wire  _parsedindexvalue2_nextIndex_T_352 = ~parsedindexvalue2_boolArray_4_1; // @[Benes3.scala 36:53]
  wire  _parsedindexvalue2_nextIndex_T_353 = parsedindexvalue2_calculation_9 == 2'h0 & ~parsedindexvalue2_boolArray_4_1; // @[Benes3.scala 36:36]
  wire  _parsedindexvalue2_nextIndex_T_354 = parsedindexvalue2_calculation_9 == 2'h1; // @[Benes3.scala 37:27]
  wire  _parsedindexvalue2_nextIndex_T_356 = parsedindexvalue2_calculation_9 == 2'h1 &
    _parsedindexvalue2_nextIndex_T_352; // @[Benes3.scala 37:36]
  wire  _parsedindexvalue2_nextIndex_T_357 = parsedindexvalue2_calculation_9 == 2'h2; // @[Benes3.scala 38:27]
  wire  _parsedindexvalue2_nextIndex_T_359 = parsedindexvalue2_calculation_9 == 2'h2 &
    _parsedindexvalue2_nextIndex_T_352; // @[Benes3.scala 38:36]
  wire  _parsedindexvalue2_nextIndex_T_360 = parsedindexvalue2_calculation_9 == 2'h3; // @[Benes3.scala 39:27]
  wire  _parsedindexvalue2_nextIndex_T_362 = parsedindexvalue2_calculation_9 == 2'h3 &
    _parsedindexvalue2_nextIndex_T_352; // @[Benes3.scala 39:36]
  wire  _parsedindexvalue2_nextIndex_T_365 = _parsedindexvalue2_nextIndex_T_351 & parsedindexvalue2_boolArray_4_1; // @[Benes3.scala 40:36]
  wire [1:0] _parsedindexvalue2_nextIndex_T_367 = parsedindexvalue2_nextIndex_8 + 2'h2; // @[Benes3.scala 40:76]
  wire  _parsedindexvalue2_nextIndex_T_370 = _parsedindexvalue2_nextIndex_T_354 & parsedindexvalue2_boolArray_4_1; // @[Benes3.scala 41:36]
  wire  _parsedindexvalue2_nextIndex_T_375 = _parsedindexvalue2_nextIndex_T_357 & parsedindexvalue2_boolArray_4_1; // @[Benes3.scala 42:36]
  wire [1:0] _parsedindexvalue2_nextIndex_T_377 = parsedindexvalue2_nextIndex_8 - 2'h2; // @[Benes3.scala 42:76]
  wire  _parsedindexvalue2_nextIndex_T_380 = _parsedindexvalue2_nextIndex_T_360 & parsedindexvalue2_boolArray_4_1; // @[Benes3.scala 43:36]
  wire [1:0] _parsedindexvalue2_nextIndex_T_383 = _parsedindexvalue2_nextIndex_T_380 ?
    _parsedindexvalue2_nextIndex_T_377 : parsedindexvalue2_nextIndex_8; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue2_nextIndex_T_384 = _parsedindexvalue2_nextIndex_T_375 ?
    _parsedindexvalue2_nextIndex_T_377 : _parsedindexvalue2_nextIndex_T_383; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue2_nextIndex_T_385 = _parsedindexvalue2_nextIndex_T_370 ?
    _parsedindexvalue2_nextIndex_T_367 : _parsedindexvalue2_nextIndex_T_384; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue2_nextIndex_T_386 = _parsedindexvalue2_nextIndex_T_365 ?
    _parsedindexvalue2_nextIndex_T_367 : _parsedindexvalue2_nextIndex_T_385; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue2_nextIndex_T_387 = _parsedindexvalue2_nextIndex_T_362 ? parsedindexvalue2_nextIndex_8 :
    _parsedindexvalue2_nextIndex_T_386; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue2_nextIndex_T_388 = _parsedindexvalue2_nextIndex_T_359 ? parsedindexvalue2_nextIndex_8 :
    _parsedindexvalue2_nextIndex_T_387; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue2_nextIndex_T_389 = _parsedindexvalue2_nextIndex_T_356 ? parsedindexvalue2_nextIndex_8 :
    _parsedindexvalue2_nextIndex_T_388; // @[Mux.scala 101:16]
  wire [1:0] parsedindexvalue2_nextIndex_9 = _parsedindexvalue2_nextIndex_T_353 ? parsedindexvalue2_nextIndex_8 :
    _parsedindexvalue2_nextIndex_T_389; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue2_third_stage_T_33 = parsedindexvalue2_nextIndex_9 % 2'h2; // @[Benes3.scala 49:61]
  wire [1:0] _parsedindexvalue2_third_stage_T_36 = parsedindexvalue2_nextIndex_9 + 2'h1; // @[Benes3.scala 49:89]
  wire [1:0] _parsedindexvalue2_third_stage_T_38 = parsedindexvalue2_nextIndex_9 - 2'h1; // @[Benes3.scala 49:109]
  wire [1:0] _parsedindexvalue2_third_stage_T_39 = _parsedindexvalue2_third_stage_T_33 == 2'h0 ?
    _parsedindexvalue2_third_stage_T_36 : _parsedindexvalue2_third_stage_T_38; // @[Benes3.scala 49:47]
  wire [1:0] parsedindexvalue2_4 = io_i_mux_bus_1_1[3] ? _parsedindexvalue2_third_stage_T_39 :
    parsedindexvalue2_nextIndex_9; // @[Benes3.scala 49:24]
  wire [2:0] _T_86 = {{1'd0}, parsedindexvalue2_4};
  wire [15:0] _GEN_135 = 3'h0 == _T_86 ? io_i_data_bus2_1 : _GEN_130; // @[Benes3.scala 100:{44,44}]
  wire [15:0] _GEN_136 = 3'h1 == _T_86 ? io_i_data_bus2_1 : _GEN_131; // @[Benes3.scala 100:{44,44}]
  wire [15:0] _GEN_137 = 3'h2 == _T_86 ? io_i_data_bus2_1 : _GEN_132; // @[Benes3.scala 100:{44,44}]
  wire [15:0] _GEN_138 = 3'h3 == _T_86 ? io_i_data_bus2_1 : _GEN_133; // @[Benes3.scala 100:{44,44}]
  wire [15:0] _GEN_140 = _T_71 & |io_i_mux_bus_1_1 ? _GEN_135 : _GEN_125; // @[Benes3.scala 92:84]
  wire [15:0] _GEN_141 = _T_71 & |io_i_mux_bus_1_1 ? _GEN_136 : _GEN_126; // @[Benes3.scala 92:84]
  wire [15:0] _GEN_142 = _T_71 & |io_i_mux_bus_1_1 ? _GEN_137 : _GEN_127; // @[Benes3.scala 92:84]
  wire [15:0] _GEN_143 = _T_71 & |io_i_mux_bus_1_1 ? _GEN_138 : _GEN_128; // @[Benes3.scala 92:84]
  wire [15:0] _GEN_145 = 3'h0 == _T_73 ? io_i_data_bus2_1 : _GEN_140; // @[Benes3.scala 117:{48,48}]
  wire [15:0] _GEN_146 = 3'h1 == _T_73 ? io_i_data_bus2_1 : _GEN_141; // @[Benes3.scala 117:{48,48}]
  wire [15:0] _GEN_147 = 3'h2 == _T_73 ? io_i_data_bus2_1 : _GEN_142; // @[Benes3.scala 117:{48,48}]
  wire [15:0] _GEN_148 = 3'h3 == _T_73 ? io_i_data_bus2_1 : _GEN_143; // @[Benes3.scala 117:{48,48}]
  wire [15:0] _GEN_150 = 3'h0 == _T_86 ? io_i_data_bus2_1 : _GEN_145; // @[Benes3.scala 122:{44,44}]
  wire [15:0] _GEN_151 = 3'h1 == _T_86 ? io_i_data_bus2_1 : _GEN_146; // @[Benes3.scala 122:{44,44}]
  wire [15:0] _GEN_152 = 3'h2 == _T_86 ? io_i_data_bus2_1 : _GEN_147; // @[Benes3.scala 122:{44,44}]
  wire [15:0] _GEN_153 = 3'h3 == _T_86 ? io_i_data_bus2_1 : _GEN_148; // @[Benes3.scala 122:{44,44}]
  wire  parsedindexvalue3_first_stage_3 = io_i_mux_bus_1_2[0] ? 1'h0 : 1'h1; // @[Benes3.scala 25:26]
  wire  parsedindexvalue3_boolArray_3_0 = io_i_mux_bus_1_2[1]; // @[Benes3.scala 29:92]
  wire  parsedindexvalue3_boolArray_3_1 = io_i_mux_bus_1_2[2]; // @[Benes3.scala 29:92]
  wire [2:0] _GEN_129 = {{2'd0}, parsedindexvalue3_first_stage_3}; // @[Benes3.scala 34:40]
  wire [2:0] _GEN_134 = _GEN_129 % 3'h4; // @[Benes3.scala 34:40]
  wire  parsedindexvalue3_calculation_6 = _GEN_134[0]; // @[Benes3.scala 34:40]
  wire  _parsedindexvalue3_nextIndex_T_234 = ~parsedindexvalue3_calculation_6; // @[Benes3.scala 36:27]
  wire  _parsedindexvalue3_nextIndex_T_235 = ~parsedindexvalue3_boolArray_3_0; // @[Benes3.scala 36:53]
  wire  _parsedindexvalue3_nextIndex_T_236 = ~parsedindexvalue3_calculation_6 & ~parsedindexvalue3_boolArray_3_0; // @[Benes3.scala 36:36]
  wire  _parsedindexvalue3_nextIndex_T_239 = parsedindexvalue3_calculation_6 & _parsedindexvalue3_nextIndex_T_235; // @[Benes3.scala 37:36]
  wire [1:0] _GEN_608 = {{1'd0}, parsedindexvalue3_calculation_6}; // @[Benes3.scala 38:27]
  wire  _parsedindexvalue3_nextIndex_T_240 = _GEN_608 == 2'h2; // @[Benes3.scala 38:27]
  wire  _parsedindexvalue3_nextIndex_T_242 = _GEN_608 == 2'h2 & _parsedindexvalue3_nextIndex_T_235; // @[Benes3.scala 38:36]
  wire  _parsedindexvalue3_nextIndex_T_243 = _GEN_608 == 2'h3; // @[Benes3.scala 39:27]
  wire  _parsedindexvalue3_nextIndex_T_245 = _GEN_608 == 2'h3 & _parsedindexvalue3_nextIndex_T_235; // @[Benes3.scala 39:36]
  wire  _parsedindexvalue3_nextIndex_T_248 = _parsedindexvalue3_nextIndex_T_234 & parsedindexvalue3_boolArray_3_0; // @[Benes3.scala 40:36]
  wire [1:0] _GEN_610 = {{1'd0}, parsedindexvalue3_first_stage_3}; // @[Benes3.scala 40:76]
  wire [1:0] _parsedindexvalue3_nextIndex_T_250 = _GEN_610 + 2'h2; // @[Benes3.scala 40:76]
  wire  _parsedindexvalue3_nextIndex_T_253 = parsedindexvalue3_calculation_6 & parsedindexvalue3_boolArray_3_0; // @[Benes3.scala 41:36]
  wire  _parsedindexvalue3_nextIndex_T_258 = _parsedindexvalue3_nextIndex_T_240 & parsedindexvalue3_boolArray_3_0; // @[Benes3.scala 42:36]
  wire [1:0] _parsedindexvalue3_nextIndex_T_260 = _GEN_610 - 2'h2; // @[Benes3.scala 42:76]
  wire  _parsedindexvalue3_nextIndex_T_263 = _parsedindexvalue3_nextIndex_T_243 & parsedindexvalue3_boolArray_3_0; // @[Benes3.scala 43:36]
  wire [1:0] _parsedindexvalue3_nextIndex_T_266 = _parsedindexvalue3_nextIndex_T_263 ?
    _parsedindexvalue3_nextIndex_T_260 : {{1'd0}, parsedindexvalue3_first_stage_3}; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue3_nextIndex_T_267 = _parsedindexvalue3_nextIndex_T_258 ?
    _parsedindexvalue3_nextIndex_T_260 : _parsedindexvalue3_nextIndex_T_266; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue3_nextIndex_T_268 = _parsedindexvalue3_nextIndex_T_253 ?
    _parsedindexvalue3_nextIndex_T_250 : _parsedindexvalue3_nextIndex_T_267; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue3_nextIndex_T_269 = _parsedindexvalue3_nextIndex_T_248 ?
    _parsedindexvalue3_nextIndex_T_250 : _parsedindexvalue3_nextIndex_T_268; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue3_nextIndex_T_270 = _parsedindexvalue3_nextIndex_T_245 ? {{1'd0},
    parsedindexvalue3_first_stage_3} : _parsedindexvalue3_nextIndex_T_269; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue3_nextIndex_T_271 = _parsedindexvalue3_nextIndex_T_242 ? {{1'd0},
    parsedindexvalue3_first_stage_3} : _parsedindexvalue3_nextIndex_T_270; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue3_nextIndex_T_272 = _parsedindexvalue3_nextIndex_T_239 ? {{1'd0},
    parsedindexvalue3_first_stage_3} : _parsedindexvalue3_nextIndex_T_271; // @[Mux.scala 101:16]
  wire [1:0] parsedindexvalue3_nextIndex_6 = _parsedindexvalue3_nextIndex_T_236 ? {{1'd0},
    parsedindexvalue3_first_stage_3} : _parsedindexvalue3_nextIndex_T_272; // @[Mux.scala 101:16]
  wire [2:0] _GEN_139 = {{1'd0}, parsedindexvalue3_nextIndex_6}; // @[Benes3.scala 34:40]
  wire [2:0] _GEN_144 = _GEN_139 % 3'h4; // @[Benes3.scala 34:40]
  wire [1:0] parsedindexvalue3_calculation_7 = _GEN_144[1:0]; // @[Benes3.scala 34:40]
  wire  _parsedindexvalue3_nextIndex_T_273 = parsedindexvalue3_calculation_7 == 2'h0; // @[Benes3.scala 36:27]
  wire  _parsedindexvalue3_nextIndex_T_274 = ~parsedindexvalue3_boolArray_3_1; // @[Benes3.scala 36:53]
  wire  _parsedindexvalue3_nextIndex_T_275 = parsedindexvalue3_calculation_7 == 2'h0 & ~parsedindexvalue3_boolArray_3_1; // @[Benes3.scala 36:36]
  wire  _parsedindexvalue3_nextIndex_T_276 = parsedindexvalue3_calculation_7 == 2'h1; // @[Benes3.scala 37:27]
  wire  _parsedindexvalue3_nextIndex_T_278 = parsedindexvalue3_calculation_7 == 2'h1 &
    _parsedindexvalue3_nextIndex_T_274; // @[Benes3.scala 37:36]
  wire  _parsedindexvalue3_nextIndex_T_279 = parsedindexvalue3_calculation_7 == 2'h2; // @[Benes3.scala 38:27]
  wire  _parsedindexvalue3_nextIndex_T_281 = parsedindexvalue3_calculation_7 == 2'h2 &
    _parsedindexvalue3_nextIndex_T_274; // @[Benes3.scala 38:36]
  wire  _parsedindexvalue3_nextIndex_T_282 = parsedindexvalue3_calculation_7 == 2'h3; // @[Benes3.scala 39:27]
  wire  _parsedindexvalue3_nextIndex_T_284 = parsedindexvalue3_calculation_7 == 2'h3 &
    _parsedindexvalue3_nextIndex_T_274; // @[Benes3.scala 39:36]
  wire  _parsedindexvalue3_nextIndex_T_287 = _parsedindexvalue3_nextIndex_T_273 & parsedindexvalue3_boolArray_3_1; // @[Benes3.scala 40:36]
  wire [1:0] _parsedindexvalue3_nextIndex_T_289 = parsedindexvalue3_nextIndex_6 + 2'h2; // @[Benes3.scala 40:76]
  wire  _parsedindexvalue3_nextIndex_T_292 = _parsedindexvalue3_nextIndex_T_276 & parsedindexvalue3_boolArray_3_1; // @[Benes3.scala 41:36]
  wire  _parsedindexvalue3_nextIndex_T_297 = _parsedindexvalue3_nextIndex_T_279 & parsedindexvalue3_boolArray_3_1; // @[Benes3.scala 42:36]
  wire [1:0] _parsedindexvalue3_nextIndex_T_299 = parsedindexvalue3_nextIndex_6 - 2'h2; // @[Benes3.scala 42:76]
  wire  _parsedindexvalue3_nextIndex_T_302 = _parsedindexvalue3_nextIndex_T_282 & parsedindexvalue3_boolArray_3_1; // @[Benes3.scala 43:36]
  wire [1:0] _parsedindexvalue3_nextIndex_T_305 = _parsedindexvalue3_nextIndex_T_302 ?
    _parsedindexvalue3_nextIndex_T_299 : parsedindexvalue3_nextIndex_6; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue3_nextIndex_T_306 = _parsedindexvalue3_nextIndex_T_297 ?
    _parsedindexvalue3_nextIndex_T_299 : _parsedindexvalue3_nextIndex_T_305; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue3_nextIndex_T_307 = _parsedindexvalue3_nextIndex_T_292 ?
    _parsedindexvalue3_nextIndex_T_289 : _parsedindexvalue3_nextIndex_T_306; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue3_nextIndex_T_308 = _parsedindexvalue3_nextIndex_T_287 ?
    _parsedindexvalue3_nextIndex_T_289 : _parsedindexvalue3_nextIndex_T_307; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue3_nextIndex_T_309 = _parsedindexvalue3_nextIndex_T_284 ? parsedindexvalue3_nextIndex_6 :
    _parsedindexvalue3_nextIndex_T_308; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue3_nextIndex_T_310 = _parsedindexvalue3_nextIndex_T_281 ? parsedindexvalue3_nextIndex_6 :
    _parsedindexvalue3_nextIndex_T_309; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue3_nextIndex_T_311 = _parsedindexvalue3_nextIndex_T_278 ? parsedindexvalue3_nextIndex_6 :
    _parsedindexvalue3_nextIndex_T_310; // @[Mux.scala 101:16]
  wire [1:0] parsedindexvalue3_nextIndex_7 = _parsedindexvalue3_nextIndex_T_275 ? parsedindexvalue3_nextIndex_6 :
    _parsedindexvalue3_nextIndex_T_311; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue3_third_stage_T_25 = parsedindexvalue3_nextIndex_7 % 2'h2; // @[Benes3.scala 49:61]
  wire [1:0] _parsedindexvalue3_third_stage_T_28 = parsedindexvalue3_nextIndex_7 + 2'h1; // @[Benes3.scala 49:89]
  wire [1:0] _parsedindexvalue3_third_stage_T_30 = parsedindexvalue3_nextIndex_7 - 2'h1; // @[Benes3.scala 49:109]
  wire [1:0] _parsedindexvalue3_third_stage_T_31 = _parsedindexvalue3_third_stage_T_25 == 2'h0 ?
    _parsedindexvalue3_third_stage_T_28 : _parsedindexvalue3_third_stage_T_30; // @[Benes3.scala 49:47]
  wire [1:0] parsedindexvalue3_3 = io_i_mux_bus_1_2[3] ? _parsedindexvalue3_third_stage_T_31 :
    parsedindexvalue3_nextIndex_7; // @[Benes3.scala 49:24]
  wire [2:0] _T_100 = {{1'd0}, parsedindexvalue3_3};
  wire [15:0] _GEN_155 = 3'h0 == _T_100 ? io_i_data_bus2_1 : _GEN_150; // @[Benes3.scala 126:{44,44}]
  wire [15:0] _GEN_156 = 3'h1 == _T_100 ? io_i_data_bus2_1 : _GEN_151; // @[Benes3.scala 126:{44,44}]
  wire [15:0] _GEN_157 = 3'h2 == _T_100 ? io_i_data_bus2_1 : _GEN_152; // @[Benes3.scala 126:{44,44}]
  wire [15:0] _GEN_158 = 3'h3 == _T_100 ? io_i_data_bus2_1 : _GEN_153; // @[Benes3.scala 126:{44,44}]
  wire [15:0] _GEN_160 = _T_83 & |io_i_mux_bus_1_2 ? _GEN_155 : _GEN_140; // @[Benes3.scala 114:120]
  wire [15:0] _GEN_161 = _T_83 & |io_i_mux_bus_1_2 ? _GEN_156 : _GEN_141; // @[Benes3.scala 114:120]
  wire [15:0] _GEN_162 = _T_83 & |io_i_mux_bus_1_2 ? _GEN_157 : _GEN_142; // @[Benes3.scala 114:120]
  wire [15:0] _GEN_163 = _T_83 & |io_i_mux_bus_1_2 ? _GEN_158 : _GEN_143; // @[Benes3.scala 114:120]
  wire [15:0] _GEN_215 = io_i_data_bus2_1 != 16'h0 ? _GEN_160 : _GEN_105; // @[Benes3.scala 62:39]
  wire [15:0] _GEN_216 = io_i_data_bus2_1 != 16'h0 ? _GEN_161 : _GEN_106; // @[Benes3.scala 62:39]
  wire [15:0] _GEN_217 = io_i_data_bus2_1 != 16'h0 ? _GEN_162 : _GEN_107; // @[Benes3.scala 62:39]
  wire [15:0] _GEN_218 = io_i_data_bus2_1 != 16'h0 ? _GEN_163 : _GEN_108; // @[Benes3.scala 62:39]
  wire  _T_141 = |io_i_mux_bus_2_0; // @[Benes3.scala 64:35]
  wire [1:0] parsedindexvalue_first_stage_4 = io_i_mux_bus_2_0[0] ? 2'h3 : 2'h2; // @[Benes3.scala 25:26]
  wire  parsedindexvalue_boolArray_4_0 = io_i_mux_bus_2_0[1]; // @[Benes3.scala 29:92]
  wire  parsedindexvalue_boolArray_4_1 = io_i_mux_bus_2_0[2]; // @[Benes3.scala 29:92]
  wire [2:0] _GEN_149 = {{1'd0}, parsedindexvalue_first_stage_4}; // @[Benes3.scala 34:40]
  wire [2:0] _GEN_154 = _GEN_149 % 3'h4; // @[Benes3.scala 34:40]
  wire [1:0] parsedindexvalue_calculation_8 = _GEN_154[1:0]; // @[Benes3.scala 34:40]
  wire  _parsedindexvalue_nextIndex_T_312 = parsedindexvalue_calculation_8 == 2'h0; // @[Benes3.scala 36:27]
  wire  _parsedindexvalue_nextIndex_T_313 = ~parsedindexvalue_boolArray_4_0; // @[Benes3.scala 36:53]
  wire  _parsedindexvalue_nextIndex_T_314 = parsedindexvalue_calculation_8 == 2'h0 & ~parsedindexvalue_boolArray_4_0; // @[Benes3.scala 36:36]
  wire  _parsedindexvalue_nextIndex_T_315 = parsedindexvalue_calculation_8 == 2'h1; // @[Benes3.scala 37:27]
  wire  _parsedindexvalue_nextIndex_T_317 = parsedindexvalue_calculation_8 == 2'h1 & _parsedindexvalue_nextIndex_T_313; // @[Benes3.scala 37:36]
  wire  _parsedindexvalue_nextIndex_T_318 = parsedindexvalue_calculation_8 == 2'h2; // @[Benes3.scala 38:27]
  wire  _parsedindexvalue_nextIndex_T_320 = parsedindexvalue_calculation_8 == 2'h2 & _parsedindexvalue_nextIndex_T_313; // @[Benes3.scala 38:36]
  wire  _parsedindexvalue_nextIndex_T_321 = parsedindexvalue_calculation_8 == 2'h3; // @[Benes3.scala 39:27]
  wire  _parsedindexvalue_nextIndex_T_323 = parsedindexvalue_calculation_8 == 2'h3 & _parsedindexvalue_nextIndex_T_313; // @[Benes3.scala 39:36]
  wire  _parsedindexvalue_nextIndex_T_326 = _parsedindexvalue_nextIndex_T_312 & parsedindexvalue_boolArray_4_0; // @[Benes3.scala 40:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_328 = parsedindexvalue_first_stage_4 + 2'h2; // @[Benes3.scala 40:76]
  wire  _parsedindexvalue_nextIndex_T_331 = _parsedindexvalue_nextIndex_T_315 & parsedindexvalue_boolArray_4_0; // @[Benes3.scala 41:36]
  wire  _parsedindexvalue_nextIndex_T_336 = _parsedindexvalue_nextIndex_T_318 & parsedindexvalue_boolArray_4_0; // @[Benes3.scala 42:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_338 = parsedindexvalue_first_stage_4 - 2'h2; // @[Benes3.scala 42:76]
  wire  _parsedindexvalue_nextIndex_T_341 = _parsedindexvalue_nextIndex_T_321 & parsedindexvalue_boolArray_4_0; // @[Benes3.scala 43:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_344 = _parsedindexvalue_nextIndex_T_341 ? _parsedindexvalue_nextIndex_T_338
     : parsedindexvalue_first_stage_4; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_345 = _parsedindexvalue_nextIndex_T_336 ? _parsedindexvalue_nextIndex_T_338
     : _parsedindexvalue_nextIndex_T_344; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_346 = _parsedindexvalue_nextIndex_T_331 ? _parsedindexvalue_nextIndex_T_328
     : _parsedindexvalue_nextIndex_T_345; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_347 = _parsedindexvalue_nextIndex_T_326 ? _parsedindexvalue_nextIndex_T_328
     : _parsedindexvalue_nextIndex_T_346; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_348 = _parsedindexvalue_nextIndex_T_323 ? parsedindexvalue_first_stage_4 :
    _parsedindexvalue_nextIndex_T_347; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_349 = _parsedindexvalue_nextIndex_T_320 ? parsedindexvalue_first_stage_4 :
    _parsedindexvalue_nextIndex_T_348; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_350 = _parsedindexvalue_nextIndex_T_317 ? parsedindexvalue_first_stage_4 :
    _parsedindexvalue_nextIndex_T_349; // @[Mux.scala 101:16]
  wire [1:0] parsedindexvalue_nextIndex_8 = _parsedindexvalue_nextIndex_T_314 ? parsedindexvalue_first_stage_4 :
    _parsedindexvalue_nextIndex_T_350; // @[Mux.scala 101:16]
  wire [2:0] _GEN_159 = {{1'd0}, parsedindexvalue_nextIndex_8}; // @[Benes3.scala 34:40]
  wire [2:0] _GEN_164 = _GEN_159 % 3'h4; // @[Benes3.scala 34:40]
  wire [1:0] parsedindexvalue_calculation_9 = _GEN_164[1:0]; // @[Benes3.scala 34:40]
  wire  _parsedindexvalue_nextIndex_T_351 = parsedindexvalue_calculation_9 == 2'h0; // @[Benes3.scala 36:27]
  wire  _parsedindexvalue_nextIndex_T_352 = ~parsedindexvalue_boolArray_4_1; // @[Benes3.scala 36:53]
  wire  _parsedindexvalue_nextIndex_T_353 = parsedindexvalue_calculation_9 == 2'h0 & ~parsedindexvalue_boolArray_4_1; // @[Benes3.scala 36:36]
  wire  _parsedindexvalue_nextIndex_T_354 = parsedindexvalue_calculation_9 == 2'h1; // @[Benes3.scala 37:27]
  wire  _parsedindexvalue_nextIndex_T_356 = parsedindexvalue_calculation_9 == 2'h1 & _parsedindexvalue_nextIndex_T_352; // @[Benes3.scala 37:36]
  wire  _parsedindexvalue_nextIndex_T_357 = parsedindexvalue_calculation_9 == 2'h2; // @[Benes3.scala 38:27]
  wire  _parsedindexvalue_nextIndex_T_359 = parsedindexvalue_calculation_9 == 2'h2 & _parsedindexvalue_nextIndex_T_352; // @[Benes3.scala 38:36]
  wire  _parsedindexvalue_nextIndex_T_360 = parsedindexvalue_calculation_9 == 2'h3; // @[Benes3.scala 39:27]
  wire  _parsedindexvalue_nextIndex_T_362 = parsedindexvalue_calculation_9 == 2'h3 & _parsedindexvalue_nextIndex_T_352; // @[Benes3.scala 39:36]
  wire  _parsedindexvalue_nextIndex_T_365 = _parsedindexvalue_nextIndex_T_351 & parsedindexvalue_boolArray_4_1; // @[Benes3.scala 40:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_367 = parsedindexvalue_nextIndex_8 + 2'h2; // @[Benes3.scala 40:76]
  wire  _parsedindexvalue_nextIndex_T_370 = _parsedindexvalue_nextIndex_T_354 & parsedindexvalue_boolArray_4_1; // @[Benes3.scala 41:36]
  wire  _parsedindexvalue_nextIndex_T_375 = _parsedindexvalue_nextIndex_T_357 & parsedindexvalue_boolArray_4_1; // @[Benes3.scala 42:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_377 = parsedindexvalue_nextIndex_8 - 2'h2; // @[Benes3.scala 42:76]
  wire  _parsedindexvalue_nextIndex_T_380 = _parsedindexvalue_nextIndex_T_360 & parsedindexvalue_boolArray_4_1; // @[Benes3.scala 43:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_383 = _parsedindexvalue_nextIndex_T_380 ? _parsedindexvalue_nextIndex_T_377
     : parsedindexvalue_nextIndex_8; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_384 = _parsedindexvalue_nextIndex_T_375 ? _parsedindexvalue_nextIndex_T_377
     : _parsedindexvalue_nextIndex_T_383; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_385 = _parsedindexvalue_nextIndex_T_370 ? _parsedindexvalue_nextIndex_T_367
     : _parsedindexvalue_nextIndex_T_384; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_386 = _parsedindexvalue_nextIndex_T_365 ? _parsedindexvalue_nextIndex_T_367
     : _parsedindexvalue_nextIndex_T_385; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_387 = _parsedindexvalue_nextIndex_T_362 ? parsedindexvalue_nextIndex_8 :
    _parsedindexvalue_nextIndex_T_386; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_388 = _parsedindexvalue_nextIndex_T_359 ? parsedindexvalue_nextIndex_8 :
    _parsedindexvalue_nextIndex_T_387; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_389 = _parsedindexvalue_nextIndex_T_356 ? parsedindexvalue_nextIndex_8 :
    _parsedindexvalue_nextIndex_T_388; // @[Mux.scala 101:16]
  wire [1:0] parsedindexvalue_nextIndex_9 = _parsedindexvalue_nextIndex_T_353 ? parsedindexvalue_nextIndex_8 :
    _parsedindexvalue_nextIndex_T_389; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_third_stage_T_33 = parsedindexvalue_nextIndex_9 % 2'h2; // @[Benes3.scala 49:61]
  wire [1:0] _parsedindexvalue_third_stage_T_36 = parsedindexvalue_nextIndex_9 + 2'h1; // @[Benes3.scala 49:89]
  wire [1:0] _parsedindexvalue_third_stage_T_38 = parsedindexvalue_nextIndex_9 - 2'h1; // @[Benes3.scala 49:109]
  wire [1:0] _parsedindexvalue_third_stage_T_39 = _parsedindexvalue_third_stage_T_33 == 2'h0 ?
    _parsedindexvalue_third_stage_T_36 : _parsedindexvalue_third_stage_T_38; // @[Benes3.scala 49:47]
  wire [1:0] parsedindexvalue_4 = io_i_mux_bus_2_0[3] ? _parsedindexvalue_third_stage_T_39 :
    parsedindexvalue_nextIndex_9; // @[Benes3.scala 49:24]
  wire [2:0] _T_143 = {{1'd0}, parsedindexvalue_4};
  wire [15:0] _GEN_220 = 3'h0 == _T_143 ? io_i_data_bus2_2 : _GEN_215; // @[Benes3.scala 67:{47,47}]
  wire [15:0] _GEN_221 = 3'h1 == _T_143 ? io_i_data_bus2_2 : _GEN_216; // @[Benes3.scala 67:{47,47}]
  wire [15:0] _GEN_222 = 3'h2 == _T_143 ? io_i_data_bus2_2 : _GEN_217; // @[Benes3.scala 67:{47,47}]
  wire [15:0] _GEN_223 = 3'h3 == _T_143 ? io_i_data_bus2_2 : _GEN_218; // @[Benes3.scala 67:{47,47}]
  wire [15:0] _GEN_225 = ~(|io_i_mux_bus_2_0) ? _GEN_220 : _GEN_215; // @[Benes3.scala 64:49]
  wire [15:0] _GEN_226 = ~(|io_i_mux_bus_2_0) ? _GEN_221 : _GEN_216; // @[Benes3.scala 64:49]
  wire [15:0] _GEN_227 = ~(|io_i_mux_bus_2_0) ? _GEN_222 : _GEN_217; // @[Benes3.scala 64:49]
  wire [15:0] _GEN_228 = ~(|io_i_mux_bus_2_0) ? _GEN_223 : _GEN_218; // @[Benes3.scala 64:49]
  wire [15:0] _GEN_230 = 3'h0 == _T_143 ? io_i_data_bus2_2 : _GEN_225; // @[Benes3.scala 77:{47,47}]
  wire [15:0] _GEN_231 = 3'h1 == _T_143 ? io_i_data_bus2_2 : _GEN_226; // @[Benes3.scala 77:{47,47}]
  wire [15:0] _GEN_232 = 3'h2 == _T_143 ? io_i_data_bus2_2 : _GEN_227; // @[Benes3.scala 77:{47,47}]
  wire [15:0] _GEN_233 = 3'h3 == _T_143 ? io_i_data_bus2_2 : _GEN_228; // @[Benes3.scala 77:{47,47}]
  wire [15:0] _GEN_235 = _T_141 ? _GEN_230 : _GEN_225; // @[Benes3.scala 74:48]
  wire [15:0] _GEN_236 = _T_141 ? _GEN_231 : _GEN_226; // @[Benes3.scala 74:48]
  wire [15:0] _GEN_237 = _T_141 ? _GEN_232 : _GEN_227; // @[Benes3.scala 74:48]
  wire [15:0] _GEN_238 = _T_141 ? _GEN_233 : _GEN_228; // @[Benes3.scala 74:48]
  wire [15:0] _GEN_240 = 3'h0 == _T_143 ? io_i_data_bus2_2 : _GEN_235; // @[Benes3.scala 95:{48,48}]
  wire [15:0] _GEN_241 = 3'h1 == _T_143 ? io_i_data_bus2_2 : _GEN_236; // @[Benes3.scala 95:{48,48}]
  wire [15:0] _GEN_242 = 3'h2 == _T_143 ? io_i_data_bus2_2 : _GEN_237; // @[Benes3.scala 95:{48,48}]
  wire [15:0] _GEN_243 = 3'h3 == _T_143 ? io_i_data_bus2_2 : _GEN_238; // @[Benes3.scala 95:{48,48}]
  wire [1:0] parsedindexvalue2_first_stage_8 = io_i_mux_bus_2_1[0] ? 2'h3 : 2'h2; // @[Benes3.scala 25:26]
  wire  parsedindexvalue2_boolArray_8_0 = io_i_mux_bus_2_1[1]; // @[Benes3.scala 29:92]
  wire  parsedindexvalue2_boolArray_8_1 = io_i_mux_bus_2_1[2]; // @[Benes3.scala 29:92]
  wire [2:0] _GEN_165 = {{1'd0}, parsedindexvalue2_first_stage_8}; // @[Benes3.scala 34:40]
  wire [2:0] _GEN_166 = _GEN_165 % 3'h4; // @[Benes3.scala 34:40]
  wire [1:0] parsedindexvalue2_calculation_16 = _GEN_166[1:0]; // @[Benes3.scala 34:40]
  wire  _parsedindexvalue2_nextIndex_T_624 = parsedindexvalue2_calculation_16 == 2'h0; // @[Benes3.scala 36:27]
  wire  _parsedindexvalue2_nextIndex_T_625 = ~parsedindexvalue2_boolArray_8_0; // @[Benes3.scala 36:53]
  wire  _parsedindexvalue2_nextIndex_T_626 = parsedindexvalue2_calculation_16 == 2'h0 & ~parsedindexvalue2_boolArray_8_0
    ; // @[Benes3.scala 36:36]
  wire  _parsedindexvalue2_nextIndex_T_627 = parsedindexvalue2_calculation_16 == 2'h1; // @[Benes3.scala 37:27]
  wire  _parsedindexvalue2_nextIndex_T_629 = parsedindexvalue2_calculation_16 == 2'h1 &
    _parsedindexvalue2_nextIndex_T_625; // @[Benes3.scala 37:36]
  wire  _parsedindexvalue2_nextIndex_T_630 = parsedindexvalue2_calculation_16 == 2'h2; // @[Benes3.scala 38:27]
  wire  _parsedindexvalue2_nextIndex_T_632 = parsedindexvalue2_calculation_16 == 2'h2 &
    _parsedindexvalue2_nextIndex_T_625; // @[Benes3.scala 38:36]
  wire  _parsedindexvalue2_nextIndex_T_633 = parsedindexvalue2_calculation_16 == 2'h3; // @[Benes3.scala 39:27]
  wire  _parsedindexvalue2_nextIndex_T_635 = parsedindexvalue2_calculation_16 == 2'h3 &
    _parsedindexvalue2_nextIndex_T_625; // @[Benes3.scala 39:36]
  wire  _parsedindexvalue2_nextIndex_T_638 = _parsedindexvalue2_nextIndex_T_624 & parsedindexvalue2_boolArray_8_0; // @[Benes3.scala 40:36]
  wire [1:0] _parsedindexvalue2_nextIndex_T_640 = parsedindexvalue2_first_stage_8 + 2'h2; // @[Benes3.scala 40:76]
  wire  _parsedindexvalue2_nextIndex_T_643 = _parsedindexvalue2_nextIndex_T_627 & parsedindexvalue2_boolArray_8_0; // @[Benes3.scala 41:36]
  wire  _parsedindexvalue2_nextIndex_T_648 = _parsedindexvalue2_nextIndex_T_630 & parsedindexvalue2_boolArray_8_0; // @[Benes3.scala 42:36]
  wire [1:0] _parsedindexvalue2_nextIndex_T_650 = parsedindexvalue2_first_stage_8 - 2'h2; // @[Benes3.scala 42:76]
  wire  _parsedindexvalue2_nextIndex_T_653 = _parsedindexvalue2_nextIndex_T_633 & parsedindexvalue2_boolArray_8_0; // @[Benes3.scala 43:36]
  wire [1:0] _parsedindexvalue2_nextIndex_T_656 = _parsedindexvalue2_nextIndex_T_653 ?
    _parsedindexvalue2_nextIndex_T_650 : parsedindexvalue2_first_stage_8; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue2_nextIndex_T_657 = _parsedindexvalue2_nextIndex_T_648 ?
    _parsedindexvalue2_nextIndex_T_650 : _parsedindexvalue2_nextIndex_T_656; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue2_nextIndex_T_658 = _parsedindexvalue2_nextIndex_T_643 ?
    _parsedindexvalue2_nextIndex_T_640 : _parsedindexvalue2_nextIndex_T_657; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue2_nextIndex_T_659 = _parsedindexvalue2_nextIndex_T_638 ?
    _parsedindexvalue2_nextIndex_T_640 : _parsedindexvalue2_nextIndex_T_658; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue2_nextIndex_T_660 = _parsedindexvalue2_nextIndex_T_635 ? parsedindexvalue2_first_stage_8
     : _parsedindexvalue2_nextIndex_T_659; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue2_nextIndex_T_661 = _parsedindexvalue2_nextIndex_T_632 ? parsedindexvalue2_first_stage_8
     : _parsedindexvalue2_nextIndex_T_660; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue2_nextIndex_T_662 = _parsedindexvalue2_nextIndex_T_629 ? parsedindexvalue2_first_stage_8
     : _parsedindexvalue2_nextIndex_T_661; // @[Mux.scala 101:16]
  wire [1:0] parsedindexvalue2_nextIndex_16 = _parsedindexvalue2_nextIndex_T_626 ? parsedindexvalue2_first_stage_8 :
    _parsedindexvalue2_nextIndex_T_662; // @[Mux.scala 101:16]
  wire [2:0] _GEN_167 = {{1'd0}, parsedindexvalue2_nextIndex_16}; // @[Benes3.scala 34:40]
  wire [2:0] _GEN_168 = _GEN_167 % 3'h4; // @[Benes3.scala 34:40]
  wire [1:0] parsedindexvalue2_calculation_17 = _GEN_168[1:0]; // @[Benes3.scala 34:40]
  wire  _parsedindexvalue2_nextIndex_T_663 = parsedindexvalue2_calculation_17 == 2'h0; // @[Benes3.scala 36:27]
  wire  _parsedindexvalue2_nextIndex_T_664 = ~parsedindexvalue2_boolArray_8_1; // @[Benes3.scala 36:53]
  wire  _parsedindexvalue2_nextIndex_T_665 = parsedindexvalue2_calculation_17 == 2'h0 & ~parsedindexvalue2_boolArray_8_1
    ; // @[Benes3.scala 36:36]
  wire  _parsedindexvalue2_nextIndex_T_666 = parsedindexvalue2_calculation_17 == 2'h1; // @[Benes3.scala 37:27]
  wire  _parsedindexvalue2_nextIndex_T_668 = parsedindexvalue2_calculation_17 == 2'h1 &
    _parsedindexvalue2_nextIndex_T_664; // @[Benes3.scala 37:36]
  wire  _parsedindexvalue2_nextIndex_T_669 = parsedindexvalue2_calculation_17 == 2'h2; // @[Benes3.scala 38:27]
  wire  _parsedindexvalue2_nextIndex_T_671 = parsedindexvalue2_calculation_17 == 2'h2 &
    _parsedindexvalue2_nextIndex_T_664; // @[Benes3.scala 38:36]
  wire  _parsedindexvalue2_nextIndex_T_672 = parsedindexvalue2_calculation_17 == 2'h3; // @[Benes3.scala 39:27]
  wire  _parsedindexvalue2_nextIndex_T_674 = parsedindexvalue2_calculation_17 == 2'h3 &
    _parsedindexvalue2_nextIndex_T_664; // @[Benes3.scala 39:36]
  wire  _parsedindexvalue2_nextIndex_T_677 = _parsedindexvalue2_nextIndex_T_663 & parsedindexvalue2_boolArray_8_1; // @[Benes3.scala 40:36]
  wire [1:0] _parsedindexvalue2_nextIndex_T_679 = parsedindexvalue2_nextIndex_16 + 2'h2; // @[Benes3.scala 40:76]
  wire  _parsedindexvalue2_nextIndex_T_682 = _parsedindexvalue2_nextIndex_T_666 & parsedindexvalue2_boolArray_8_1; // @[Benes3.scala 41:36]
  wire  _parsedindexvalue2_nextIndex_T_687 = _parsedindexvalue2_nextIndex_T_669 & parsedindexvalue2_boolArray_8_1; // @[Benes3.scala 42:36]
  wire [1:0] _parsedindexvalue2_nextIndex_T_689 = parsedindexvalue2_nextIndex_16 - 2'h2; // @[Benes3.scala 42:76]
  wire  _parsedindexvalue2_nextIndex_T_692 = _parsedindexvalue2_nextIndex_T_672 & parsedindexvalue2_boolArray_8_1; // @[Benes3.scala 43:36]
  wire [1:0] _parsedindexvalue2_nextIndex_T_695 = _parsedindexvalue2_nextIndex_T_692 ?
    _parsedindexvalue2_nextIndex_T_689 : parsedindexvalue2_nextIndex_16; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue2_nextIndex_T_696 = _parsedindexvalue2_nextIndex_T_687 ?
    _parsedindexvalue2_nextIndex_T_689 : _parsedindexvalue2_nextIndex_T_695; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue2_nextIndex_T_697 = _parsedindexvalue2_nextIndex_T_682 ?
    _parsedindexvalue2_nextIndex_T_679 : _parsedindexvalue2_nextIndex_T_696; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue2_nextIndex_T_698 = _parsedindexvalue2_nextIndex_T_677 ?
    _parsedindexvalue2_nextIndex_T_679 : _parsedindexvalue2_nextIndex_T_697; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue2_nextIndex_T_699 = _parsedindexvalue2_nextIndex_T_674 ? parsedindexvalue2_nextIndex_16 :
    _parsedindexvalue2_nextIndex_T_698; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue2_nextIndex_T_700 = _parsedindexvalue2_nextIndex_T_671 ? parsedindexvalue2_nextIndex_16 :
    _parsedindexvalue2_nextIndex_T_699; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue2_nextIndex_T_701 = _parsedindexvalue2_nextIndex_T_668 ? parsedindexvalue2_nextIndex_16 :
    _parsedindexvalue2_nextIndex_T_700; // @[Mux.scala 101:16]
  wire [1:0] parsedindexvalue2_nextIndex_17 = _parsedindexvalue2_nextIndex_T_665 ? parsedindexvalue2_nextIndex_16 :
    _parsedindexvalue2_nextIndex_T_701; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue2_third_stage_T_65 = parsedindexvalue2_nextIndex_17 % 2'h2; // @[Benes3.scala 49:61]
  wire [1:0] _parsedindexvalue2_third_stage_T_68 = parsedindexvalue2_nextIndex_17 + 2'h1; // @[Benes3.scala 49:89]
  wire [1:0] _parsedindexvalue2_third_stage_T_70 = parsedindexvalue2_nextIndex_17 - 2'h1; // @[Benes3.scala 49:109]
  wire [1:0] _parsedindexvalue2_third_stage_T_71 = _parsedindexvalue2_third_stage_T_65 == 2'h0 ?
    _parsedindexvalue2_third_stage_T_68 : _parsedindexvalue2_third_stage_T_70; // @[Benes3.scala 49:47]
  wire [1:0] parsedindexvalue2_8 = io_i_mux_bus_2_1[3] ? _parsedindexvalue2_third_stage_T_71 :
    parsedindexvalue2_nextIndex_17; // @[Benes3.scala 49:24]
  wire [2:0] _T_156 = {{1'd0}, parsedindexvalue2_8};
  wire [15:0] _GEN_245 = 3'h0 == _T_156 ? io_i_data_bus2_2 : _GEN_240; // @[Benes3.scala 100:{44,44}]
  wire [15:0] _GEN_246 = 3'h1 == _T_156 ? io_i_data_bus2_2 : _GEN_241; // @[Benes3.scala 100:{44,44}]
  wire [15:0] _GEN_247 = 3'h2 == _T_156 ? io_i_data_bus2_2 : _GEN_242; // @[Benes3.scala 100:{44,44}]
  wire [15:0] _GEN_248 = 3'h3 == _T_156 ? io_i_data_bus2_2 : _GEN_243; // @[Benes3.scala 100:{44,44}]
  wire [15:0] _GEN_250 = _T_141 & |io_i_mux_bus_2_1 ? _GEN_245 : _GEN_235; // @[Benes3.scala 92:84]
  wire [15:0] _GEN_251 = _T_141 & |io_i_mux_bus_2_1 ? _GEN_246 : _GEN_236; // @[Benes3.scala 92:84]
  wire [15:0] _GEN_252 = _T_141 & |io_i_mux_bus_2_1 ? _GEN_247 : _GEN_237; // @[Benes3.scala 92:84]
  wire [15:0] _GEN_253 = _T_141 & |io_i_mux_bus_2_1 ? _GEN_248 : _GEN_238; // @[Benes3.scala 92:84]
  wire [15:0] _GEN_325 = io_i_data_bus2_2 != 16'h0 ? _GEN_250 : _GEN_215; // @[Benes3.scala 62:39]
  wire [15:0] _GEN_326 = io_i_data_bus2_2 != 16'h0 ? _GEN_251 : _GEN_216; // @[Benes3.scala 62:39]
  wire [15:0] _GEN_327 = io_i_data_bus2_2 != 16'h0 ? _GEN_252 : _GEN_217; // @[Benes3.scala 62:39]
  wire [15:0] _GEN_328 = io_i_data_bus2_2 != 16'h0 ? _GEN_253 : _GEN_218; // @[Benes3.scala 62:39]
  wire  _T_211 = |io_i_mux_bus_3_0; // @[Benes3.scala 64:35]
  wire [1:0] _parsedindexvalue_first_stage_T_49 = 2'h3 % 2'h2; // @[Benes3.scala 25:52]
  wire [1:0] _parsedindexvalue_first_stage_T_54 = 2'h3 - 2'h1; // @[Benes3.scala 25:96]
  wire [1:0] _parsedindexvalue_first_stage_T_55 = _parsedindexvalue_first_stage_T_49 == 2'h0 ? 2'h0 :
    _parsedindexvalue_first_stage_T_54; // @[Benes3.scala 25:40]
  wire [1:0] parsedindexvalue_first_stage_6 = io_i_mux_bus_3_0[0] ? _parsedindexvalue_first_stage_T_55 : 2'h3; // @[Benes3.scala 25:26]
  wire  parsedindexvalue_boolArray_6_0 = io_i_mux_bus_3_0[1]; // @[Benes3.scala 29:92]
  wire  parsedindexvalue_boolArray_6_1 = io_i_mux_bus_3_0[2]; // @[Benes3.scala 29:92]
  wire [2:0] _GEN_169 = {{1'd0}, parsedindexvalue_first_stage_6}; // @[Benes3.scala 34:40]
  wire [2:0] _GEN_170 = _GEN_169 % 3'h4; // @[Benes3.scala 34:40]
  wire [1:0] parsedindexvalue_calculation_12 = _GEN_170[1:0]; // @[Benes3.scala 34:40]
  wire  _parsedindexvalue_nextIndex_T_468 = parsedindexvalue_calculation_12 == 2'h0; // @[Benes3.scala 36:27]
  wire  _parsedindexvalue_nextIndex_T_469 = ~parsedindexvalue_boolArray_6_0; // @[Benes3.scala 36:53]
  wire  _parsedindexvalue_nextIndex_T_470 = parsedindexvalue_calculation_12 == 2'h0 & ~parsedindexvalue_boolArray_6_0; // @[Benes3.scala 36:36]
  wire  _parsedindexvalue_nextIndex_T_471 = parsedindexvalue_calculation_12 == 2'h1; // @[Benes3.scala 37:27]
  wire  _parsedindexvalue_nextIndex_T_473 = parsedindexvalue_calculation_12 == 2'h1 & _parsedindexvalue_nextIndex_T_469; // @[Benes3.scala 37:36]
  wire  _parsedindexvalue_nextIndex_T_474 = parsedindexvalue_calculation_12 == 2'h2; // @[Benes3.scala 38:27]
  wire  _parsedindexvalue_nextIndex_T_476 = parsedindexvalue_calculation_12 == 2'h2 & _parsedindexvalue_nextIndex_T_469; // @[Benes3.scala 38:36]
  wire  _parsedindexvalue_nextIndex_T_477 = parsedindexvalue_calculation_12 == 2'h3; // @[Benes3.scala 39:27]
  wire  _parsedindexvalue_nextIndex_T_479 = parsedindexvalue_calculation_12 == 2'h3 & _parsedindexvalue_nextIndex_T_469; // @[Benes3.scala 39:36]
  wire  _parsedindexvalue_nextIndex_T_482 = _parsedindexvalue_nextIndex_T_468 & parsedindexvalue_boolArray_6_0; // @[Benes3.scala 40:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_484 = parsedindexvalue_first_stage_6 + 2'h2; // @[Benes3.scala 40:76]
  wire  _parsedindexvalue_nextIndex_T_487 = _parsedindexvalue_nextIndex_T_471 & parsedindexvalue_boolArray_6_0; // @[Benes3.scala 41:36]
  wire  _parsedindexvalue_nextIndex_T_492 = _parsedindexvalue_nextIndex_T_474 & parsedindexvalue_boolArray_6_0; // @[Benes3.scala 42:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_494 = parsedindexvalue_first_stage_6 - 2'h2; // @[Benes3.scala 42:76]
  wire  _parsedindexvalue_nextIndex_T_497 = _parsedindexvalue_nextIndex_T_477 & parsedindexvalue_boolArray_6_0; // @[Benes3.scala 43:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_500 = _parsedindexvalue_nextIndex_T_497 ? _parsedindexvalue_nextIndex_T_494
     : parsedindexvalue_first_stage_6; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_501 = _parsedindexvalue_nextIndex_T_492 ? _parsedindexvalue_nextIndex_T_494
     : _parsedindexvalue_nextIndex_T_500; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_502 = _parsedindexvalue_nextIndex_T_487 ? _parsedindexvalue_nextIndex_T_484
     : _parsedindexvalue_nextIndex_T_501; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_503 = _parsedindexvalue_nextIndex_T_482 ? _parsedindexvalue_nextIndex_T_484
     : _parsedindexvalue_nextIndex_T_502; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_504 = _parsedindexvalue_nextIndex_T_479 ? parsedindexvalue_first_stage_6 :
    _parsedindexvalue_nextIndex_T_503; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_505 = _parsedindexvalue_nextIndex_T_476 ? parsedindexvalue_first_stage_6 :
    _parsedindexvalue_nextIndex_T_504; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_506 = _parsedindexvalue_nextIndex_T_473 ? parsedindexvalue_first_stage_6 :
    _parsedindexvalue_nextIndex_T_505; // @[Mux.scala 101:16]
  wire [1:0] parsedindexvalue_nextIndex_12 = _parsedindexvalue_nextIndex_T_470 ? parsedindexvalue_first_stage_6 :
    _parsedindexvalue_nextIndex_T_506; // @[Mux.scala 101:16]
  wire [2:0] _GEN_171 = {{1'd0}, parsedindexvalue_nextIndex_12}; // @[Benes3.scala 34:40]
  wire [2:0] _GEN_172 = _GEN_171 % 3'h4; // @[Benes3.scala 34:40]
  wire [1:0] parsedindexvalue_calculation_13 = _GEN_172[1:0]; // @[Benes3.scala 34:40]
  wire  _parsedindexvalue_nextIndex_T_507 = parsedindexvalue_calculation_13 == 2'h0; // @[Benes3.scala 36:27]
  wire  _parsedindexvalue_nextIndex_T_508 = ~parsedindexvalue_boolArray_6_1; // @[Benes3.scala 36:53]
  wire  _parsedindexvalue_nextIndex_T_509 = parsedindexvalue_calculation_13 == 2'h0 & ~parsedindexvalue_boolArray_6_1; // @[Benes3.scala 36:36]
  wire  _parsedindexvalue_nextIndex_T_510 = parsedindexvalue_calculation_13 == 2'h1; // @[Benes3.scala 37:27]
  wire  _parsedindexvalue_nextIndex_T_512 = parsedindexvalue_calculation_13 == 2'h1 & _parsedindexvalue_nextIndex_T_508; // @[Benes3.scala 37:36]
  wire  _parsedindexvalue_nextIndex_T_513 = parsedindexvalue_calculation_13 == 2'h2; // @[Benes3.scala 38:27]
  wire  _parsedindexvalue_nextIndex_T_515 = parsedindexvalue_calculation_13 == 2'h2 & _parsedindexvalue_nextIndex_T_508; // @[Benes3.scala 38:36]
  wire  _parsedindexvalue_nextIndex_T_516 = parsedindexvalue_calculation_13 == 2'h3; // @[Benes3.scala 39:27]
  wire  _parsedindexvalue_nextIndex_T_518 = parsedindexvalue_calculation_13 == 2'h3 & _parsedindexvalue_nextIndex_T_508; // @[Benes3.scala 39:36]
  wire  _parsedindexvalue_nextIndex_T_521 = _parsedindexvalue_nextIndex_T_507 & parsedindexvalue_boolArray_6_1; // @[Benes3.scala 40:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_523 = parsedindexvalue_nextIndex_12 + 2'h2; // @[Benes3.scala 40:76]
  wire  _parsedindexvalue_nextIndex_T_526 = _parsedindexvalue_nextIndex_T_510 & parsedindexvalue_boolArray_6_1; // @[Benes3.scala 41:36]
  wire  _parsedindexvalue_nextIndex_T_531 = _parsedindexvalue_nextIndex_T_513 & parsedindexvalue_boolArray_6_1; // @[Benes3.scala 42:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_533 = parsedindexvalue_nextIndex_12 - 2'h2; // @[Benes3.scala 42:76]
  wire  _parsedindexvalue_nextIndex_T_536 = _parsedindexvalue_nextIndex_T_516 & parsedindexvalue_boolArray_6_1; // @[Benes3.scala 43:36]
  wire [1:0] _parsedindexvalue_nextIndex_T_539 = _parsedindexvalue_nextIndex_T_536 ? _parsedindexvalue_nextIndex_T_533
     : parsedindexvalue_nextIndex_12; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_540 = _parsedindexvalue_nextIndex_T_531 ? _parsedindexvalue_nextIndex_T_533
     : _parsedindexvalue_nextIndex_T_539; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_541 = _parsedindexvalue_nextIndex_T_526 ? _parsedindexvalue_nextIndex_T_523
     : _parsedindexvalue_nextIndex_T_540; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_542 = _parsedindexvalue_nextIndex_T_521 ? _parsedindexvalue_nextIndex_T_523
     : _parsedindexvalue_nextIndex_T_541; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_543 = _parsedindexvalue_nextIndex_T_518 ? parsedindexvalue_nextIndex_12 :
    _parsedindexvalue_nextIndex_T_542; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_544 = _parsedindexvalue_nextIndex_T_515 ? parsedindexvalue_nextIndex_12 :
    _parsedindexvalue_nextIndex_T_543; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_nextIndex_T_545 = _parsedindexvalue_nextIndex_T_512 ? parsedindexvalue_nextIndex_12 :
    _parsedindexvalue_nextIndex_T_544; // @[Mux.scala 101:16]
  wire [1:0] parsedindexvalue_nextIndex_13 = _parsedindexvalue_nextIndex_T_509 ? parsedindexvalue_nextIndex_12 :
    _parsedindexvalue_nextIndex_T_545; // @[Mux.scala 101:16]
  wire [1:0] _parsedindexvalue_third_stage_T_49 = parsedindexvalue_nextIndex_13 % 2'h2; // @[Benes3.scala 49:61]
  wire [1:0] _parsedindexvalue_third_stage_T_52 = parsedindexvalue_nextIndex_13 + 2'h1; // @[Benes3.scala 49:89]
  wire [1:0] _parsedindexvalue_third_stage_T_54 = parsedindexvalue_nextIndex_13 - 2'h1; // @[Benes3.scala 49:109]
  wire [1:0] _parsedindexvalue_third_stage_T_55 = _parsedindexvalue_third_stage_T_49 == 2'h0 ?
    _parsedindexvalue_third_stage_T_52 : _parsedindexvalue_third_stage_T_54; // @[Benes3.scala 49:47]
  wire [1:0] parsedindexvalue_6 = io_i_mux_bus_3_0[3] ? _parsedindexvalue_third_stage_T_55 :
    parsedindexvalue_nextIndex_13; // @[Benes3.scala 49:24]
  wire [2:0] _T_213 = {{1'd0}, parsedindexvalue_6};
  wire [15:0] _GEN_330 = 3'h0 == _T_213 ? io_i_data_bus2_3 : _GEN_325; // @[Benes3.scala 67:{47,47}]
  wire [15:0] _GEN_331 = 3'h1 == _T_213 ? io_i_data_bus2_3 : _GEN_326; // @[Benes3.scala 67:{47,47}]
  wire [15:0] _GEN_332 = 3'h2 == _T_213 ? io_i_data_bus2_3 : _GEN_327; // @[Benes3.scala 67:{47,47}]
  wire [15:0] _GEN_333 = 3'h3 == _T_213 ? io_i_data_bus2_3 : _GEN_328; // @[Benes3.scala 67:{47,47}]
  wire [15:0] _GEN_335 = ~(|io_i_mux_bus_3_0) ? _GEN_330 : _GEN_325; // @[Benes3.scala 64:49]
  wire [15:0] _GEN_336 = ~(|io_i_mux_bus_3_0) ? _GEN_331 : _GEN_326; // @[Benes3.scala 64:49]
  wire [15:0] _GEN_337 = ~(|io_i_mux_bus_3_0) ? _GEN_332 : _GEN_327; // @[Benes3.scala 64:49]
  wire [15:0] _GEN_338 = ~(|io_i_mux_bus_3_0) ? _GEN_333 : _GEN_328; // @[Benes3.scala 64:49]
  wire [15:0] _GEN_340 = 3'h0 == _T_213 ? io_i_data_bus2_3 : _GEN_335; // @[Benes3.scala 77:{47,47}]
  wire [15:0] _GEN_341 = 3'h1 == _T_213 ? io_i_data_bus2_3 : _GEN_336; // @[Benes3.scala 77:{47,47}]
  wire [15:0] _GEN_342 = 3'h2 == _T_213 ? io_i_data_bus2_3 : _GEN_337; // @[Benes3.scala 77:{47,47}]
  wire [15:0] _GEN_343 = 3'h3 == _T_213 ? io_i_data_bus2_3 : _GEN_338; // @[Benes3.scala 77:{47,47}]
  wire [15:0] _GEN_345 = _T_211 ? _GEN_340 : _GEN_335; // @[Benes3.scala 74:48]
  wire [15:0] _GEN_346 = _T_211 ? _GEN_341 : _GEN_336; // @[Benes3.scala 74:48]
  wire [15:0] _GEN_347 = _T_211 ? _GEN_342 : _GEN_337; // @[Benes3.scala 74:48]
  wire [15:0] _GEN_348 = _T_211 ? _GEN_343 : _GEN_338; // @[Benes3.scala 74:48]
  assign io_o_dist_bus1_0 = io_i_data_bus1_0; // @[Benes3.scala 17:18]
  assign io_o_dist_bus1_1 = io_i_data_bus1_1; // @[Benes3.scala 17:18]
  assign io_o_dist_bus1_2 = io_i_data_bus1_2; // @[Benes3.scala 17:18]
  assign io_o_dist_bus1_3 = io_i_data_bus1_3; // @[Benes3.scala 17:18]
  assign io_o_dist_bus2_0 = io_i_data_bus2_3 != 16'h0 ? _GEN_345 : _GEN_325; // @[Benes3.scala 62:39]
  assign io_o_dist_bus2_1 = io_i_data_bus2_3 != 16'h0 ? _GEN_346 : _GEN_326; // @[Benes3.scala 62:39]
  assign io_o_dist_bus2_2 = io_i_data_bus2_3 != 16'h0 ? _GEN_347 : _GEN_327; // @[Benes3.scala 62:39]
  assign io_o_dist_bus2_3 = io_i_data_bus2_3 != 16'h0 ? _GEN_348 : _GEN_328; // @[Benes3.scala 62:39]
endmodule
module buffer_multiplication(
  input  [15:0] io_buffer1_0,
  input  [15:0] io_buffer1_1,
  input  [15:0] io_buffer1_2,
  input  [15:0] io_buffer1_3,
  input  [15:0] io_buffer2_0,
  input  [15:0] io_buffer2_1,
  input  [15:0] io_buffer2_2,
  input  [15:0] io_buffer2_3,
  output [15:0] io_out_0,
  output [15:0] io_out_1,
  output [15:0] io_out_2,
  output [15:0] io_out_3
);
  wire [31:0] elementMul = io_buffer1_0 * io_buffer2_0; // @[buffer_multiplication.scala 17:42]
  wire [31:0] result_elementMul = io_buffer1_1 * io_buffer2_1; // @[buffer_multiplication.scala 17:42]
  wire [31:0] result_result_elementMul = io_buffer1_2 * io_buffer2_2; // @[buffer_multiplication.scala 17:42]
  wire [31:0] result_result_result_elementMul = io_buffer1_3 * io_buffer2_3; // @[buffer_multiplication.scala 17:42]
  assign io_out_0 = elementMul[15:0]; // @[buffer_multiplication.scala 15:20 19:27]
  assign io_out_1 = result_elementMul[15:0]; // @[buffer_multiplication.scala 15:20 19:27]
  assign io_out_2 = result_result_elementMul[15:0]; // @[buffer_multiplication.scala 15:20 19:27]
  assign io_out_3 = result_result_result_elementMul[15:0]; // @[buffer_multiplication.scala 15:20 19:27]
endmodule
module ReductionMux(
  input  [31:0] io_i_data_0,
  input  [31:0] io_i_data_1,
  output [31:0] io_o_data_0,
  output [31:0] io_o_data_1
);
  assign io_o_data_0 = io_i_data_0; // @[ReductionMux.scala 31:39 33:18 35:18]
  assign io_o_data_1 = io_i_data_1; // @[ReductionMux.scala 37:22]
endmodule
module SimpleAdder(
  input  [31:0] io_A,
  input  [31:0] io_B,
  output [31:0] io_O
);
  assign io_O = io_A + io_B; // @[SimpleAdder.scala 14:18]
endmodule
module EdgeAdderSwitch(
  input         clock,
  input         reset,
  input         io_i_valid,
  input  [63:0] io_i_data_bus_0,
  input  [63:0] io_i_data_bus_1,
  input  [2:0]  io_i_add_en,
  input  [4:0]  io_i_cmd,
  output [31:0] io_o_adder
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] reductionMux_io_i_data_0; // @[EdgeAdderSwitch.scala 19:28]
  wire [31:0] reductionMux_io_i_data_1; // @[EdgeAdderSwitch.scala 19:28]
  wire [31:0] reductionMux_io_o_data_0; // @[EdgeAdderSwitch.scala 19:28]
  wire [31:0] reductionMux_io_o_data_1; // @[EdgeAdderSwitch.scala 19:28]
  wire [31:0] adder32_io_A; // @[EdgeAdderSwitch.scala 23:23]
  wire [31:0] adder32_io_B; // @[EdgeAdderSwitch.scala 23:23]
  wire [31:0] adder32_io_O; // @[EdgeAdderSwitch.scala 23:23]
  reg  r_valid; // @[EdgeAdderSwitch.scala 27:24]
  reg [31:0] r_adder; // @[EdgeAdderSwitch.scala 28:24]
  reg [2:0] r_add_en; // @[EdgeAdderSwitch.scala 31:25]
  wire [31:0] _GEN_3 = 5'h4 == io_i_cmd ? reductionMux_io_o_data_0 : r_adder; // @[EdgeAdderSwitch.scala 38:23 45:17 28:24]
  wire [31:0] _GEN_15 = r_add_en == 3'h0 ? r_adder : adder32_io_O; // @[EdgeAdderSwitch.scala 64:22 65:18 67:18]
  ReductionMux reductionMux ( // @[EdgeAdderSwitch.scala 19:28]
    .io_i_data_0(reductionMux_io_i_data_0),
    .io_i_data_1(reductionMux_io_i_data_1),
    .io_o_data_0(reductionMux_io_o_data_0),
    .io_o_data_1(reductionMux_io_o_data_1)
  );
  SimpleAdder adder32 ( // @[EdgeAdderSwitch.scala 23:23]
    .io_A(adder32_io_A),
    .io_B(adder32_io_B),
    .io_O(adder32_io_O)
  );
  assign io_o_adder = reset ? 32'h0 : _GEN_15; // @[EdgeAdderSwitch.scala 59:14 60:16]
  assign reductionMux_io_i_data_0 = io_i_data_bus_0[31:0]; // @[EdgeAdderSwitch.scala 20:26]
  assign reductionMux_io_i_data_1 = io_i_data_bus_1[31:0]; // @[EdgeAdderSwitch.scala 20:26]
  assign adder32_io_A = reductionMux_io_o_data_1; // @[EdgeAdderSwitch.scala 24:16]
  assign adder32_io_B = reductionMux_io_o_data_0; // @[EdgeAdderSwitch.scala 25:16]
  always @(posedge clock) begin
    if (reset) begin // @[EdgeAdderSwitch.scala 27:24]
      r_valid <= 1'h0; // @[EdgeAdderSwitch.scala 27:24]
    end else begin
      r_valid <= io_i_valid; // @[EdgeAdderSwitch.scala 27:24]
    end
    if (reset) begin // @[EdgeAdderSwitch.scala 28:24]
      r_adder <= 32'h0; // @[EdgeAdderSwitch.scala 28:24]
    end else if (reset) begin // @[EdgeAdderSwitch.scala 33:14]
      r_adder <= 32'h0; // @[EdgeAdderSwitch.scala 34:13]
    end else if (r_valid) begin // @[EdgeAdderSwitch.scala 37:25]
      if (5'h3 == io_i_cmd) begin // @[EdgeAdderSwitch.scala 38:23]
        r_adder <= reductionMux_io_o_data_1; // @[EdgeAdderSwitch.scala 40:17]
      end else begin
        r_adder <= _GEN_3;
      end
    end
    if (reset) begin // @[EdgeAdderSwitch.scala 31:25]
      r_add_en <= 3'h0; // @[EdgeAdderSwitch.scala 31:25]
    end else begin
      r_add_en <= io_i_add_en; // @[EdgeAdderSwitch.scala 31:25]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  r_adder = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  r_add_en = _RAND_2[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Fan4(
  input         clock,
  input         reset,
  input         io_i_valid,
  input  [31:0] io_i_data_bus_0,
  input  [31:0] io_i_data_bus_1,
  input  [31:0] io_i_data_bus_2,
  input  [31:0] io_i_data_bus_3,
  input         io_i_add_en_bus_0,
  input         io_i_add_en_bus_1,
  input         io_i_add_en_bus_2,
  input  [2:0]  io_i_cmd_bus_0,
  input  [2:0]  io_i_cmd_bus_1,
  input  [2:0]  io_i_cmd_bus_2,
  output [31:0] io_o_adder_0,
  output [31:0] io_o_adder_1,
  output [31:0] io_o_adder_2
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  my_adder_0_clock; // @[FanNetwork.scala 119:28]
  wire  my_adder_0_reset; // @[FanNetwork.scala 119:28]
  wire  my_adder_0_io_i_valid; // @[FanNetwork.scala 119:28]
  wire [63:0] my_adder_0_io_i_data_bus_0; // @[FanNetwork.scala 119:28]
  wire [63:0] my_adder_0_io_i_data_bus_1; // @[FanNetwork.scala 119:28]
  wire [2:0] my_adder_0_io_i_add_en; // @[FanNetwork.scala 119:28]
  wire [4:0] my_adder_0_io_i_cmd; // @[FanNetwork.scala 119:28]
  wire [31:0] my_adder_0_io_o_adder; // @[FanNetwork.scala 119:28]
  wire  my_adder_1_clock; // @[FanNetwork.scala 132:28]
  wire  my_adder_1_reset; // @[FanNetwork.scala 132:28]
  wire  my_adder_1_io_i_valid; // @[FanNetwork.scala 132:28]
  wire [63:0] my_adder_1_io_i_data_bus_0; // @[FanNetwork.scala 132:28]
  wire [63:0] my_adder_1_io_i_data_bus_1; // @[FanNetwork.scala 132:28]
  wire [2:0] my_adder_1_io_i_add_en; // @[FanNetwork.scala 132:28]
  wire [4:0] my_adder_1_io_i_cmd; // @[FanNetwork.scala 132:28]
  wire [31:0] my_adder_1_io_o_adder; // @[FanNetwork.scala 132:28]
  wire  my_adder_2_clock; // @[FanNetwork.scala 145:28]
  wire  my_adder_2_reset; // @[FanNetwork.scala 145:28]
  wire  my_adder_2_io_i_valid; // @[FanNetwork.scala 145:28]
  wire [63:0] my_adder_2_io_i_data_bus_0; // @[FanNetwork.scala 145:28]
  wire [63:0] my_adder_2_io_i_data_bus_1; // @[FanNetwork.scala 145:28]
  wire [2:0] my_adder_2_io_i_add_en; // @[FanNetwork.scala 145:28]
  wire [4:0] my_adder_2_io_i_cmd; // @[FanNetwork.scala 145:28]
  wire [31:0] my_adder_2_io_o_adder; // @[FanNetwork.scala 145:28]
  reg  r_valid_0; // @[FanNetwork.scala 30:26]
  reg  r_valid_1; // @[FanNetwork.scala 30:26]
  wire [63:0] w_fan_lvl_0_0 = {{32'd0}, my_adder_0_io_o_adder};
  wire [63:0] w_fan_lvl_0_1 = {{32'd0}, my_adder_2_io_o_adder};
  EdgeAdderSwitch my_adder_0 ( // @[FanNetwork.scala 119:28]
    .clock(my_adder_0_clock),
    .reset(my_adder_0_reset),
    .io_i_valid(my_adder_0_io_i_valid),
    .io_i_data_bus_0(my_adder_0_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_0_io_i_data_bus_1),
    .io_i_add_en(my_adder_0_io_i_add_en),
    .io_i_cmd(my_adder_0_io_i_cmd),
    .io_o_adder(my_adder_0_io_o_adder)
  );
  EdgeAdderSwitch my_adder_1 ( // @[FanNetwork.scala 132:28]
    .clock(my_adder_1_clock),
    .reset(my_adder_1_reset),
    .io_i_valid(my_adder_1_io_i_valid),
    .io_i_data_bus_0(my_adder_1_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_1_io_i_data_bus_1),
    .io_i_add_en(my_adder_1_io_i_add_en),
    .io_i_cmd(my_adder_1_io_i_cmd),
    .io_o_adder(my_adder_1_io_o_adder)
  );
  EdgeAdderSwitch my_adder_2 ( // @[FanNetwork.scala 145:28]
    .clock(my_adder_2_clock),
    .reset(my_adder_2_reset),
    .io_i_valid(my_adder_2_io_i_valid),
    .io_i_data_bus_0(my_adder_2_io_i_data_bus_0),
    .io_i_data_bus_1(my_adder_2_io_i_data_bus_1),
    .io_i_add_en(my_adder_2_io_i_add_en),
    .io_i_cmd(my_adder_2_io_i_cmd),
    .io_o_adder(my_adder_2_io_o_adder)
  );
  assign io_o_adder_0 = w_fan_lvl_0_0[31:0]; // @[FanNetwork.scala 207:19]
  assign io_o_adder_1 = my_adder_1_io_o_adder; // @[FanNetwork.scala 208:19]
  assign io_o_adder_2 = w_fan_lvl_0_1[31:0]; // @[FanNetwork.scala 209:19]
  assign my_adder_0_clock = clock;
  assign my_adder_0_reset = reset;
  assign my_adder_0_io_i_valid = r_valid_0; // @[FanNetwork.scala 121:27]
  assign my_adder_0_io_i_data_bus_0 = {{32'd0}, io_i_data_bus_1}; // @[FanNetwork.scala 122:30]
  assign my_adder_0_io_i_data_bus_1 = {{32'd0}, io_i_data_bus_0}; // @[FanNetwork.scala 122:30]
  assign my_adder_0_io_i_add_en = {{2'd0}, io_i_add_en_bus_0}; // @[FanNetwork.scala 123:28]
  assign my_adder_0_io_i_cmd = {{2'd0}, io_i_cmd_bus_0}; // @[FanNetwork.scala 124:25]
  assign my_adder_1_clock = clock;
  assign my_adder_1_reset = reset;
  assign my_adder_1_io_i_valid = r_valid_1; // @[FanNetwork.scala 134:27]
  assign my_adder_1_io_i_data_bus_0 = {{32'd0}, my_adder_2_io_o_adder}; // @[FanNetwork.scala 135:{40,40}]
  assign my_adder_1_io_i_data_bus_1 = {{32'd0}, my_adder_0_io_o_adder}; // @[FanNetwork.scala 135:{40,40}]
  assign my_adder_1_io_i_add_en = {{2'd0}, io_i_add_en_bus_2}; // @[FanNetwork.scala 136:28]
  assign my_adder_1_io_i_cmd = {{2'd0}, io_i_cmd_bus_2}; // @[FanNetwork.scala 137:26]
  assign my_adder_2_clock = clock;
  assign my_adder_2_reset = reset;
  assign my_adder_2_io_i_valid = r_valid_0; // @[FanNetwork.scala 147:27]
  assign my_adder_2_io_i_data_bus_0 = {{32'd0}, io_i_data_bus_3}; // @[FanNetwork.scala 148:30]
  assign my_adder_2_io_i_data_bus_1 = {{32'd0}, io_i_data_bus_2}; // @[FanNetwork.scala 148:30]
  assign my_adder_2_io_i_add_en = {{2'd0}, io_i_add_en_bus_1}; // @[FanNetwork.scala 149:28]
  assign my_adder_2_io_i_cmd = {{2'd0}, io_i_cmd_bus_1}; // @[FanNetwork.scala 150:25]
  always @(posedge clock) begin
    if (reset) begin // @[FanNetwork.scala 30:26]
      r_valid_0 <= 1'h0; // @[FanNetwork.scala 30:26]
    end else begin
      r_valid_0 <= io_i_valid;
    end
    if (reset) begin // @[FanNetwork.scala 30:26]
      r_valid_1 <= 1'h0; // @[FanNetwork.scala 30:26]
    end else begin
      r_valid_1 <= r_valid_0; // @[FanNetwork.scala 114:24]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_valid_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  r_valid_1 = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module flexdpecom4(
  input         clock,
  input         reset,
  input         io_i_data_valid,
  input  [15:0] io_i_data_bus_0,
  input  [15:0] io_i_data_bus_1,
  input  [15:0] io_i_data_bus_2,
  input  [15:0] io_i_data_bus_3,
  input  [15:0] io_i_data_bus2_0,
  input  [15:0] io_i_data_bus2_1,
  input  [15:0] io_i_data_bus2_2,
  input  [15:0] io_i_data_bus2_3,
  input  [4:0]  io_i_vn_0,
  input  [4:0]  io_i_vn_1,
  input  [4:0]  io_i_vn_2,
  input  [4:0]  io_i_vn_3,
  output [15:0] io_o_adder_0,
  output [15:0] io_o_adder_1,
  output [15:0] io_o_adder_2,
  input  [3:0]  io_i_mux_bus_0_0,
  input  [3:0]  io_i_mux_bus_0_1,
  input  [3:0]  io_i_mux_bus_0_2,
  input  [3:0]  io_i_mux_bus_0_3,
  input  [3:0]  io_i_mux_bus_1_0,
  input  [3:0]  io_i_mux_bus_1_1,
  input  [3:0]  io_i_mux_bus_1_2,
  input  [3:0]  io_i_mux_bus_2_0,
  input  [3:0]  io_i_mux_bus_2_1,
  input  [3:0]  io_i_mux_bus_3_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
`endif // RANDOMIZE_REG_INIT
  wire  my_controller_clock; // @[FlexDPE.scala 55:31]
  wire  my_controller_reset; // @[FlexDPE.scala 55:31]
  wire [4:0] my_controller_io_i_vn_0; // @[FlexDPE.scala 55:31]
  wire [4:0] my_controller_io_i_vn_1; // @[FlexDPE.scala 55:31]
  wire [4:0] my_controller_io_i_vn_2; // @[FlexDPE.scala 55:31]
  wire [4:0] my_controller_io_i_vn_3; // @[FlexDPE.scala 55:31]
  wire  my_controller_io_i_data_valid; // @[FlexDPE.scala 55:31]
  wire  my_controller_io_o_reduction_add_0; // @[FlexDPE.scala 55:31]
  wire  my_controller_io_o_reduction_add_1; // @[FlexDPE.scala 55:31]
  wire  my_controller_io_o_reduction_add_2; // @[FlexDPE.scala 55:31]
  wire [2:0] my_controller_io_o_reduction_cmd_0; // @[FlexDPE.scala 55:31]
  wire [2:0] my_controller_io_o_reduction_cmd_1; // @[FlexDPE.scala 55:31]
  wire [2:0] my_controller_io_o_reduction_cmd_2; // @[FlexDPE.scala 55:31]
  wire  my_controller_io_o_reduction_valid; // @[FlexDPE.scala 55:31]
  wire [15:0] my_Benes_io_i_data_bus2_0; // @[FlexDPE.scala 64:26]
  wire [15:0] my_Benes_io_i_data_bus2_1; // @[FlexDPE.scala 64:26]
  wire [15:0] my_Benes_io_i_data_bus2_2; // @[FlexDPE.scala 64:26]
  wire [15:0] my_Benes_io_i_data_bus2_3; // @[FlexDPE.scala 64:26]
  wire [15:0] my_Benes_io_i_data_bus1_0; // @[FlexDPE.scala 64:26]
  wire [15:0] my_Benes_io_i_data_bus1_1; // @[FlexDPE.scala 64:26]
  wire [15:0] my_Benes_io_i_data_bus1_2; // @[FlexDPE.scala 64:26]
  wire [15:0] my_Benes_io_i_data_bus1_3; // @[FlexDPE.scala 64:26]
  wire [3:0] my_Benes_io_i_mux_bus_0_0; // @[FlexDPE.scala 64:26]
  wire [3:0] my_Benes_io_i_mux_bus_0_1; // @[FlexDPE.scala 64:26]
  wire [3:0] my_Benes_io_i_mux_bus_0_2; // @[FlexDPE.scala 64:26]
  wire [3:0] my_Benes_io_i_mux_bus_0_3; // @[FlexDPE.scala 64:26]
  wire [3:0] my_Benes_io_i_mux_bus_1_0; // @[FlexDPE.scala 64:26]
  wire [3:0] my_Benes_io_i_mux_bus_1_1; // @[FlexDPE.scala 64:26]
  wire [3:0] my_Benes_io_i_mux_bus_1_2; // @[FlexDPE.scala 64:26]
  wire [3:0] my_Benes_io_i_mux_bus_2_0; // @[FlexDPE.scala 64:26]
  wire [3:0] my_Benes_io_i_mux_bus_2_1; // @[FlexDPE.scala 64:26]
  wire [3:0] my_Benes_io_i_mux_bus_3_0; // @[FlexDPE.scala 64:26]
  wire [15:0] my_Benes_io_o_dist_bus1_0; // @[FlexDPE.scala 64:26]
  wire [15:0] my_Benes_io_o_dist_bus1_1; // @[FlexDPE.scala 64:26]
  wire [15:0] my_Benes_io_o_dist_bus1_2; // @[FlexDPE.scala 64:26]
  wire [15:0] my_Benes_io_o_dist_bus1_3; // @[FlexDPE.scala 64:26]
  wire [15:0] my_Benes_io_o_dist_bus2_0; // @[FlexDPE.scala 64:26]
  wire [15:0] my_Benes_io_o_dist_bus2_1; // @[FlexDPE.scala 64:26]
  wire [15:0] my_Benes_io_o_dist_bus2_2; // @[FlexDPE.scala 64:26]
  wire [15:0] my_Benes_io_o_dist_bus2_3; // @[FlexDPE.scala 64:26]
  wire [15:0] buffer_mult_io_buffer1_0; // @[FlexDPE.scala 75:30]
  wire [15:0] buffer_mult_io_buffer1_1; // @[FlexDPE.scala 75:30]
  wire [15:0] buffer_mult_io_buffer1_2; // @[FlexDPE.scala 75:30]
  wire [15:0] buffer_mult_io_buffer1_3; // @[FlexDPE.scala 75:30]
  wire [15:0] buffer_mult_io_buffer2_0; // @[FlexDPE.scala 75:30]
  wire [15:0] buffer_mult_io_buffer2_1; // @[FlexDPE.scala 75:30]
  wire [15:0] buffer_mult_io_buffer2_2; // @[FlexDPE.scala 75:30]
  wire [15:0] buffer_mult_io_buffer2_3; // @[FlexDPE.scala 75:30]
  wire [15:0] buffer_mult_io_out_0; // @[FlexDPE.scala 75:30]
  wire [15:0] buffer_mult_io_out_1; // @[FlexDPE.scala 75:30]
  wire [15:0] buffer_mult_io_out_2; // @[FlexDPE.scala 75:30]
  wire [15:0] buffer_mult_io_out_3; // @[FlexDPE.scala 75:30]
  wire  my_fan_network_clock; // @[FlexDPE.scala 87:32]
  wire  my_fan_network_reset; // @[FlexDPE.scala 87:32]
  wire  my_fan_network_io_i_valid; // @[FlexDPE.scala 87:32]
  wire [31:0] my_fan_network_io_i_data_bus_0; // @[FlexDPE.scala 87:32]
  wire [31:0] my_fan_network_io_i_data_bus_1; // @[FlexDPE.scala 87:32]
  wire [31:0] my_fan_network_io_i_data_bus_2; // @[FlexDPE.scala 87:32]
  wire [31:0] my_fan_network_io_i_data_bus_3; // @[FlexDPE.scala 87:32]
  wire  my_fan_network_io_i_add_en_bus_0; // @[FlexDPE.scala 87:32]
  wire  my_fan_network_io_i_add_en_bus_1; // @[FlexDPE.scala 87:32]
  wire  my_fan_network_io_i_add_en_bus_2; // @[FlexDPE.scala 87:32]
  wire [2:0] my_fan_network_io_i_cmd_bus_0; // @[FlexDPE.scala 87:32]
  wire [2:0] my_fan_network_io_i_cmd_bus_1; // @[FlexDPE.scala 87:32]
  wire [2:0] my_fan_network_io_i_cmd_bus_2; // @[FlexDPE.scala 87:32]
  wire [31:0] my_fan_network_io_o_adder_0; // @[FlexDPE.scala 87:32]
  wire [31:0] my_fan_network_io_o_adder_1; // @[FlexDPE.scala 87:32]
  wire [31:0] my_fan_network_io_o_adder_2; // @[FlexDPE.scala 87:32]
  reg [14:0] r_mult_0; // @[FlexDPE.scala 32:26]
  reg [14:0] r_mult_1; // @[FlexDPE.scala 32:26]
  reg [14:0] r_mult_2; // @[FlexDPE.scala 32:26]
  reg [14:0] r_mult_3; // @[FlexDPE.scala 32:26]
  reg [15:0] matrix_0_0; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_0_1; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_0_2; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_0_3; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_0_4; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_0_5; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_0_6; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_0_7; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_1_0; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_1_1; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_1_2; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_1_3; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_1_4; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_1_5; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_1_6; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_1_7; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_2_0; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_2_1; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_2_2; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_2_3; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_2_4; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_2_5; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_2_6; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_2_7; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_3_0; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_3_1; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_3_2; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_3_3; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_3_4; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_3_5; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_3_6; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_3_7; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_4_0; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_4_1; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_4_2; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_4_3; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_4_4; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_4_5; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_4_6; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_4_7; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_5_0; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_5_1; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_5_2; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_5_3; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_5_4; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_5_5; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_5_6; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_5_7; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_6_0; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_6_1; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_6_2; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_6_3; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_6_4; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_6_5; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_6_6; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_6_7; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_7_0; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_7_1; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_7_2; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_7_3; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_7_4; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_7_5; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_7_6; // @[FlexDPE.scala 33:21]
  reg [15:0] matrix_7_7; // @[FlexDPE.scala 33:21]
  wire [15:0] _GEN_0 = reset ? 16'h0 : buffer_mult_io_out_0; // @[FlexDPE.scala 32:{26,26} 81:14]
  wire [15:0] _GEN_1 = reset ? 16'h0 : buffer_mult_io_out_1; // @[FlexDPE.scala 32:{26,26} 81:14]
  wire [15:0] _GEN_2 = reset ? 16'h0 : buffer_mult_io_out_2; // @[FlexDPE.scala 32:{26,26} 81:14]
  wire [15:0] _GEN_3 = reset ? 16'h0 : buffer_mult_io_out_3; // @[FlexDPE.scala 32:{26,26} 81:14]
  fancontrol4 my_controller ( // @[FlexDPE.scala 55:31]
    .clock(my_controller_clock),
    .reset(my_controller_reset),
    .io_i_vn_0(my_controller_io_i_vn_0),
    .io_i_vn_1(my_controller_io_i_vn_1),
    .io_i_vn_2(my_controller_io_i_vn_2),
    .io_i_vn_3(my_controller_io_i_vn_3),
    .io_i_data_valid(my_controller_io_i_data_valid),
    .io_o_reduction_add_0(my_controller_io_o_reduction_add_0),
    .io_o_reduction_add_1(my_controller_io_o_reduction_add_1),
    .io_o_reduction_add_2(my_controller_io_o_reduction_add_2),
    .io_o_reduction_cmd_0(my_controller_io_o_reduction_cmd_0),
    .io_o_reduction_cmd_1(my_controller_io_o_reduction_cmd_1),
    .io_o_reduction_cmd_2(my_controller_io_o_reduction_cmd_2),
    .io_o_reduction_valid(my_controller_io_o_reduction_valid)
  );
  Benes3 my_Benes ( // @[FlexDPE.scala 64:26]
    .io_i_data_bus2_0(my_Benes_io_i_data_bus2_0),
    .io_i_data_bus2_1(my_Benes_io_i_data_bus2_1),
    .io_i_data_bus2_2(my_Benes_io_i_data_bus2_2),
    .io_i_data_bus2_3(my_Benes_io_i_data_bus2_3),
    .io_i_data_bus1_0(my_Benes_io_i_data_bus1_0),
    .io_i_data_bus1_1(my_Benes_io_i_data_bus1_1),
    .io_i_data_bus1_2(my_Benes_io_i_data_bus1_2),
    .io_i_data_bus1_3(my_Benes_io_i_data_bus1_3),
    .io_i_mux_bus_0_0(my_Benes_io_i_mux_bus_0_0),
    .io_i_mux_bus_0_1(my_Benes_io_i_mux_bus_0_1),
    .io_i_mux_bus_0_2(my_Benes_io_i_mux_bus_0_2),
    .io_i_mux_bus_0_3(my_Benes_io_i_mux_bus_0_3),
    .io_i_mux_bus_1_0(my_Benes_io_i_mux_bus_1_0),
    .io_i_mux_bus_1_1(my_Benes_io_i_mux_bus_1_1),
    .io_i_mux_bus_1_2(my_Benes_io_i_mux_bus_1_2),
    .io_i_mux_bus_2_0(my_Benes_io_i_mux_bus_2_0),
    .io_i_mux_bus_2_1(my_Benes_io_i_mux_bus_2_1),
    .io_i_mux_bus_3_0(my_Benes_io_i_mux_bus_3_0),
    .io_o_dist_bus1_0(my_Benes_io_o_dist_bus1_0),
    .io_o_dist_bus1_1(my_Benes_io_o_dist_bus1_1),
    .io_o_dist_bus1_2(my_Benes_io_o_dist_bus1_2),
    .io_o_dist_bus1_3(my_Benes_io_o_dist_bus1_3),
    .io_o_dist_bus2_0(my_Benes_io_o_dist_bus2_0),
    .io_o_dist_bus2_1(my_Benes_io_o_dist_bus2_1),
    .io_o_dist_bus2_2(my_Benes_io_o_dist_bus2_2),
    .io_o_dist_bus2_3(my_Benes_io_o_dist_bus2_3)
  );
  buffer_multiplication buffer_mult ( // @[FlexDPE.scala 75:30]
    .io_buffer1_0(buffer_mult_io_buffer1_0),
    .io_buffer1_1(buffer_mult_io_buffer1_1),
    .io_buffer1_2(buffer_mult_io_buffer1_2),
    .io_buffer1_3(buffer_mult_io_buffer1_3),
    .io_buffer2_0(buffer_mult_io_buffer2_0),
    .io_buffer2_1(buffer_mult_io_buffer2_1),
    .io_buffer2_2(buffer_mult_io_buffer2_2),
    .io_buffer2_3(buffer_mult_io_buffer2_3),
    .io_out_0(buffer_mult_io_out_0),
    .io_out_1(buffer_mult_io_out_1),
    .io_out_2(buffer_mult_io_out_2),
    .io_out_3(buffer_mult_io_out_3)
  );
  Fan4 my_fan_network ( // @[FlexDPE.scala 87:32]
    .clock(my_fan_network_clock),
    .reset(my_fan_network_reset),
    .io_i_valid(my_fan_network_io_i_valid),
    .io_i_data_bus_0(my_fan_network_io_i_data_bus_0),
    .io_i_data_bus_1(my_fan_network_io_i_data_bus_1),
    .io_i_data_bus_2(my_fan_network_io_i_data_bus_2),
    .io_i_data_bus_3(my_fan_network_io_i_data_bus_3),
    .io_i_add_en_bus_0(my_fan_network_io_i_add_en_bus_0),
    .io_i_add_en_bus_1(my_fan_network_io_i_add_en_bus_1),
    .io_i_add_en_bus_2(my_fan_network_io_i_add_en_bus_2),
    .io_i_cmd_bus_0(my_fan_network_io_i_cmd_bus_0),
    .io_i_cmd_bus_1(my_fan_network_io_i_cmd_bus_1),
    .io_i_cmd_bus_2(my_fan_network_io_i_cmd_bus_2),
    .io_o_adder_0(my_fan_network_io_o_adder_0),
    .io_o_adder_1(my_fan_network_io_o_adder_1),
    .io_o_adder_2(my_fan_network_io_o_adder_2)
  );
  assign io_o_adder_0 = my_fan_network_io_o_adder_0[15:0]; // @[FlexDPE.scala 96:16]
  assign io_o_adder_1 = my_fan_network_io_o_adder_1[15:0]; // @[FlexDPE.scala 96:16]
  assign io_o_adder_2 = my_fan_network_io_o_adder_2[15:0]; // @[FlexDPE.scala 96:16]
  assign my_controller_clock = clock;
  assign my_controller_reset = reset;
  assign my_controller_io_i_vn_0 = io_i_vn_0; // @[FlexDPE.scala 57:27]
  assign my_controller_io_i_vn_1 = io_i_vn_1; // @[FlexDPE.scala 57:27]
  assign my_controller_io_i_vn_2 = io_i_vn_2; // @[FlexDPE.scala 57:27]
  assign my_controller_io_i_vn_3 = io_i_vn_3; // @[FlexDPE.scala 57:27]
  assign my_controller_io_i_data_valid = io_i_data_valid; // @[FlexDPE.scala 59:35]
  assign my_Benes_io_i_data_bus2_0 = io_i_data_bus2_0; // @[FlexDPE.scala 67:29]
  assign my_Benes_io_i_data_bus2_1 = io_i_data_bus2_1; // @[FlexDPE.scala 67:29]
  assign my_Benes_io_i_data_bus2_2 = io_i_data_bus2_2; // @[FlexDPE.scala 67:29]
  assign my_Benes_io_i_data_bus2_3 = io_i_data_bus2_3; // @[FlexDPE.scala 67:29]
  assign my_Benes_io_i_data_bus1_0 = io_i_data_bus_0; // @[FlexDPE.scala 66:29]
  assign my_Benes_io_i_data_bus1_1 = io_i_data_bus_1; // @[FlexDPE.scala 66:29]
  assign my_Benes_io_i_data_bus1_2 = io_i_data_bus_2; // @[FlexDPE.scala 66:29]
  assign my_Benes_io_i_data_bus1_3 = io_i_data_bus_3; // @[FlexDPE.scala 66:29]
  assign my_Benes_io_i_mux_bus_0_0 = io_i_mux_bus_0_0; // @[FlexDPE.scala 68:27]
  assign my_Benes_io_i_mux_bus_0_1 = io_i_mux_bus_0_1; // @[FlexDPE.scala 68:27]
  assign my_Benes_io_i_mux_bus_0_2 = io_i_mux_bus_0_2; // @[FlexDPE.scala 68:27]
  assign my_Benes_io_i_mux_bus_0_3 = io_i_mux_bus_0_3; // @[FlexDPE.scala 68:27]
  assign my_Benes_io_i_mux_bus_1_0 = io_i_mux_bus_1_0; // @[FlexDPE.scala 68:27]
  assign my_Benes_io_i_mux_bus_1_1 = io_i_mux_bus_1_1; // @[FlexDPE.scala 68:27]
  assign my_Benes_io_i_mux_bus_1_2 = io_i_mux_bus_1_2; // @[FlexDPE.scala 68:27]
  assign my_Benes_io_i_mux_bus_2_0 = io_i_mux_bus_2_0; // @[FlexDPE.scala 68:27]
  assign my_Benes_io_i_mux_bus_2_1 = io_i_mux_bus_2_1; // @[FlexDPE.scala 68:27]
  assign my_Benes_io_i_mux_bus_3_0 = io_i_mux_bus_3_0; // @[FlexDPE.scala 68:27]
  assign buffer_mult_io_buffer1_0 = my_Benes_io_o_dist_bus1_0; // @[FlexDPE.scala 78:30]
  assign buffer_mult_io_buffer1_1 = my_Benes_io_o_dist_bus1_1; // @[FlexDPE.scala 78:30]
  assign buffer_mult_io_buffer1_2 = my_Benes_io_o_dist_bus1_2; // @[FlexDPE.scala 78:30]
  assign buffer_mult_io_buffer1_3 = my_Benes_io_o_dist_bus1_3; // @[FlexDPE.scala 78:30]
  assign buffer_mult_io_buffer2_0 = my_Benes_io_o_dist_bus2_0; // @[FlexDPE.scala 79:30]
  assign buffer_mult_io_buffer2_1 = my_Benes_io_o_dist_bus2_1; // @[FlexDPE.scala 79:30]
  assign buffer_mult_io_buffer2_2 = my_Benes_io_o_dist_bus2_2; // @[FlexDPE.scala 79:30]
  assign buffer_mult_io_buffer2_3 = my_Benes_io_o_dist_bus2_3; // @[FlexDPE.scala 79:30]
  assign my_fan_network_clock = clock;
  assign my_fan_network_reset = reset;
  assign my_fan_network_io_i_valid = my_controller_io_o_reduction_valid; // @[FlexDPE.scala 89:31]
  assign my_fan_network_io_i_data_bus_0 = {{17'd0}, r_mult_0}; // @[FlexDPE.scala 90:34]
  assign my_fan_network_io_i_data_bus_1 = {{17'd0}, r_mult_1}; // @[FlexDPE.scala 90:34]
  assign my_fan_network_io_i_data_bus_2 = {{17'd0}, r_mult_2}; // @[FlexDPE.scala 90:34]
  assign my_fan_network_io_i_data_bus_3 = {{17'd0}, r_mult_3}; // @[FlexDPE.scala 90:34]
  assign my_fan_network_io_i_add_en_bus_0 = my_controller_io_o_reduction_add_0; // @[FlexDPE.scala 91:36]
  assign my_fan_network_io_i_add_en_bus_1 = my_controller_io_o_reduction_add_1; // @[FlexDPE.scala 91:36]
  assign my_fan_network_io_i_add_en_bus_2 = my_controller_io_o_reduction_add_2; // @[FlexDPE.scala 91:36]
  assign my_fan_network_io_i_cmd_bus_0 = my_controller_io_o_reduction_cmd_0; // @[FlexDPE.scala 92:33]
  assign my_fan_network_io_i_cmd_bus_1 = my_controller_io_o_reduction_cmd_1; // @[FlexDPE.scala 92:33]
  assign my_fan_network_io_i_cmd_bus_2 = my_controller_io_o_reduction_cmd_2; // @[FlexDPE.scala 92:33]
  always @(posedge clock) begin
    r_mult_0 <= _GEN_0[14:0]; // @[FlexDPE.scala 32:{26,26} 81:14]
    r_mult_1 <= _GEN_1[14:0]; // @[FlexDPE.scala 32:{26,26} 81:14]
    r_mult_2 <= _GEN_2[14:0]; // @[FlexDPE.scala 32:{26,26} 81:14]
    r_mult_3 <= _GEN_3[14:0]; // @[FlexDPE.scala 32:{26,26} 81:14]
    matrix_0_0 <= matrix_0_0; // @[FlexDPE.scala 33:21]
    matrix_0_1 <= matrix_0_1; // @[FlexDPE.scala 33:21]
    matrix_0_2 <= matrix_0_2; // @[FlexDPE.scala 33:21]
    matrix_0_3 <= matrix_0_3; // @[FlexDPE.scala 33:21]
    matrix_0_4 <= matrix_0_4; // @[FlexDPE.scala 33:21]
    matrix_0_5 <= matrix_0_5; // @[FlexDPE.scala 33:21]
    matrix_0_6 <= matrix_0_6; // @[FlexDPE.scala 33:21]
    matrix_0_7 <= matrix_0_7; // @[FlexDPE.scala 33:21]
    matrix_1_0 <= matrix_1_0; // @[FlexDPE.scala 33:21]
    matrix_1_1 <= matrix_1_1; // @[FlexDPE.scala 33:21]
    matrix_1_2 <= matrix_1_2; // @[FlexDPE.scala 33:21]
    matrix_1_3 <= matrix_1_3; // @[FlexDPE.scala 33:21]
    matrix_1_4 <= matrix_1_4; // @[FlexDPE.scala 33:21]
    matrix_1_5 <= matrix_1_5; // @[FlexDPE.scala 33:21]
    matrix_1_6 <= matrix_1_6; // @[FlexDPE.scala 33:21]
    matrix_1_7 <= matrix_1_7; // @[FlexDPE.scala 33:21]
    matrix_2_0 <= matrix_2_0; // @[FlexDPE.scala 33:21]
    matrix_2_1 <= matrix_2_1; // @[FlexDPE.scala 33:21]
    matrix_2_2 <= matrix_2_2; // @[FlexDPE.scala 33:21]
    matrix_2_3 <= matrix_2_3; // @[FlexDPE.scala 33:21]
    matrix_2_4 <= matrix_2_4; // @[FlexDPE.scala 33:21]
    matrix_2_5 <= matrix_2_5; // @[FlexDPE.scala 33:21]
    matrix_2_6 <= matrix_2_6; // @[FlexDPE.scala 33:21]
    matrix_2_7 <= matrix_2_7; // @[FlexDPE.scala 33:21]
    matrix_3_0 <= matrix_3_0; // @[FlexDPE.scala 33:21]
    matrix_3_1 <= matrix_3_1; // @[FlexDPE.scala 33:21]
    matrix_3_2 <= matrix_3_2; // @[FlexDPE.scala 33:21]
    matrix_3_3 <= matrix_3_3; // @[FlexDPE.scala 33:21]
    matrix_3_4 <= matrix_3_4; // @[FlexDPE.scala 33:21]
    matrix_3_5 <= matrix_3_5; // @[FlexDPE.scala 33:21]
    matrix_3_6 <= matrix_3_6; // @[FlexDPE.scala 33:21]
    matrix_3_7 <= matrix_3_7; // @[FlexDPE.scala 33:21]
    matrix_4_0 <= matrix_4_0; // @[FlexDPE.scala 33:21]
    matrix_4_1 <= matrix_4_1; // @[FlexDPE.scala 33:21]
    matrix_4_2 <= matrix_4_2; // @[FlexDPE.scala 33:21]
    matrix_4_3 <= matrix_4_3; // @[FlexDPE.scala 33:21]
    matrix_4_4 <= matrix_4_4; // @[FlexDPE.scala 33:21]
    matrix_4_5 <= matrix_4_5; // @[FlexDPE.scala 33:21]
    matrix_4_6 <= matrix_4_6; // @[FlexDPE.scala 33:21]
    matrix_4_7 <= matrix_4_7; // @[FlexDPE.scala 33:21]
    matrix_5_0 <= matrix_5_0; // @[FlexDPE.scala 33:21]
    matrix_5_1 <= matrix_5_1; // @[FlexDPE.scala 33:21]
    matrix_5_2 <= matrix_5_2; // @[FlexDPE.scala 33:21]
    matrix_5_3 <= matrix_5_3; // @[FlexDPE.scala 33:21]
    matrix_5_4 <= matrix_5_4; // @[FlexDPE.scala 33:21]
    matrix_5_5 <= matrix_5_5; // @[FlexDPE.scala 33:21]
    matrix_5_6 <= matrix_5_6; // @[FlexDPE.scala 33:21]
    matrix_5_7 <= matrix_5_7; // @[FlexDPE.scala 33:21]
    matrix_6_0 <= matrix_6_0; // @[FlexDPE.scala 33:21]
    matrix_6_1 <= matrix_6_1; // @[FlexDPE.scala 33:21]
    matrix_6_2 <= matrix_6_2; // @[FlexDPE.scala 33:21]
    matrix_6_3 <= matrix_6_3; // @[FlexDPE.scala 33:21]
    matrix_6_4 <= matrix_6_4; // @[FlexDPE.scala 33:21]
    matrix_6_5 <= matrix_6_5; // @[FlexDPE.scala 33:21]
    matrix_6_6 <= matrix_6_6; // @[FlexDPE.scala 33:21]
    matrix_6_7 <= matrix_6_7; // @[FlexDPE.scala 33:21]
    matrix_7_0 <= matrix_7_0; // @[FlexDPE.scala 33:21]
    matrix_7_1 <= matrix_7_1; // @[FlexDPE.scala 33:21]
    matrix_7_2 <= matrix_7_2; // @[FlexDPE.scala 33:21]
    matrix_7_3 <= matrix_7_3; // @[FlexDPE.scala 33:21]
    matrix_7_4 <= matrix_7_4; // @[FlexDPE.scala 33:21]
    matrix_7_5 <= matrix_7_5; // @[FlexDPE.scala 33:21]
    matrix_7_6 <= matrix_7_6; // @[FlexDPE.scala 33:21]
    matrix_7_7 <= matrix_7_7; // @[FlexDPE.scala 33:21]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_mult_0 = _RAND_0[14:0];
  _RAND_1 = {1{`RANDOM}};
  r_mult_1 = _RAND_1[14:0];
  _RAND_2 = {1{`RANDOM}};
  r_mult_2 = _RAND_2[14:0];
  _RAND_3 = {1{`RANDOM}};
  r_mult_3 = _RAND_3[14:0];
  _RAND_4 = {1{`RANDOM}};
  matrix_0_0 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  matrix_0_1 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  matrix_0_2 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  matrix_0_3 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  matrix_0_4 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  matrix_0_5 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  matrix_0_6 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  matrix_0_7 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  matrix_1_0 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  matrix_1_1 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  matrix_1_2 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  matrix_1_3 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  matrix_1_4 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  matrix_1_5 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  matrix_1_6 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  matrix_1_7 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  matrix_2_0 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  matrix_2_1 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  matrix_2_2 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  matrix_2_3 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  matrix_2_4 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  matrix_2_5 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  matrix_2_6 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  matrix_2_7 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  matrix_3_0 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  matrix_3_1 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  matrix_3_2 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  matrix_3_3 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  matrix_3_4 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  matrix_3_5 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  matrix_3_6 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  matrix_3_7 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  matrix_4_0 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  matrix_4_1 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  matrix_4_2 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  matrix_4_3 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  matrix_4_4 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  matrix_4_5 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  matrix_4_6 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  matrix_4_7 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  matrix_5_0 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  matrix_5_1 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  matrix_5_2 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  matrix_5_3 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  matrix_5_4 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  matrix_5_5 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  matrix_5_6 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  matrix_5_7 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  matrix_6_0 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  matrix_6_1 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  matrix_6_2 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  matrix_6_3 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  matrix_6_4 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  matrix_6_5 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  matrix_6_6 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  matrix_6_7 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  matrix_7_0 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  matrix_7_1 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  matrix_7_2 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  matrix_7_3 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  matrix_7_4 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  matrix_7_5 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  matrix_7_6 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  matrix_7_7 = _RAND_67[15:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FlexDPU(
  input         clock,
  input         reset,
  input  [15:0] io_Stationary_matrix_0_0,
  input  [15:0] io_Stationary_matrix_0_1,
  input  [15:0] io_Stationary_matrix_0_2,
  input  [15:0] io_Stationary_matrix_0_3,
  input  [15:0] io_Stationary_matrix_0_4,
  input  [15:0] io_Stationary_matrix_0_5,
  input  [15:0] io_Stationary_matrix_0_6,
  input  [15:0] io_Stationary_matrix_0_7,
  input  [15:0] io_Stationary_matrix_1_0,
  input  [15:0] io_Stationary_matrix_1_1,
  input  [15:0] io_Stationary_matrix_1_2,
  input  [15:0] io_Stationary_matrix_1_3,
  input  [15:0] io_Stationary_matrix_1_4,
  input  [15:0] io_Stationary_matrix_1_5,
  input  [15:0] io_Stationary_matrix_1_6,
  input  [15:0] io_Stationary_matrix_1_7,
  input  [15:0] io_Stationary_matrix_2_0,
  input  [15:0] io_Stationary_matrix_2_1,
  input  [15:0] io_Stationary_matrix_2_2,
  input  [15:0] io_Stationary_matrix_2_3,
  input  [15:0] io_Stationary_matrix_2_4,
  input  [15:0] io_Stationary_matrix_2_5,
  input  [15:0] io_Stationary_matrix_2_6,
  input  [15:0] io_Stationary_matrix_2_7,
  input  [15:0] io_Stationary_matrix_3_0,
  input  [15:0] io_Stationary_matrix_3_1,
  input  [15:0] io_Stationary_matrix_3_2,
  input  [15:0] io_Stationary_matrix_3_3,
  input  [15:0] io_Stationary_matrix_3_4,
  input  [15:0] io_Stationary_matrix_3_5,
  input  [15:0] io_Stationary_matrix_3_6,
  input  [15:0] io_Stationary_matrix_3_7,
  input  [15:0] io_Stationary_matrix_4_0,
  input  [15:0] io_Stationary_matrix_4_1,
  input  [15:0] io_Stationary_matrix_4_2,
  input  [15:0] io_Stationary_matrix_4_3,
  input  [15:0] io_Stationary_matrix_4_4,
  input  [15:0] io_Stationary_matrix_4_5,
  input  [15:0] io_Stationary_matrix_4_6,
  input  [15:0] io_Stationary_matrix_4_7,
  input  [15:0] io_Stationary_matrix_5_0,
  input  [15:0] io_Stationary_matrix_5_1,
  input  [15:0] io_Stationary_matrix_5_2,
  input  [15:0] io_Stationary_matrix_5_3,
  input  [15:0] io_Stationary_matrix_5_4,
  input  [15:0] io_Stationary_matrix_5_5,
  input  [15:0] io_Stationary_matrix_5_6,
  input  [15:0] io_Stationary_matrix_5_7,
  input  [15:0] io_Stationary_matrix_6_0,
  input  [15:0] io_Stationary_matrix_6_1,
  input  [15:0] io_Stationary_matrix_6_2,
  input  [15:0] io_Stationary_matrix_6_3,
  input  [15:0] io_Stationary_matrix_6_4,
  input  [15:0] io_Stationary_matrix_6_5,
  input  [15:0] io_Stationary_matrix_6_6,
  input  [15:0] io_Stationary_matrix_6_7,
  input  [15:0] io_Stationary_matrix_7_0,
  input  [15:0] io_Stationary_matrix_7_1,
  input  [15:0] io_Stationary_matrix_7_2,
  input  [15:0] io_Stationary_matrix_7_3,
  input  [15:0] io_Stationary_matrix_7_4,
  input  [15:0] io_Stationary_matrix_7_5,
  input  [15:0] io_Stationary_matrix_7_6,
  input  [15:0] io_Stationary_matrix_7_7,
  input  [15:0] io_Streaming_matrix_0_0,
  input  [15:0] io_Streaming_matrix_0_1,
  input  [15:0] io_Streaming_matrix_0_2,
  input  [15:0] io_Streaming_matrix_0_3,
  input  [15:0] io_Streaming_matrix_0_4,
  input  [15:0] io_Streaming_matrix_0_5,
  input  [15:0] io_Streaming_matrix_0_6,
  input  [15:0] io_Streaming_matrix_0_7,
  input  [15:0] io_Streaming_matrix_1_0,
  input  [15:0] io_Streaming_matrix_1_1,
  input  [15:0] io_Streaming_matrix_1_2,
  input  [15:0] io_Streaming_matrix_1_3,
  input  [15:0] io_Streaming_matrix_1_4,
  input  [15:0] io_Streaming_matrix_1_5,
  input  [15:0] io_Streaming_matrix_1_6,
  input  [15:0] io_Streaming_matrix_1_7,
  input  [15:0] io_Streaming_matrix_2_0,
  input  [15:0] io_Streaming_matrix_2_1,
  input  [15:0] io_Streaming_matrix_2_2,
  input  [15:0] io_Streaming_matrix_2_3,
  input  [15:0] io_Streaming_matrix_2_4,
  input  [15:0] io_Streaming_matrix_2_5,
  input  [15:0] io_Streaming_matrix_2_6,
  input  [15:0] io_Streaming_matrix_2_7,
  input  [15:0] io_Streaming_matrix_3_0,
  input  [15:0] io_Streaming_matrix_3_1,
  input  [15:0] io_Streaming_matrix_3_2,
  input  [15:0] io_Streaming_matrix_3_3,
  input  [15:0] io_Streaming_matrix_3_4,
  input  [15:0] io_Streaming_matrix_3_5,
  input  [15:0] io_Streaming_matrix_3_6,
  input  [15:0] io_Streaming_matrix_3_7,
  input  [15:0] io_Streaming_matrix_4_0,
  input  [15:0] io_Streaming_matrix_4_1,
  input  [15:0] io_Streaming_matrix_4_2,
  input  [15:0] io_Streaming_matrix_4_3,
  input  [15:0] io_Streaming_matrix_4_4,
  input  [15:0] io_Streaming_matrix_4_5,
  input  [15:0] io_Streaming_matrix_4_6,
  input  [15:0] io_Streaming_matrix_4_7,
  input  [15:0] io_Streaming_matrix_5_0,
  input  [15:0] io_Streaming_matrix_5_1,
  input  [15:0] io_Streaming_matrix_5_2,
  input  [15:0] io_Streaming_matrix_5_3,
  input  [15:0] io_Streaming_matrix_5_4,
  input  [15:0] io_Streaming_matrix_5_5,
  input  [15:0] io_Streaming_matrix_5_6,
  input  [15:0] io_Streaming_matrix_5_7,
  input  [15:0] io_Streaming_matrix_6_0,
  input  [15:0] io_Streaming_matrix_6_1,
  input  [15:0] io_Streaming_matrix_6_2,
  input  [15:0] io_Streaming_matrix_6_3,
  input  [15:0] io_Streaming_matrix_6_4,
  input  [15:0] io_Streaming_matrix_6_5,
  input  [15:0] io_Streaming_matrix_6_6,
  input  [15:0] io_Streaming_matrix_6_7,
  input  [15:0] io_Streaming_matrix_7_0,
  input  [15:0] io_Streaming_matrix_7_1,
  input  [15:0] io_Streaming_matrix_7_2,
  input  [15:0] io_Streaming_matrix_7_3,
  input  [15:0] io_Streaming_matrix_7_4,
  input  [15:0] io_Streaming_matrix_7_5,
  input  [15:0] io_Streaming_matrix_7_6,
  input  [15:0] io_Streaming_matrix_7_7
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
`endif // RANDOMIZE_REG_INIT
  wire  PathFinder_clock; // @[FlexDPU.scala 77:41]
  wire  PathFinder_reset; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_0_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_0_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_0_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_0_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_0_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_0_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_0_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_0_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_1_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_1_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_1_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_1_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_1_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_1_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_1_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_1_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_2_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_2_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_2_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_2_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_2_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_2_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_2_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_2_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_3_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_3_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_3_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_3_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_3_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_3_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_3_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_3_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_4_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_4_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_4_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_4_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_4_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_4_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_4_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_4_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_5_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_5_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_5_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_5_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_5_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_5_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_5_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_5_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_6_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_6_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_6_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_6_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_6_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_6_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_6_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_6_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_7_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_7_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_7_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_7_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_7_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_7_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_7_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Stationary_matrix_7_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Streaming_matrix_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Streaming_matrix_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Streaming_matrix_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Streaming_matrix_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Streaming_matrix_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Streaming_matrix_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Streaming_matrix_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Streaming_matrix_7; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_io_i_mux_bus_0; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_io_i_mux_bus_1; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_io_i_mux_bus_2; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_io_i_mux_bus_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Source_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Source_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Source_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_io_Source_3; // @[FlexDPU.scala 77:41]
  wire  PathFinder_io_PF_Valid; // @[FlexDPU.scala 77:41]
  wire [31:0] PathFinder_io_NoDPE; // @[FlexDPU.scala 77:41]
  wire  PathFinder_io_DataValid; // @[FlexDPU.scala 77:41]
  wire  PathFinder_1_clock; // @[FlexDPU.scala 77:41]
  wire  PathFinder_1_reset; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_0_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_0_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_0_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_0_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_0_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_0_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_0_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_0_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_1_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_1_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_1_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_1_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_1_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_1_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_1_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_1_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_2_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_2_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_2_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_2_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_2_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_2_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_2_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_2_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_3_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_3_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_3_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_3_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_3_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_3_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_3_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_3_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_4_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_4_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_4_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_4_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_4_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_4_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_4_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_4_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_5_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_5_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_5_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_5_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_5_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_5_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_5_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_5_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_6_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_6_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_6_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_6_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_6_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_6_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_6_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_6_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_7_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_7_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_7_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_7_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_7_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_7_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_7_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Stationary_matrix_7_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Streaming_matrix_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Streaming_matrix_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Streaming_matrix_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Streaming_matrix_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Streaming_matrix_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Streaming_matrix_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Streaming_matrix_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Streaming_matrix_7; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_1_io_i_mux_bus_0; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_1_io_i_mux_bus_1; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_1_io_i_mux_bus_2; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_1_io_i_mux_bus_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Source_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Source_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Source_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_1_io_Source_3; // @[FlexDPU.scala 77:41]
  wire  PathFinder_1_io_PF_Valid; // @[FlexDPU.scala 77:41]
  wire [31:0] PathFinder_1_io_NoDPE; // @[FlexDPU.scala 77:41]
  wire  PathFinder_1_io_DataValid; // @[FlexDPU.scala 77:41]
  wire  PathFinder_2_clock; // @[FlexDPU.scala 77:41]
  wire  PathFinder_2_reset; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_0_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_0_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_0_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_0_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_0_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_0_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_0_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_0_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_1_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_1_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_1_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_1_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_1_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_1_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_1_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_1_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_2_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_2_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_2_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_2_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_2_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_2_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_2_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_2_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_3_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_3_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_3_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_3_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_3_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_3_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_3_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_3_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_4_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_4_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_4_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_4_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_4_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_4_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_4_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_4_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_5_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_5_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_5_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_5_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_5_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_5_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_5_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_5_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_6_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_6_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_6_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_6_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_6_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_6_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_6_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_6_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_7_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_7_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_7_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_7_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_7_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_7_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_7_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Stationary_matrix_7_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Streaming_matrix_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Streaming_matrix_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Streaming_matrix_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Streaming_matrix_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Streaming_matrix_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Streaming_matrix_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Streaming_matrix_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Streaming_matrix_7; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_2_io_i_mux_bus_0; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_2_io_i_mux_bus_1; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_2_io_i_mux_bus_2; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_2_io_i_mux_bus_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Source_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Source_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Source_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_2_io_Source_3; // @[FlexDPU.scala 77:41]
  wire  PathFinder_2_io_PF_Valid; // @[FlexDPU.scala 77:41]
  wire [31:0] PathFinder_2_io_NoDPE; // @[FlexDPU.scala 77:41]
  wire  PathFinder_2_io_DataValid; // @[FlexDPU.scala 77:41]
  wire  PathFinder_3_clock; // @[FlexDPU.scala 77:41]
  wire  PathFinder_3_reset; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_0_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_0_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_0_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_0_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_0_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_0_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_0_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_0_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_1_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_1_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_1_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_1_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_1_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_1_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_1_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_1_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_2_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_2_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_2_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_2_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_2_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_2_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_2_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_2_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_3_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_3_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_3_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_3_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_3_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_3_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_3_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_3_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_4_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_4_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_4_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_4_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_4_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_4_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_4_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_4_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_5_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_5_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_5_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_5_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_5_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_5_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_5_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_5_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_6_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_6_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_6_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_6_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_6_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_6_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_6_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_6_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_7_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_7_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_7_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_7_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_7_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_7_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_7_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Stationary_matrix_7_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Streaming_matrix_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Streaming_matrix_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Streaming_matrix_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Streaming_matrix_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Streaming_matrix_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Streaming_matrix_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Streaming_matrix_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Streaming_matrix_7; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_3_io_i_mux_bus_0; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_3_io_i_mux_bus_1; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_3_io_i_mux_bus_2; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_3_io_i_mux_bus_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Source_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Source_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Source_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_3_io_Source_3; // @[FlexDPU.scala 77:41]
  wire  PathFinder_3_io_PF_Valid; // @[FlexDPU.scala 77:41]
  wire [31:0] PathFinder_3_io_NoDPE; // @[FlexDPU.scala 77:41]
  wire  PathFinder_3_io_DataValid; // @[FlexDPU.scala 77:41]
  wire  PathFinder_4_clock; // @[FlexDPU.scala 77:41]
  wire  PathFinder_4_reset; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_0_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_0_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_0_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_0_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_0_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_0_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_0_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_0_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_1_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_1_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_1_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_1_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_1_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_1_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_1_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_1_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_2_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_2_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_2_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_2_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_2_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_2_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_2_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_2_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_3_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_3_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_3_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_3_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_3_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_3_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_3_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_3_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_4_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_4_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_4_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_4_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_4_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_4_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_4_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_4_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_5_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_5_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_5_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_5_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_5_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_5_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_5_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_5_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_6_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_6_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_6_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_6_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_6_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_6_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_6_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_6_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_7_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_7_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_7_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_7_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_7_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_7_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_7_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Stationary_matrix_7_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Streaming_matrix_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Streaming_matrix_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Streaming_matrix_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Streaming_matrix_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Streaming_matrix_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Streaming_matrix_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Streaming_matrix_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Streaming_matrix_7; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_4_io_i_mux_bus_0; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_4_io_i_mux_bus_1; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_4_io_i_mux_bus_2; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_4_io_i_mux_bus_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Source_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Source_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Source_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_4_io_Source_3; // @[FlexDPU.scala 77:41]
  wire  PathFinder_4_io_PF_Valid; // @[FlexDPU.scala 77:41]
  wire [31:0] PathFinder_4_io_NoDPE; // @[FlexDPU.scala 77:41]
  wire  PathFinder_4_io_DataValid; // @[FlexDPU.scala 77:41]
  wire  PathFinder_5_clock; // @[FlexDPU.scala 77:41]
  wire  PathFinder_5_reset; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_0_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_0_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_0_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_0_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_0_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_0_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_0_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_0_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_1_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_1_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_1_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_1_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_1_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_1_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_1_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_1_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_2_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_2_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_2_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_2_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_2_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_2_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_2_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_2_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_3_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_3_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_3_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_3_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_3_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_3_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_3_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_3_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_4_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_4_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_4_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_4_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_4_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_4_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_4_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_4_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_5_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_5_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_5_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_5_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_5_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_5_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_5_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_5_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_6_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_6_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_6_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_6_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_6_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_6_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_6_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_6_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_7_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_7_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_7_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_7_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_7_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_7_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_7_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Stationary_matrix_7_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Streaming_matrix_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Streaming_matrix_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Streaming_matrix_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Streaming_matrix_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Streaming_matrix_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Streaming_matrix_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Streaming_matrix_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Streaming_matrix_7; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_5_io_i_mux_bus_0; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_5_io_i_mux_bus_1; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_5_io_i_mux_bus_2; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_5_io_i_mux_bus_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Source_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Source_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Source_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_5_io_Source_3; // @[FlexDPU.scala 77:41]
  wire  PathFinder_5_io_PF_Valid; // @[FlexDPU.scala 77:41]
  wire [31:0] PathFinder_5_io_NoDPE; // @[FlexDPU.scala 77:41]
  wire  PathFinder_5_io_DataValid; // @[FlexDPU.scala 77:41]
  wire  PathFinder_6_clock; // @[FlexDPU.scala 77:41]
  wire  PathFinder_6_reset; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_0_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_0_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_0_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_0_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_0_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_0_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_0_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_0_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_1_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_1_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_1_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_1_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_1_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_1_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_1_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_1_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_2_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_2_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_2_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_2_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_2_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_2_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_2_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_2_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_3_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_3_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_3_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_3_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_3_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_3_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_3_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_3_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_4_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_4_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_4_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_4_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_4_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_4_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_4_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_4_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_5_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_5_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_5_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_5_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_5_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_5_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_5_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_5_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_6_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_6_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_6_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_6_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_6_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_6_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_6_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_6_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_7_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_7_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_7_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_7_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_7_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_7_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_7_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Stationary_matrix_7_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Streaming_matrix_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Streaming_matrix_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Streaming_matrix_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Streaming_matrix_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Streaming_matrix_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Streaming_matrix_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Streaming_matrix_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Streaming_matrix_7; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_6_io_i_mux_bus_0; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_6_io_i_mux_bus_1; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_6_io_i_mux_bus_2; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_6_io_i_mux_bus_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Source_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Source_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Source_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_6_io_Source_3; // @[FlexDPU.scala 77:41]
  wire  PathFinder_6_io_PF_Valid; // @[FlexDPU.scala 77:41]
  wire [31:0] PathFinder_6_io_NoDPE; // @[FlexDPU.scala 77:41]
  wire  PathFinder_6_io_DataValid; // @[FlexDPU.scala 77:41]
  wire  PathFinder_7_clock; // @[FlexDPU.scala 77:41]
  wire  PathFinder_7_reset; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_0_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_0_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_0_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_0_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_0_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_0_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_0_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_0_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_1_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_1_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_1_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_1_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_1_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_1_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_1_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_1_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_2_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_2_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_2_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_2_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_2_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_2_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_2_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_2_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_3_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_3_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_3_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_3_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_3_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_3_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_3_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_3_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_4_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_4_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_4_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_4_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_4_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_4_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_4_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_4_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_5_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_5_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_5_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_5_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_5_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_5_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_5_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_5_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_6_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_6_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_6_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_6_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_6_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_6_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_6_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_6_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_7_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_7_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_7_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_7_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_7_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_7_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_7_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Stationary_matrix_7_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Streaming_matrix_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Streaming_matrix_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Streaming_matrix_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Streaming_matrix_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Streaming_matrix_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Streaming_matrix_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Streaming_matrix_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Streaming_matrix_7; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_7_io_i_mux_bus_0; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_7_io_i_mux_bus_1; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_7_io_i_mux_bus_2; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_7_io_i_mux_bus_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Source_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Source_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Source_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_7_io_Source_3; // @[FlexDPU.scala 77:41]
  wire  PathFinder_7_io_PF_Valid; // @[FlexDPU.scala 77:41]
  wire [31:0] PathFinder_7_io_NoDPE; // @[FlexDPU.scala 77:41]
  wire  PathFinder_7_io_DataValid; // @[FlexDPU.scala 77:41]
  wire  PathFinder_8_clock; // @[FlexDPU.scala 77:41]
  wire  PathFinder_8_reset; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_0_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_0_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_0_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_0_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_0_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_0_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_0_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_0_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_1_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_1_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_1_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_1_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_1_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_1_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_1_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_1_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_2_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_2_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_2_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_2_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_2_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_2_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_2_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_2_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_3_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_3_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_3_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_3_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_3_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_3_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_3_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_3_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_4_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_4_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_4_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_4_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_4_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_4_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_4_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_4_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_5_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_5_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_5_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_5_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_5_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_5_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_5_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_5_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_6_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_6_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_6_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_6_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_6_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_6_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_6_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_6_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_7_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_7_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_7_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_7_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_7_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_7_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_7_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Stationary_matrix_7_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Streaming_matrix_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Streaming_matrix_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Streaming_matrix_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Streaming_matrix_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Streaming_matrix_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Streaming_matrix_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Streaming_matrix_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Streaming_matrix_7; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_8_io_i_mux_bus_0; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_8_io_i_mux_bus_1; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_8_io_i_mux_bus_2; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_8_io_i_mux_bus_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Source_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Source_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Source_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_8_io_Source_3; // @[FlexDPU.scala 77:41]
  wire  PathFinder_8_io_PF_Valid; // @[FlexDPU.scala 77:41]
  wire [31:0] PathFinder_8_io_NoDPE; // @[FlexDPU.scala 77:41]
  wire  PathFinder_8_io_DataValid; // @[FlexDPU.scala 77:41]
  wire  PathFinder_9_clock; // @[FlexDPU.scala 77:41]
  wire  PathFinder_9_reset; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_0_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_0_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_0_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_0_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_0_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_0_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_0_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_0_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_1_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_1_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_1_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_1_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_1_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_1_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_1_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_1_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_2_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_2_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_2_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_2_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_2_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_2_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_2_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_2_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_3_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_3_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_3_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_3_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_3_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_3_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_3_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_3_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_4_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_4_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_4_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_4_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_4_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_4_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_4_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_4_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_5_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_5_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_5_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_5_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_5_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_5_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_5_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_5_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_6_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_6_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_6_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_6_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_6_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_6_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_6_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_6_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_7_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_7_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_7_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_7_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_7_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_7_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_7_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Stationary_matrix_7_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Streaming_matrix_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Streaming_matrix_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Streaming_matrix_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Streaming_matrix_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Streaming_matrix_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Streaming_matrix_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Streaming_matrix_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Streaming_matrix_7; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_9_io_i_mux_bus_0; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_9_io_i_mux_bus_1; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_9_io_i_mux_bus_2; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_9_io_i_mux_bus_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Source_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Source_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Source_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_9_io_Source_3; // @[FlexDPU.scala 77:41]
  wire  PathFinder_9_io_PF_Valid; // @[FlexDPU.scala 77:41]
  wire [31:0] PathFinder_9_io_NoDPE; // @[FlexDPU.scala 77:41]
  wire  PathFinder_9_io_DataValid; // @[FlexDPU.scala 77:41]
  wire  PathFinder_10_clock; // @[FlexDPU.scala 77:41]
  wire  PathFinder_10_reset; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_0_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_0_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_0_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_0_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_0_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_0_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_0_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_0_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_1_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_1_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_1_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_1_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_1_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_1_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_1_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_1_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_2_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_2_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_2_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_2_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_2_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_2_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_2_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_2_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_3_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_3_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_3_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_3_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_3_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_3_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_3_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_3_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_4_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_4_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_4_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_4_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_4_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_4_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_4_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_4_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_5_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_5_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_5_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_5_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_5_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_5_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_5_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_5_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_6_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_6_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_6_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_6_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_6_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_6_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_6_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_6_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_7_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_7_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_7_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_7_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_7_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_7_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_7_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Stationary_matrix_7_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Streaming_matrix_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Streaming_matrix_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Streaming_matrix_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Streaming_matrix_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Streaming_matrix_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Streaming_matrix_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Streaming_matrix_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Streaming_matrix_7; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_10_io_i_mux_bus_0; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_10_io_i_mux_bus_1; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_10_io_i_mux_bus_2; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_10_io_i_mux_bus_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Source_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Source_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Source_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_10_io_Source_3; // @[FlexDPU.scala 77:41]
  wire  PathFinder_10_io_PF_Valid; // @[FlexDPU.scala 77:41]
  wire [31:0] PathFinder_10_io_NoDPE; // @[FlexDPU.scala 77:41]
  wire  PathFinder_10_io_DataValid; // @[FlexDPU.scala 77:41]
  wire  PathFinder_11_clock; // @[FlexDPU.scala 77:41]
  wire  PathFinder_11_reset; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_0_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_0_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_0_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_0_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_0_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_0_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_0_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_0_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_1_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_1_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_1_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_1_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_1_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_1_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_1_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_1_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_2_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_2_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_2_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_2_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_2_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_2_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_2_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_2_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_3_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_3_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_3_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_3_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_3_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_3_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_3_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_3_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_4_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_4_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_4_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_4_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_4_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_4_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_4_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_4_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_5_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_5_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_5_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_5_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_5_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_5_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_5_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_5_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_6_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_6_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_6_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_6_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_6_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_6_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_6_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_6_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_7_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_7_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_7_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_7_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_7_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_7_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_7_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Stationary_matrix_7_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Streaming_matrix_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Streaming_matrix_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Streaming_matrix_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Streaming_matrix_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Streaming_matrix_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Streaming_matrix_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Streaming_matrix_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Streaming_matrix_7; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_11_io_i_mux_bus_0; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_11_io_i_mux_bus_1; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_11_io_i_mux_bus_2; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_11_io_i_mux_bus_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Source_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Source_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Source_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_11_io_Source_3; // @[FlexDPU.scala 77:41]
  wire  PathFinder_11_io_PF_Valid; // @[FlexDPU.scala 77:41]
  wire [31:0] PathFinder_11_io_NoDPE; // @[FlexDPU.scala 77:41]
  wire  PathFinder_11_io_DataValid; // @[FlexDPU.scala 77:41]
  wire  PathFinder_12_clock; // @[FlexDPU.scala 77:41]
  wire  PathFinder_12_reset; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_0_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_0_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_0_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_0_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_0_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_0_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_0_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_0_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_1_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_1_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_1_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_1_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_1_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_1_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_1_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_1_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_2_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_2_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_2_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_2_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_2_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_2_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_2_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_2_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_3_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_3_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_3_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_3_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_3_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_3_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_3_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_3_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_4_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_4_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_4_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_4_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_4_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_4_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_4_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_4_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_5_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_5_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_5_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_5_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_5_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_5_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_5_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_5_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_6_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_6_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_6_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_6_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_6_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_6_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_6_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_6_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_7_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_7_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_7_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_7_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_7_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_7_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_7_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Stationary_matrix_7_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Streaming_matrix_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Streaming_matrix_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Streaming_matrix_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Streaming_matrix_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Streaming_matrix_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Streaming_matrix_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Streaming_matrix_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Streaming_matrix_7; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_12_io_i_mux_bus_0; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_12_io_i_mux_bus_1; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_12_io_i_mux_bus_2; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_12_io_i_mux_bus_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Source_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Source_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Source_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_12_io_Source_3; // @[FlexDPU.scala 77:41]
  wire  PathFinder_12_io_PF_Valid; // @[FlexDPU.scala 77:41]
  wire [31:0] PathFinder_12_io_NoDPE; // @[FlexDPU.scala 77:41]
  wire  PathFinder_12_io_DataValid; // @[FlexDPU.scala 77:41]
  wire  PathFinder_13_clock; // @[FlexDPU.scala 77:41]
  wire  PathFinder_13_reset; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_0_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_0_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_0_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_0_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_0_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_0_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_0_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_0_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_1_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_1_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_1_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_1_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_1_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_1_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_1_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_1_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_2_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_2_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_2_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_2_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_2_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_2_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_2_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_2_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_3_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_3_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_3_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_3_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_3_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_3_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_3_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_3_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_4_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_4_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_4_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_4_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_4_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_4_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_4_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_4_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_5_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_5_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_5_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_5_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_5_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_5_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_5_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_5_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_6_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_6_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_6_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_6_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_6_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_6_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_6_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_6_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_7_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_7_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_7_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_7_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_7_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_7_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_7_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Stationary_matrix_7_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Streaming_matrix_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Streaming_matrix_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Streaming_matrix_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Streaming_matrix_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Streaming_matrix_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Streaming_matrix_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Streaming_matrix_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Streaming_matrix_7; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_13_io_i_mux_bus_0; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_13_io_i_mux_bus_1; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_13_io_i_mux_bus_2; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_13_io_i_mux_bus_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Source_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Source_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Source_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_13_io_Source_3; // @[FlexDPU.scala 77:41]
  wire  PathFinder_13_io_PF_Valid; // @[FlexDPU.scala 77:41]
  wire [31:0] PathFinder_13_io_NoDPE; // @[FlexDPU.scala 77:41]
  wire  PathFinder_13_io_DataValid; // @[FlexDPU.scala 77:41]
  wire  PathFinder_14_clock; // @[FlexDPU.scala 77:41]
  wire  PathFinder_14_reset; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_0_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_0_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_0_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_0_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_0_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_0_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_0_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_0_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_1_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_1_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_1_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_1_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_1_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_1_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_1_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_1_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_2_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_2_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_2_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_2_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_2_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_2_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_2_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_2_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_3_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_3_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_3_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_3_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_3_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_3_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_3_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_3_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_4_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_4_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_4_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_4_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_4_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_4_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_4_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_4_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_5_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_5_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_5_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_5_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_5_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_5_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_5_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_5_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_6_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_6_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_6_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_6_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_6_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_6_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_6_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_6_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_7_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_7_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_7_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_7_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_7_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_7_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_7_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Stationary_matrix_7_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Streaming_matrix_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Streaming_matrix_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Streaming_matrix_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Streaming_matrix_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Streaming_matrix_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Streaming_matrix_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Streaming_matrix_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Streaming_matrix_7; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_14_io_i_mux_bus_0; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_14_io_i_mux_bus_1; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_14_io_i_mux_bus_2; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_14_io_i_mux_bus_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Source_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Source_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Source_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_14_io_Source_3; // @[FlexDPU.scala 77:41]
  wire  PathFinder_14_io_PF_Valid; // @[FlexDPU.scala 77:41]
  wire [31:0] PathFinder_14_io_NoDPE; // @[FlexDPU.scala 77:41]
  wire  PathFinder_14_io_DataValid; // @[FlexDPU.scala 77:41]
  wire  PathFinder_15_clock; // @[FlexDPU.scala 77:41]
  wire  PathFinder_15_reset; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_0_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_0_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_0_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_0_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_0_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_0_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_0_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_0_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_1_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_1_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_1_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_1_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_1_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_1_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_1_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_1_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_2_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_2_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_2_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_2_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_2_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_2_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_2_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_2_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_3_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_3_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_3_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_3_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_3_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_3_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_3_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_3_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_4_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_4_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_4_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_4_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_4_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_4_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_4_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_4_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_5_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_5_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_5_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_5_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_5_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_5_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_5_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_5_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_6_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_6_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_6_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_6_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_6_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_6_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_6_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_6_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_7_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_7_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_7_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_7_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_7_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_7_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_7_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Stationary_matrix_7_7; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Streaming_matrix_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Streaming_matrix_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Streaming_matrix_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Streaming_matrix_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Streaming_matrix_4; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Streaming_matrix_5; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Streaming_matrix_6; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Streaming_matrix_7; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_15_io_i_mux_bus_0; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_15_io_i_mux_bus_1; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_15_io_i_mux_bus_2; // @[FlexDPU.scala 77:41]
  wire [3:0] PathFinder_15_io_i_mux_bus_3; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Source_0; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Source_1; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Source_2; // @[FlexDPU.scala 77:41]
  wire [15:0] PathFinder_15_io_Source_3; // @[FlexDPU.scala 77:41]
  wire  PathFinder_15_io_PF_Valid; // @[FlexDPU.scala 77:41]
  wire [31:0] PathFinder_15_io_NoDPE; // @[FlexDPU.scala 77:41]
  wire  PathFinder_15_io_DataValid; // @[FlexDPU.scala 77:41]
  wire  ivntop_clock; // @[FlexDPU.scala 87:21]
  wire  ivntop_reset; // @[FlexDPU.scala 87:21]
  wire  ivntop_io_ProcessValid; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_0_0; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_0_1; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_0_2; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_0_3; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_0_4; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_0_5; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_0_6; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_0_7; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_1_0; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_1_1; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_1_2; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_1_3; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_1_4; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_1_5; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_1_6; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_1_7; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_2_0; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_2_1; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_2_2; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_2_3; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_2_4; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_2_5; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_2_6; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_2_7; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_3_0; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_3_1; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_3_2; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_3_3; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_3_4; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_3_5; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_3_6; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_3_7; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_4_0; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_4_1; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_4_2; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_4_3; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_4_4; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_4_5; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_4_6; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_4_7; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_5_0; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_5_1; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_5_2; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_5_3; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_5_4; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_5_5; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_5_6; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_5_7; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_6_0; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_6_1; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_6_2; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_6_3; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_6_4; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_6_5; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_6_6; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_6_7; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_7_0; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_7_1; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_7_2; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_7_3; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_7_4; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_7_5; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_7_6; // @[FlexDPU.scala 87:21]
  wire [15:0] ivntop_io_Stationary_matrix_7_7; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_0_0; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_0_1; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_0_2; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_0_3; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_1_0; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_1_1; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_1_2; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_1_3; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_2_0; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_2_1; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_2_2; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_2_3; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_3_0; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_3_1; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_3_2; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_3_3; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_4_0; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_4_1; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_4_2; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_4_3; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_5_0; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_5_1; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_5_2; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_5_3; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_6_0; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_6_1; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_6_2; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_6_3; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_7_0; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_7_1; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_7_2; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_7_3; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_8_0; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_8_1; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_8_2; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_8_3; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_9_0; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_9_1; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_9_2; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_9_3; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_10_0; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_10_1; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_10_2; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_10_3; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_11_0; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_11_1; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_11_2; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_11_3; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_12_0; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_12_1; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_12_2; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_12_3; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_13_0; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_13_1; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_13_2; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_13_3; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_14_0; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_14_1; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_14_2; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_14_3; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_15_0; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_15_1; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_15_2; // @[FlexDPU.scala 87:21]
  wire [4:0] ivntop_io_o_vn_15_3; // @[FlexDPU.scala 87:21]
  wire  MuxesWrapper_io_valid; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_io_src_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_io_src_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_io_src_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_io_src_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_io_muxes_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_io_muxes_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_io_muxes_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_io_muxes_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_io_Osrc_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_io_Osrc_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_io_Osrc_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_io_Osrc_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_io_Omuxes_0_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_io_Omuxes_0_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_io_Omuxes_0_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_io_Omuxes_0_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_io_Omuxes_1_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_io_Omuxes_1_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_io_Omuxes_1_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_io_Omuxes_2_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_io_Omuxes_2_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_io_Omuxes_3_0; // @[FlexDPU.scala 124:53]
  wire  MuxesWrapper_1_io_valid; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_1_io_src_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_1_io_src_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_1_io_src_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_1_io_src_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_1_io_muxes_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_1_io_muxes_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_1_io_muxes_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_1_io_muxes_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_1_io_Osrc_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_1_io_Osrc_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_1_io_Osrc_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_1_io_Osrc_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_1_io_Omuxes_0_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_1_io_Omuxes_0_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_1_io_Omuxes_0_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_1_io_Omuxes_0_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_1_io_Omuxes_1_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_1_io_Omuxes_1_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_1_io_Omuxes_1_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_1_io_Omuxes_2_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_1_io_Omuxes_2_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_1_io_Omuxes_3_0; // @[FlexDPU.scala 124:53]
  wire  MuxesWrapper_2_io_valid; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_2_io_src_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_2_io_src_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_2_io_src_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_2_io_src_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_2_io_muxes_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_2_io_muxes_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_2_io_muxes_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_2_io_muxes_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_2_io_Osrc_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_2_io_Osrc_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_2_io_Osrc_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_2_io_Osrc_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_2_io_Omuxes_0_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_2_io_Omuxes_0_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_2_io_Omuxes_0_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_2_io_Omuxes_0_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_2_io_Omuxes_1_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_2_io_Omuxes_1_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_2_io_Omuxes_1_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_2_io_Omuxes_2_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_2_io_Omuxes_2_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_2_io_Omuxes_3_0; // @[FlexDPU.scala 124:53]
  wire  MuxesWrapper_3_io_valid; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_3_io_src_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_3_io_src_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_3_io_src_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_3_io_src_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_3_io_muxes_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_3_io_muxes_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_3_io_muxes_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_3_io_muxes_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_3_io_Osrc_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_3_io_Osrc_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_3_io_Osrc_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_3_io_Osrc_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_3_io_Omuxes_0_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_3_io_Omuxes_0_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_3_io_Omuxes_0_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_3_io_Omuxes_0_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_3_io_Omuxes_1_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_3_io_Omuxes_1_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_3_io_Omuxes_1_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_3_io_Omuxes_2_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_3_io_Omuxes_2_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_3_io_Omuxes_3_0; // @[FlexDPU.scala 124:53]
  wire  MuxesWrapper_4_io_valid; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_4_io_src_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_4_io_src_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_4_io_src_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_4_io_src_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_4_io_muxes_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_4_io_muxes_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_4_io_muxes_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_4_io_muxes_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_4_io_Osrc_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_4_io_Osrc_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_4_io_Osrc_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_4_io_Osrc_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_4_io_Omuxes_0_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_4_io_Omuxes_0_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_4_io_Omuxes_0_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_4_io_Omuxes_0_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_4_io_Omuxes_1_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_4_io_Omuxes_1_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_4_io_Omuxes_1_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_4_io_Omuxes_2_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_4_io_Omuxes_2_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_4_io_Omuxes_3_0; // @[FlexDPU.scala 124:53]
  wire  MuxesWrapper_5_io_valid; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_5_io_src_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_5_io_src_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_5_io_src_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_5_io_src_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_5_io_muxes_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_5_io_muxes_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_5_io_muxes_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_5_io_muxes_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_5_io_Osrc_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_5_io_Osrc_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_5_io_Osrc_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_5_io_Osrc_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_5_io_Omuxes_0_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_5_io_Omuxes_0_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_5_io_Omuxes_0_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_5_io_Omuxes_0_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_5_io_Omuxes_1_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_5_io_Omuxes_1_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_5_io_Omuxes_1_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_5_io_Omuxes_2_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_5_io_Omuxes_2_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_5_io_Omuxes_3_0; // @[FlexDPU.scala 124:53]
  wire  MuxesWrapper_6_io_valid; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_6_io_src_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_6_io_src_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_6_io_src_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_6_io_src_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_6_io_muxes_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_6_io_muxes_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_6_io_muxes_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_6_io_muxes_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_6_io_Osrc_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_6_io_Osrc_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_6_io_Osrc_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_6_io_Osrc_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_6_io_Omuxes_0_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_6_io_Omuxes_0_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_6_io_Omuxes_0_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_6_io_Omuxes_0_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_6_io_Omuxes_1_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_6_io_Omuxes_1_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_6_io_Omuxes_1_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_6_io_Omuxes_2_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_6_io_Omuxes_2_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_6_io_Omuxes_3_0; // @[FlexDPU.scala 124:53]
  wire  MuxesWrapper_7_io_valid; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_7_io_src_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_7_io_src_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_7_io_src_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_7_io_src_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_7_io_muxes_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_7_io_muxes_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_7_io_muxes_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_7_io_muxes_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_7_io_Osrc_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_7_io_Osrc_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_7_io_Osrc_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_7_io_Osrc_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_7_io_Omuxes_0_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_7_io_Omuxes_0_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_7_io_Omuxes_0_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_7_io_Omuxes_0_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_7_io_Omuxes_1_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_7_io_Omuxes_1_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_7_io_Omuxes_1_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_7_io_Omuxes_2_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_7_io_Omuxes_2_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_7_io_Omuxes_3_0; // @[FlexDPU.scala 124:53]
  wire  MuxesWrapper_8_io_valid; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_8_io_src_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_8_io_src_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_8_io_src_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_8_io_src_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_8_io_muxes_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_8_io_muxes_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_8_io_muxes_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_8_io_muxes_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_8_io_Osrc_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_8_io_Osrc_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_8_io_Osrc_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_8_io_Osrc_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_8_io_Omuxes_0_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_8_io_Omuxes_0_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_8_io_Omuxes_0_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_8_io_Omuxes_0_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_8_io_Omuxes_1_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_8_io_Omuxes_1_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_8_io_Omuxes_1_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_8_io_Omuxes_2_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_8_io_Omuxes_2_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_8_io_Omuxes_3_0; // @[FlexDPU.scala 124:53]
  wire  MuxesWrapper_9_io_valid; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_9_io_src_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_9_io_src_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_9_io_src_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_9_io_src_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_9_io_muxes_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_9_io_muxes_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_9_io_muxes_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_9_io_muxes_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_9_io_Osrc_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_9_io_Osrc_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_9_io_Osrc_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_9_io_Osrc_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_9_io_Omuxes_0_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_9_io_Omuxes_0_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_9_io_Omuxes_0_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_9_io_Omuxes_0_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_9_io_Omuxes_1_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_9_io_Omuxes_1_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_9_io_Omuxes_1_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_9_io_Omuxes_2_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_9_io_Omuxes_2_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_9_io_Omuxes_3_0; // @[FlexDPU.scala 124:53]
  wire  MuxesWrapper_10_io_valid; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_10_io_src_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_10_io_src_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_10_io_src_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_10_io_src_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_10_io_muxes_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_10_io_muxes_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_10_io_muxes_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_10_io_muxes_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_10_io_Osrc_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_10_io_Osrc_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_10_io_Osrc_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_10_io_Osrc_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_10_io_Omuxes_0_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_10_io_Omuxes_0_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_10_io_Omuxes_0_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_10_io_Omuxes_0_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_10_io_Omuxes_1_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_10_io_Omuxes_1_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_10_io_Omuxes_1_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_10_io_Omuxes_2_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_10_io_Omuxes_2_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_10_io_Omuxes_3_0; // @[FlexDPU.scala 124:53]
  wire  MuxesWrapper_11_io_valid; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_11_io_src_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_11_io_src_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_11_io_src_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_11_io_src_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_11_io_muxes_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_11_io_muxes_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_11_io_muxes_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_11_io_muxes_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_11_io_Osrc_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_11_io_Osrc_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_11_io_Osrc_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_11_io_Osrc_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_11_io_Omuxes_0_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_11_io_Omuxes_0_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_11_io_Omuxes_0_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_11_io_Omuxes_0_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_11_io_Omuxes_1_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_11_io_Omuxes_1_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_11_io_Omuxes_1_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_11_io_Omuxes_2_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_11_io_Omuxes_2_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_11_io_Omuxes_3_0; // @[FlexDPU.scala 124:53]
  wire  MuxesWrapper_12_io_valid; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_12_io_src_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_12_io_src_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_12_io_src_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_12_io_src_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_12_io_muxes_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_12_io_muxes_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_12_io_muxes_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_12_io_muxes_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_12_io_Osrc_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_12_io_Osrc_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_12_io_Osrc_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_12_io_Osrc_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_12_io_Omuxes_0_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_12_io_Omuxes_0_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_12_io_Omuxes_0_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_12_io_Omuxes_0_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_12_io_Omuxes_1_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_12_io_Omuxes_1_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_12_io_Omuxes_1_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_12_io_Omuxes_2_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_12_io_Omuxes_2_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_12_io_Omuxes_3_0; // @[FlexDPU.scala 124:53]
  wire  MuxesWrapper_13_io_valid; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_13_io_src_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_13_io_src_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_13_io_src_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_13_io_src_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_13_io_muxes_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_13_io_muxes_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_13_io_muxes_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_13_io_muxes_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_13_io_Osrc_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_13_io_Osrc_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_13_io_Osrc_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_13_io_Osrc_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_13_io_Omuxes_0_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_13_io_Omuxes_0_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_13_io_Omuxes_0_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_13_io_Omuxes_0_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_13_io_Omuxes_1_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_13_io_Omuxes_1_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_13_io_Omuxes_1_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_13_io_Omuxes_2_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_13_io_Omuxes_2_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_13_io_Omuxes_3_0; // @[FlexDPU.scala 124:53]
  wire  MuxesWrapper_14_io_valid; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_14_io_src_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_14_io_src_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_14_io_src_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_14_io_src_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_14_io_muxes_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_14_io_muxes_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_14_io_muxes_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_14_io_muxes_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_14_io_Osrc_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_14_io_Osrc_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_14_io_Osrc_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_14_io_Osrc_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_14_io_Omuxes_0_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_14_io_Omuxes_0_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_14_io_Omuxes_0_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_14_io_Omuxes_0_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_14_io_Omuxes_1_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_14_io_Omuxes_1_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_14_io_Omuxes_1_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_14_io_Omuxes_2_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_14_io_Omuxes_2_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_14_io_Omuxes_3_0; // @[FlexDPU.scala 124:53]
  wire  MuxesWrapper_15_io_valid; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_15_io_src_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_15_io_src_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_15_io_src_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_15_io_src_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_15_io_muxes_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_15_io_muxes_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_15_io_muxes_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_15_io_muxes_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_15_io_Osrc_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_15_io_Osrc_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_15_io_Osrc_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_15_io_Osrc_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_15_io_Omuxes_0_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_15_io_Omuxes_0_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_15_io_Omuxes_0_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_15_io_Omuxes_0_3; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_15_io_Omuxes_1_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_15_io_Omuxes_1_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_15_io_Omuxes_1_2; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_15_io_Omuxes_2_0; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_15_io_Omuxes_2_1; // @[FlexDPU.scala 124:53]
  wire [31:0] MuxesWrapper_15_io_Omuxes_3_0; // @[FlexDPU.scala 124:53]
  wire  flexdpecom4_clock; // @[FlexDPU.scala 132:47]
  wire  flexdpecom4_reset; // @[FlexDPU.scala 132:47]
  wire  flexdpecom4_io_i_data_valid; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_io_i_data_bus_0; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_io_i_data_bus_1; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_io_i_data_bus_2; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_io_i_data_bus_3; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_io_i_data_bus2_0; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_io_i_data_bus2_1; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_io_i_data_bus2_2; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_io_i_data_bus2_3; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_io_i_vn_0; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_io_i_vn_1; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_io_i_vn_2; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_io_i_vn_3; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_io_o_adder_0; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_io_o_adder_1; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_io_o_adder_2; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_io_i_mux_bus_0_0; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_io_i_mux_bus_0_1; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_io_i_mux_bus_0_2; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_io_i_mux_bus_0_3; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_io_i_mux_bus_1_0; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_io_i_mux_bus_1_1; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_io_i_mux_bus_1_2; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_io_i_mux_bus_2_0; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_io_i_mux_bus_2_1; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_io_i_mux_bus_3_0; // @[FlexDPU.scala 132:47]
  wire  flexdpecom4_1_clock; // @[FlexDPU.scala 132:47]
  wire  flexdpecom4_1_reset; // @[FlexDPU.scala 132:47]
  wire  flexdpecom4_1_io_i_data_valid; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_1_io_i_data_bus_0; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_1_io_i_data_bus_1; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_1_io_i_data_bus_2; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_1_io_i_data_bus_3; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_1_io_i_data_bus2_0; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_1_io_i_data_bus2_1; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_1_io_i_data_bus2_2; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_1_io_i_data_bus2_3; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_1_io_i_vn_0; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_1_io_i_vn_1; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_1_io_i_vn_2; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_1_io_i_vn_3; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_1_io_o_adder_0; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_1_io_o_adder_1; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_1_io_o_adder_2; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_1_io_i_mux_bus_0_0; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_1_io_i_mux_bus_0_1; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_1_io_i_mux_bus_0_2; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_1_io_i_mux_bus_0_3; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_1_io_i_mux_bus_1_0; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_1_io_i_mux_bus_1_1; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_1_io_i_mux_bus_1_2; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_1_io_i_mux_bus_2_0; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_1_io_i_mux_bus_2_1; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_1_io_i_mux_bus_3_0; // @[FlexDPU.scala 132:47]
  wire  flexdpecom4_2_clock; // @[FlexDPU.scala 132:47]
  wire  flexdpecom4_2_reset; // @[FlexDPU.scala 132:47]
  wire  flexdpecom4_2_io_i_data_valid; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_2_io_i_data_bus_0; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_2_io_i_data_bus_1; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_2_io_i_data_bus_2; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_2_io_i_data_bus_3; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_2_io_i_data_bus2_0; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_2_io_i_data_bus2_1; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_2_io_i_data_bus2_2; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_2_io_i_data_bus2_3; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_2_io_i_vn_0; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_2_io_i_vn_1; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_2_io_i_vn_2; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_2_io_i_vn_3; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_2_io_o_adder_0; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_2_io_o_adder_1; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_2_io_o_adder_2; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_2_io_i_mux_bus_0_0; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_2_io_i_mux_bus_0_1; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_2_io_i_mux_bus_0_2; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_2_io_i_mux_bus_0_3; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_2_io_i_mux_bus_1_0; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_2_io_i_mux_bus_1_1; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_2_io_i_mux_bus_1_2; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_2_io_i_mux_bus_2_0; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_2_io_i_mux_bus_2_1; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_2_io_i_mux_bus_3_0; // @[FlexDPU.scala 132:47]
  wire  flexdpecom4_3_clock; // @[FlexDPU.scala 132:47]
  wire  flexdpecom4_3_reset; // @[FlexDPU.scala 132:47]
  wire  flexdpecom4_3_io_i_data_valid; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_3_io_i_data_bus_0; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_3_io_i_data_bus_1; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_3_io_i_data_bus_2; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_3_io_i_data_bus_3; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_3_io_i_data_bus2_0; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_3_io_i_data_bus2_1; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_3_io_i_data_bus2_2; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_3_io_i_data_bus2_3; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_3_io_i_vn_0; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_3_io_i_vn_1; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_3_io_i_vn_2; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_3_io_i_vn_3; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_3_io_o_adder_0; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_3_io_o_adder_1; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_3_io_o_adder_2; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_3_io_i_mux_bus_0_0; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_3_io_i_mux_bus_0_1; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_3_io_i_mux_bus_0_2; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_3_io_i_mux_bus_0_3; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_3_io_i_mux_bus_1_0; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_3_io_i_mux_bus_1_1; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_3_io_i_mux_bus_1_2; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_3_io_i_mux_bus_2_0; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_3_io_i_mux_bus_2_1; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_3_io_i_mux_bus_3_0; // @[FlexDPU.scala 132:47]
  wire  flexdpecom4_4_clock; // @[FlexDPU.scala 132:47]
  wire  flexdpecom4_4_reset; // @[FlexDPU.scala 132:47]
  wire  flexdpecom4_4_io_i_data_valid; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_4_io_i_data_bus_0; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_4_io_i_data_bus_1; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_4_io_i_data_bus_2; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_4_io_i_data_bus_3; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_4_io_i_data_bus2_0; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_4_io_i_data_bus2_1; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_4_io_i_data_bus2_2; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_4_io_i_data_bus2_3; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_4_io_i_vn_0; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_4_io_i_vn_1; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_4_io_i_vn_2; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_4_io_i_vn_3; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_4_io_o_adder_0; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_4_io_o_adder_1; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_4_io_o_adder_2; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_4_io_i_mux_bus_0_0; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_4_io_i_mux_bus_0_1; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_4_io_i_mux_bus_0_2; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_4_io_i_mux_bus_0_3; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_4_io_i_mux_bus_1_0; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_4_io_i_mux_bus_1_1; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_4_io_i_mux_bus_1_2; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_4_io_i_mux_bus_2_0; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_4_io_i_mux_bus_2_1; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_4_io_i_mux_bus_3_0; // @[FlexDPU.scala 132:47]
  wire  flexdpecom4_5_clock; // @[FlexDPU.scala 132:47]
  wire  flexdpecom4_5_reset; // @[FlexDPU.scala 132:47]
  wire  flexdpecom4_5_io_i_data_valid; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_5_io_i_data_bus_0; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_5_io_i_data_bus_1; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_5_io_i_data_bus_2; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_5_io_i_data_bus_3; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_5_io_i_data_bus2_0; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_5_io_i_data_bus2_1; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_5_io_i_data_bus2_2; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_5_io_i_data_bus2_3; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_5_io_i_vn_0; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_5_io_i_vn_1; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_5_io_i_vn_2; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_5_io_i_vn_3; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_5_io_o_adder_0; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_5_io_o_adder_1; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_5_io_o_adder_2; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_5_io_i_mux_bus_0_0; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_5_io_i_mux_bus_0_1; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_5_io_i_mux_bus_0_2; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_5_io_i_mux_bus_0_3; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_5_io_i_mux_bus_1_0; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_5_io_i_mux_bus_1_1; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_5_io_i_mux_bus_1_2; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_5_io_i_mux_bus_2_0; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_5_io_i_mux_bus_2_1; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_5_io_i_mux_bus_3_0; // @[FlexDPU.scala 132:47]
  wire  flexdpecom4_6_clock; // @[FlexDPU.scala 132:47]
  wire  flexdpecom4_6_reset; // @[FlexDPU.scala 132:47]
  wire  flexdpecom4_6_io_i_data_valid; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_6_io_i_data_bus_0; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_6_io_i_data_bus_1; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_6_io_i_data_bus_2; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_6_io_i_data_bus_3; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_6_io_i_data_bus2_0; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_6_io_i_data_bus2_1; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_6_io_i_data_bus2_2; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_6_io_i_data_bus2_3; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_6_io_i_vn_0; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_6_io_i_vn_1; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_6_io_i_vn_2; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_6_io_i_vn_3; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_6_io_o_adder_0; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_6_io_o_adder_1; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_6_io_o_adder_2; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_6_io_i_mux_bus_0_0; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_6_io_i_mux_bus_0_1; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_6_io_i_mux_bus_0_2; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_6_io_i_mux_bus_0_3; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_6_io_i_mux_bus_1_0; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_6_io_i_mux_bus_1_1; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_6_io_i_mux_bus_1_2; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_6_io_i_mux_bus_2_0; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_6_io_i_mux_bus_2_1; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_6_io_i_mux_bus_3_0; // @[FlexDPU.scala 132:47]
  wire  flexdpecom4_7_clock; // @[FlexDPU.scala 132:47]
  wire  flexdpecom4_7_reset; // @[FlexDPU.scala 132:47]
  wire  flexdpecom4_7_io_i_data_valid; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_7_io_i_data_bus_0; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_7_io_i_data_bus_1; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_7_io_i_data_bus_2; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_7_io_i_data_bus_3; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_7_io_i_data_bus2_0; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_7_io_i_data_bus2_1; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_7_io_i_data_bus2_2; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_7_io_i_data_bus2_3; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_7_io_i_vn_0; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_7_io_i_vn_1; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_7_io_i_vn_2; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_7_io_i_vn_3; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_7_io_o_adder_0; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_7_io_o_adder_1; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_7_io_o_adder_2; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_7_io_i_mux_bus_0_0; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_7_io_i_mux_bus_0_1; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_7_io_i_mux_bus_0_2; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_7_io_i_mux_bus_0_3; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_7_io_i_mux_bus_1_0; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_7_io_i_mux_bus_1_1; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_7_io_i_mux_bus_1_2; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_7_io_i_mux_bus_2_0; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_7_io_i_mux_bus_2_1; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_7_io_i_mux_bus_3_0; // @[FlexDPU.scala 132:47]
  wire  flexdpecom4_8_clock; // @[FlexDPU.scala 132:47]
  wire  flexdpecom4_8_reset; // @[FlexDPU.scala 132:47]
  wire  flexdpecom4_8_io_i_data_valid; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_8_io_i_data_bus_0; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_8_io_i_data_bus_1; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_8_io_i_data_bus_2; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_8_io_i_data_bus_3; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_8_io_i_data_bus2_0; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_8_io_i_data_bus2_1; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_8_io_i_data_bus2_2; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_8_io_i_data_bus2_3; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_8_io_i_vn_0; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_8_io_i_vn_1; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_8_io_i_vn_2; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_8_io_i_vn_3; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_8_io_o_adder_0; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_8_io_o_adder_1; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_8_io_o_adder_2; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_8_io_i_mux_bus_0_0; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_8_io_i_mux_bus_0_1; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_8_io_i_mux_bus_0_2; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_8_io_i_mux_bus_0_3; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_8_io_i_mux_bus_1_0; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_8_io_i_mux_bus_1_1; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_8_io_i_mux_bus_1_2; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_8_io_i_mux_bus_2_0; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_8_io_i_mux_bus_2_1; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_8_io_i_mux_bus_3_0; // @[FlexDPU.scala 132:47]
  wire  flexdpecom4_9_clock; // @[FlexDPU.scala 132:47]
  wire  flexdpecom4_9_reset; // @[FlexDPU.scala 132:47]
  wire  flexdpecom4_9_io_i_data_valid; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_9_io_i_data_bus_0; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_9_io_i_data_bus_1; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_9_io_i_data_bus_2; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_9_io_i_data_bus_3; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_9_io_i_data_bus2_0; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_9_io_i_data_bus2_1; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_9_io_i_data_bus2_2; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_9_io_i_data_bus2_3; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_9_io_i_vn_0; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_9_io_i_vn_1; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_9_io_i_vn_2; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_9_io_i_vn_3; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_9_io_o_adder_0; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_9_io_o_adder_1; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_9_io_o_adder_2; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_9_io_i_mux_bus_0_0; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_9_io_i_mux_bus_0_1; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_9_io_i_mux_bus_0_2; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_9_io_i_mux_bus_0_3; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_9_io_i_mux_bus_1_0; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_9_io_i_mux_bus_1_1; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_9_io_i_mux_bus_1_2; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_9_io_i_mux_bus_2_0; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_9_io_i_mux_bus_2_1; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_9_io_i_mux_bus_3_0; // @[FlexDPU.scala 132:47]
  wire  flexdpecom4_10_clock; // @[FlexDPU.scala 132:47]
  wire  flexdpecom4_10_reset; // @[FlexDPU.scala 132:47]
  wire  flexdpecom4_10_io_i_data_valid; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_10_io_i_data_bus_0; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_10_io_i_data_bus_1; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_10_io_i_data_bus_2; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_10_io_i_data_bus_3; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_10_io_i_data_bus2_0; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_10_io_i_data_bus2_1; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_10_io_i_data_bus2_2; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_10_io_i_data_bus2_3; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_10_io_i_vn_0; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_10_io_i_vn_1; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_10_io_i_vn_2; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_10_io_i_vn_3; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_10_io_o_adder_0; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_10_io_o_adder_1; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_10_io_o_adder_2; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_10_io_i_mux_bus_0_0; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_10_io_i_mux_bus_0_1; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_10_io_i_mux_bus_0_2; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_10_io_i_mux_bus_0_3; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_10_io_i_mux_bus_1_0; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_10_io_i_mux_bus_1_1; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_10_io_i_mux_bus_1_2; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_10_io_i_mux_bus_2_0; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_10_io_i_mux_bus_2_1; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_10_io_i_mux_bus_3_0; // @[FlexDPU.scala 132:47]
  wire  flexdpecom4_11_clock; // @[FlexDPU.scala 132:47]
  wire  flexdpecom4_11_reset; // @[FlexDPU.scala 132:47]
  wire  flexdpecom4_11_io_i_data_valid; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_11_io_i_data_bus_0; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_11_io_i_data_bus_1; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_11_io_i_data_bus_2; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_11_io_i_data_bus_3; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_11_io_i_data_bus2_0; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_11_io_i_data_bus2_1; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_11_io_i_data_bus2_2; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_11_io_i_data_bus2_3; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_11_io_i_vn_0; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_11_io_i_vn_1; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_11_io_i_vn_2; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_11_io_i_vn_3; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_11_io_o_adder_0; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_11_io_o_adder_1; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_11_io_o_adder_2; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_11_io_i_mux_bus_0_0; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_11_io_i_mux_bus_0_1; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_11_io_i_mux_bus_0_2; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_11_io_i_mux_bus_0_3; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_11_io_i_mux_bus_1_0; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_11_io_i_mux_bus_1_1; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_11_io_i_mux_bus_1_2; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_11_io_i_mux_bus_2_0; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_11_io_i_mux_bus_2_1; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_11_io_i_mux_bus_3_0; // @[FlexDPU.scala 132:47]
  wire  flexdpecom4_12_clock; // @[FlexDPU.scala 132:47]
  wire  flexdpecom4_12_reset; // @[FlexDPU.scala 132:47]
  wire  flexdpecom4_12_io_i_data_valid; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_12_io_i_data_bus_0; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_12_io_i_data_bus_1; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_12_io_i_data_bus_2; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_12_io_i_data_bus_3; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_12_io_i_data_bus2_0; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_12_io_i_data_bus2_1; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_12_io_i_data_bus2_2; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_12_io_i_data_bus2_3; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_12_io_i_vn_0; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_12_io_i_vn_1; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_12_io_i_vn_2; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_12_io_i_vn_3; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_12_io_o_adder_0; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_12_io_o_adder_1; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_12_io_o_adder_2; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_12_io_i_mux_bus_0_0; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_12_io_i_mux_bus_0_1; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_12_io_i_mux_bus_0_2; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_12_io_i_mux_bus_0_3; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_12_io_i_mux_bus_1_0; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_12_io_i_mux_bus_1_1; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_12_io_i_mux_bus_1_2; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_12_io_i_mux_bus_2_0; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_12_io_i_mux_bus_2_1; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_12_io_i_mux_bus_3_0; // @[FlexDPU.scala 132:47]
  wire  flexdpecom4_13_clock; // @[FlexDPU.scala 132:47]
  wire  flexdpecom4_13_reset; // @[FlexDPU.scala 132:47]
  wire  flexdpecom4_13_io_i_data_valid; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_13_io_i_data_bus_0; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_13_io_i_data_bus_1; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_13_io_i_data_bus_2; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_13_io_i_data_bus_3; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_13_io_i_data_bus2_0; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_13_io_i_data_bus2_1; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_13_io_i_data_bus2_2; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_13_io_i_data_bus2_3; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_13_io_i_vn_0; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_13_io_i_vn_1; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_13_io_i_vn_2; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_13_io_i_vn_3; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_13_io_o_adder_0; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_13_io_o_adder_1; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_13_io_o_adder_2; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_13_io_i_mux_bus_0_0; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_13_io_i_mux_bus_0_1; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_13_io_i_mux_bus_0_2; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_13_io_i_mux_bus_0_3; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_13_io_i_mux_bus_1_0; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_13_io_i_mux_bus_1_1; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_13_io_i_mux_bus_1_2; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_13_io_i_mux_bus_2_0; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_13_io_i_mux_bus_2_1; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_13_io_i_mux_bus_3_0; // @[FlexDPU.scala 132:47]
  wire  flexdpecom4_14_clock; // @[FlexDPU.scala 132:47]
  wire  flexdpecom4_14_reset; // @[FlexDPU.scala 132:47]
  wire  flexdpecom4_14_io_i_data_valid; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_14_io_i_data_bus_0; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_14_io_i_data_bus_1; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_14_io_i_data_bus_2; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_14_io_i_data_bus_3; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_14_io_i_data_bus2_0; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_14_io_i_data_bus2_1; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_14_io_i_data_bus2_2; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_14_io_i_data_bus2_3; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_14_io_i_vn_0; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_14_io_i_vn_1; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_14_io_i_vn_2; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_14_io_i_vn_3; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_14_io_o_adder_0; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_14_io_o_adder_1; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_14_io_o_adder_2; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_14_io_i_mux_bus_0_0; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_14_io_i_mux_bus_0_1; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_14_io_i_mux_bus_0_2; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_14_io_i_mux_bus_0_3; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_14_io_i_mux_bus_1_0; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_14_io_i_mux_bus_1_1; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_14_io_i_mux_bus_1_2; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_14_io_i_mux_bus_2_0; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_14_io_i_mux_bus_2_1; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_14_io_i_mux_bus_3_0; // @[FlexDPU.scala 132:47]
  wire  flexdpecom4_15_clock; // @[FlexDPU.scala 132:47]
  wire  flexdpecom4_15_reset; // @[FlexDPU.scala 132:47]
  wire  flexdpecom4_15_io_i_data_valid; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_15_io_i_data_bus_0; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_15_io_i_data_bus_1; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_15_io_i_data_bus_2; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_15_io_i_data_bus_3; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_15_io_i_data_bus2_0; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_15_io_i_data_bus2_1; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_15_io_i_data_bus2_2; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_15_io_i_data_bus2_3; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_15_io_i_vn_0; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_15_io_i_vn_1; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_15_io_i_vn_2; // @[FlexDPU.scala 132:47]
  wire [4:0] flexdpecom4_15_io_i_vn_3; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_15_io_o_adder_0; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_15_io_o_adder_1; // @[FlexDPU.scala 132:47]
  wire [15:0] flexdpecom4_15_io_o_adder_2; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_15_io_i_mux_bus_0_0; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_15_io_i_mux_bus_0_1; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_15_io_i_mux_bus_0_2; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_15_io_i_mux_bus_0_3; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_15_io_i_mux_bus_1_0; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_15_io_i_mux_bus_1_1; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_15_io_i_mux_bus_1_2; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_15_io_i_mux_bus_2_0; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_15_io_i_mux_bus_2_1; // @[FlexDPU.scala 132:47]
  wire [3:0] flexdpecom4_15_io_i_mux_bus_3_0; // @[FlexDPU.scala 132:47]
  reg [31:0] used_FlexDPE_0; // @[FlexDPU.scala 19:27]
  reg [31:0] used_FlexDPE_1; // @[FlexDPU.scala 19:27]
  reg [31:0] used_FlexDPE_2; // @[FlexDPU.scala 19:27]
  reg [31:0] used_FlexDPE_3; // @[FlexDPU.scala 19:27]
  reg [31:0] used_FlexDPE_4; // @[FlexDPU.scala 19:27]
  reg [31:0] used_FlexDPE_5; // @[FlexDPU.scala 19:27]
  reg [31:0] used_FlexDPE_6; // @[FlexDPU.scala 19:27]
  reg [31:0] used_FlexDPE_7; // @[FlexDPU.scala 19:27]
  reg [31:0] used_FlexDPE_8; // @[FlexDPU.scala 19:27]
  reg [31:0] used_FlexDPE_9; // @[FlexDPU.scala 19:27]
  reg [31:0] used_FlexDPE_10; // @[FlexDPU.scala 19:27]
  reg [31:0] used_FlexDPE_11; // @[FlexDPU.scala 19:27]
  reg [31:0] used_FlexDPE_12; // @[FlexDPU.scala 19:27]
  reg [31:0] used_FlexDPE_13; // @[FlexDPU.scala 19:27]
  reg [31:0] used_FlexDPE_14; // @[FlexDPU.scala 19:27]
  reg [31:0] used_FlexDPE_15; // @[FlexDPU.scala 19:27]
  wire [31:0] equalDistribution = 32'h10 / 5'h10; // @[FlexDPU.scala 21:39]
  wire [31:0] _GEN_0 = 32'h10 % 32'h10; // @[FlexDPU.scala 22:43]
  wire [4:0] remainingDistribution = _GEN_0[4:0]; // @[FlexDPU.scala 22:43]
  wire [31:0] _used_FlexDPE_0_T_2 = equalDistribution + 32'h1; // @[FlexDPU.scala 25:73]
  reg [31:0] nonZeroValues_0; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_1; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_2; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_3; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_4; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_5; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_6; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_7; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_8; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_9; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_10; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_11; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_12; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_13; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_14; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_15; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_16; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_17; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_18; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_19; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_20; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_21; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_22; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_23; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_24; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_25; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_26; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_27; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_28; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_29; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_30; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_31; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_32; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_33; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_34; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_35; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_36; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_37; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_38; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_39; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_40; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_41; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_42; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_43; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_44; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_45; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_46; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_47; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_48; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_49; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_50; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_51; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_52; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_53; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_54; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_55; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_56; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_57; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_58; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_59; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_60; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_61; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_62; // @[FlexDPU.scala 31:32]
  reg [31:0] nonZeroValues_63; // @[FlexDPU.scala 31:32]
  reg [31:0] index; // @[FlexDPU.scala 32:24]
  reg [31:0] iloop; // @[FlexDPU.scala 33:24]
  reg [31:0] jloop; // @[FlexDPU.scala 34:24]
  reg  Statvalid; // @[FlexDPU.scala 35:28]
  wire  _Statvalid_T_1 = jloop == 32'h7; // @[FlexDPU.scala 37:61]
  wire  _Statvalid_T_2 = iloop == 32'h7 & jloop == 32'h7; // @[FlexDPU.scala 37:51]
  wire [15:0] _GEN_1 = 3'h0 == iloop[2:0] & 3'h1 == jloop[2:0] ? io_Stationary_matrix_0_1 : io_Stationary_matrix_0_0; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_2 = 3'h0 == iloop[2:0] & 3'h2 == jloop[2:0] ? io_Stationary_matrix_0_2 : _GEN_1; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_3 = 3'h0 == iloop[2:0] & 3'h3 == jloop[2:0] ? io_Stationary_matrix_0_3 : _GEN_2; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_4 = 3'h0 == iloop[2:0] & 3'h4 == jloop[2:0] ? io_Stationary_matrix_0_4 : _GEN_3; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_5 = 3'h0 == iloop[2:0] & 3'h5 == jloop[2:0] ? io_Stationary_matrix_0_5 : _GEN_4; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_6 = 3'h0 == iloop[2:0] & 3'h6 == jloop[2:0] ? io_Stationary_matrix_0_6 : _GEN_5; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_7 = 3'h0 == iloop[2:0] & 3'h7 == jloop[2:0] ? io_Stationary_matrix_0_7 : _GEN_6; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_8 = 3'h1 == iloop[2:0] & 3'h0 == jloop[2:0] ? io_Stationary_matrix_1_0 : _GEN_7; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_9 = 3'h1 == iloop[2:0] & 3'h1 == jloop[2:0] ? io_Stationary_matrix_1_1 : _GEN_8; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_10 = 3'h1 == iloop[2:0] & 3'h2 == jloop[2:0] ? io_Stationary_matrix_1_2 : _GEN_9; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_11 = 3'h1 == iloop[2:0] & 3'h3 == jloop[2:0] ? io_Stationary_matrix_1_3 : _GEN_10; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_12 = 3'h1 == iloop[2:0] & 3'h4 == jloop[2:0] ? io_Stationary_matrix_1_4 : _GEN_11; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_13 = 3'h1 == iloop[2:0] & 3'h5 == jloop[2:0] ? io_Stationary_matrix_1_5 : _GEN_12; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_14 = 3'h1 == iloop[2:0] & 3'h6 == jloop[2:0] ? io_Stationary_matrix_1_6 : _GEN_13; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_15 = 3'h1 == iloop[2:0] & 3'h7 == jloop[2:0] ? io_Stationary_matrix_1_7 : _GEN_14; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_16 = 3'h2 == iloop[2:0] & 3'h0 == jloop[2:0] ? io_Stationary_matrix_2_0 : _GEN_15; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_17 = 3'h2 == iloop[2:0] & 3'h1 == jloop[2:0] ? io_Stationary_matrix_2_1 : _GEN_16; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_18 = 3'h2 == iloop[2:0] & 3'h2 == jloop[2:0] ? io_Stationary_matrix_2_2 : _GEN_17; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_19 = 3'h2 == iloop[2:0] & 3'h3 == jloop[2:0] ? io_Stationary_matrix_2_3 : _GEN_18; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_20 = 3'h2 == iloop[2:0] & 3'h4 == jloop[2:0] ? io_Stationary_matrix_2_4 : _GEN_19; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_21 = 3'h2 == iloop[2:0] & 3'h5 == jloop[2:0] ? io_Stationary_matrix_2_5 : _GEN_20; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_22 = 3'h2 == iloop[2:0] & 3'h6 == jloop[2:0] ? io_Stationary_matrix_2_6 : _GEN_21; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_23 = 3'h2 == iloop[2:0] & 3'h7 == jloop[2:0] ? io_Stationary_matrix_2_7 : _GEN_22; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_24 = 3'h3 == iloop[2:0] & 3'h0 == jloop[2:0] ? io_Stationary_matrix_3_0 : _GEN_23; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_25 = 3'h3 == iloop[2:0] & 3'h1 == jloop[2:0] ? io_Stationary_matrix_3_1 : _GEN_24; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_26 = 3'h3 == iloop[2:0] & 3'h2 == jloop[2:0] ? io_Stationary_matrix_3_2 : _GEN_25; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_27 = 3'h3 == iloop[2:0] & 3'h3 == jloop[2:0] ? io_Stationary_matrix_3_3 : _GEN_26; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_28 = 3'h3 == iloop[2:0] & 3'h4 == jloop[2:0] ? io_Stationary_matrix_3_4 : _GEN_27; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_29 = 3'h3 == iloop[2:0] & 3'h5 == jloop[2:0] ? io_Stationary_matrix_3_5 : _GEN_28; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_30 = 3'h3 == iloop[2:0] & 3'h6 == jloop[2:0] ? io_Stationary_matrix_3_6 : _GEN_29; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_31 = 3'h3 == iloop[2:0] & 3'h7 == jloop[2:0] ? io_Stationary_matrix_3_7 : _GEN_30; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_32 = 3'h4 == iloop[2:0] & 3'h0 == jloop[2:0] ? io_Stationary_matrix_4_0 : _GEN_31; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_33 = 3'h4 == iloop[2:0] & 3'h1 == jloop[2:0] ? io_Stationary_matrix_4_1 : _GEN_32; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_34 = 3'h4 == iloop[2:0] & 3'h2 == jloop[2:0] ? io_Stationary_matrix_4_2 : _GEN_33; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_35 = 3'h4 == iloop[2:0] & 3'h3 == jloop[2:0] ? io_Stationary_matrix_4_3 : _GEN_34; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_36 = 3'h4 == iloop[2:0] & 3'h4 == jloop[2:0] ? io_Stationary_matrix_4_4 : _GEN_35; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_37 = 3'h4 == iloop[2:0] & 3'h5 == jloop[2:0] ? io_Stationary_matrix_4_5 : _GEN_36; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_38 = 3'h4 == iloop[2:0] & 3'h6 == jloop[2:0] ? io_Stationary_matrix_4_6 : _GEN_37; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_39 = 3'h4 == iloop[2:0] & 3'h7 == jloop[2:0] ? io_Stationary_matrix_4_7 : _GEN_38; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_40 = 3'h5 == iloop[2:0] & 3'h0 == jloop[2:0] ? io_Stationary_matrix_5_0 : _GEN_39; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_41 = 3'h5 == iloop[2:0] & 3'h1 == jloop[2:0] ? io_Stationary_matrix_5_1 : _GEN_40; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_42 = 3'h5 == iloop[2:0] & 3'h2 == jloop[2:0] ? io_Stationary_matrix_5_2 : _GEN_41; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_43 = 3'h5 == iloop[2:0] & 3'h3 == jloop[2:0] ? io_Stationary_matrix_5_3 : _GEN_42; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_44 = 3'h5 == iloop[2:0] & 3'h4 == jloop[2:0] ? io_Stationary_matrix_5_4 : _GEN_43; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_45 = 3'h5 == iloop[2:0] & 3'h5 == jloop[2:0] ? io_Stationary_matrix_5_5 : _GEN_44; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_46 = 3'h5 == iloop[2:0] & 3'h6 == jloop[2:0] ? io_Stationary_matrix_5_6 : _GEN_45; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_47 = 3'h5 == iloop[2:0] & 3'h7 == jloop[2:0] ? io_Stationary_matrix_5_7 : _GEN_46; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_48 = 3'h6 == iloop[2:0] & 3'h0 == jloop[2:0] ? io_Stationary_matrix_6_0 : _GEN_47; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_49 = 3'h6 == iloop[2:0] & 3'h1 == jloop[2:0] ? io_Stationary_matrix_6_1 : _GEN_48; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_50 = 3'h6 == iloop[2:0] & 3'h2 == jloop[2:0] ? io_Stationary_matrix_6_2 : _GEN_49; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_51 = 3'h6 == iloop[2:0] & 3'h3 == jloop[2:0] ? io_Stationary_matrix_6_3 : _GEN_50; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_52 = 3'h6 == iloop[2:0] & 3'h4 == jloop[2:0] ? io_Stationary_matrix_6_4 : _GEN_51; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_53 = 3'h6 == iloop[2:0] & 3'h5 == jloop[2:0] ? io_Stationary_matrix_6_5 : _GEN_52; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_54 = 3'h6 == iloop[2:0] & 3'h6 == jloop[2:0] ? io_Stationary_matrix_6_6 : _GEN_53; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_55 = 3'h6 == iloop[2:0] & 3'h7 == jloop[2:0] ? io_Stationary_matrix_6_7 : _GEN_54; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_56 = 3'h7 == iloop[2:0] & 3'h0 == jloop[2:0] ? io_Stationary_matrix_7_0 : _GEN_55; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_57 = 3'h7 == iloop[2:0] & 3'h1 == jloop[2:0] ? io_Stationary_matrix_7_1 : _GEN_56; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_58 = 3'h7 == iloop[2:0] & 3'h2 == jloop[2:0] ? io_Stationary_matrix_7_2 : _GEN_57; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_59 = 3'h7 == iloop[2:0] & 3'h3 == jloop[2:0] ? io_Stationary_matrix_7_3 : _GEN_58; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_60 = 3'h7 == iloop[2:0] & 3'h4 == jloop[2:0] ? io_Stationary_matrix_7_4 : _GEN_59; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_61 = 3'h7 == iloop[2:0] & 3'h5 == jloop[2:0] ? io_Stationary_matrix_7_5 : _GEN_60; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_62 = 3'h7 == iloop[2:0] & 3'h6 == jloop[2:0] ? io_Stationary_matrix_7_6 : _GEN_61; // @[FlexDPU.scala 38:{46,46}]
  wire [15:0] _GEN_63 = 3'h7 == iloop[2:0] & 3'h7 == jloop[2:0] ? io_Stationary_matrix_7_7 : _GEN_62; // @[FlexDPU.scala 38:{46,46}]
  wire [31:0] _nonZeroValues_T_3 = {{16'd0}, _GEN_63}; // @[FlexDPU.scala 39:{30,30}]
  wire [31:0] _index_T_1 = index + 32'h1; // @[FlexDPU.scala 40:24]
  wire [31:0] _iloop_T_1 = iloop + 32'h1; // @[FlexDPU.scala 44:24]
  wire [31:0] _jloop_T_1 = jloop + 32'h1; // @[FlexDPU.scala 48:24]
  reg [31:0] PF1_Stream_Col_0; // @[FlexDPU.scala 61:33]
  reg [31:0] PF1_Stream_Col_1; // @[FlexDPU.scala 61:33]
  reg [31:0] PF1_Stream_Col_2; // @[FlexDPU.scala 61:33]
  reg [31:0] PF1_Stream_Col_3; // @[FlexDPU.scala 61:33]
  reg [31:0] PF1_Stream_Col_4; // @[FlexDPU.scala 61:33]
  reg [31:0] PF1_Stream_Col_5; // @[FlexDPU.scala 61:33]
  reg [31:0] PF1_Stream_Col_6; // @[FlexDPU.scala 61:33]
  reg [31:0] PF1_Stream_Col_7; // @[FlexDPU.scala 61:33]
  reg [31:0] ModuleIndex; // @[FlexDPU.scala 62:30]
  reg [31:0] delay; // @[FlexDPU.scala 99:24]
  wire  _GEN_260 = ivntop_io_ProcessValid; // @[FlexDPU.scala 101:28 102:15]
  wire [31:0] _delay_T_1 = delay + 32'h1; // @[FlexDPU.scala 107:20]
  wire  _GEN_262 = delay < 32'hbb8 | _GEN_260; // @[FlexDPU.scala 106:32 108:11]
  wire  check = ivntop_io_ProcessValid | _GEN_262; // @[FlexDPU.scala 104:29 105:11]
  wire  _T_14 = Statvalid & check; // @[FlexDPU.scala 112:20]
  wire [31:0] MuxWrapper_0_Omuxes_0_0 = MuxesWrapper_io_Omuxes_0_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_0_i_mux_bus_0_0_rev_T_2 = {MuxWrapper_0_Omuxes_0_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_0_i_mux_bus_0_0_rev_T_4 = {{1'd0}, MuxWrapper_0_Omuxes_0_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_1788 = {_FDPE_0_i_mux_bus_0_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_0_i_mux_bus_0_0_rev_T_6 = {{1'd0}, _GEN_1788}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_0_i_mux_bus_0_0_rev_T_7 = _FDPE_0_i_mux_bus_0_0_rev_T_2 | _FDPE_0_i_mux_bus_0_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_0_i_mux_bus_0_0_rev_T_8 = {{2'd0}, MuxWrapper_0_Omuxes_0_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_0_i_mux_bus_0_0_rev_T_10 = {_FDPE_0_i_mux_bus_0_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1790 = {{2'd0}, _FDPE_0_i_mux_bus_0_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_0_i_mux_bus_0_0_rev_T_11 = _FDPE_0_i_mux_bus_0_0_rev_T_7 | _GEN_1790; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_0_i_mux_bus_0_0_rev_T_12 = {{3'd0}, MuxWrapper_0_Omuxes_0_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_0_i_mux_bus_0_0_rev_T_14 = {{1'd0}, _FDPE_0_i_mux_bus_0_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1792 = {{2'd0}, _FDPE_0_i_mux_bus_0_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_0_Omuxes_0_1 = MuxesWrapper_io_Omuxes_0_1; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_0_i_mux_bus_0_1_rev_T_2 = {MuxWrapper_0_Omuxes_0_1[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_0_i_mux_bus_0_1_rev_T_4 = {{1'd0}, MuxWrapper_0_Omuxes_0_1[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_1794 = {_FDPE_0_i_mux_bus_0_1_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_0_i_mux_bus_0_1_rev_T_6 = {{1'd0}, _GEN_1794}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_0_i_mux_bus_0_1_rev_T_7 = _FDPE_0_i_mux_bus_0_1_rev_T_2 | _FDPE_0_i_mux_bus_0_1_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_0_i_mux_bus_0_1_rev_T_8 = {{2'd0}, MuxWrapper_0_Omuxes_0_1[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_0_i_mux_bus_0_1_rev_T_10 = {_FDPE_0_i_mux_bus_0_1_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1796 = {{2'd0}, _FDPE_0_i_mux_bus_0_1_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_0_i_mux_bus_0_1_rev_T_11 = _FDPE_0_i_mux_bus_0_1_rev_T_7 | _GEN_1796; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_0_i_mux_bus_0_1_rev_T_12 = {{3'd0}, MuxWrapper_0_Omuxes_0_1[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_0_i_mux_bus_0_1_rev_T_14 = {{1'd0}, _FDPE_0_i_mux_bus_0_1_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1798 = {{2'd0}, _FDPE_0_i_mux_bus_0_1_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_0_Omuxes_0_2 = MuxesWrapper_io_Omuxes_0_2; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_0_i_mux_bus_0_2_rev_T_2 = {MuxWrapper_0_Omuxes_0_2[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_0_i_mux_bus_0_2_rev_T_4 = {{1'd0}, MuxWrapper_0_Omuxes_0_2[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_1800 = {_FDPE_0_i_mux_bus_0_2_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_0_i_mux_bus_0_2_rev_T_6 = {{1'd0}, _GEN_1800}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_0_i_mux_bus_0_2_rev_T_7 = _FDPE_0_i_mux_bus_0_2_rev_T_2 | _FDPE_0_i_mux_bus_0_2_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_0_i_mux_bus_0_2_rev_T_8 = {{2'd0}, MuxWrapper_0_Omuxes_0_2[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_0_i_mux_bus_0_2_rev_T_10 = {_FDPE_0_i_mux_bus_0_2_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1802 = {{2'd0}, _FDPE_0_i_mux_bus_0_2_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_0_i_mux_bus_0_2_rev_T_11 = _FDPE_0_i_mux_bus_0_2_rev_T_7 | _GEN_1802; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_0_i_mux_bus_0_2_rev_T_12 = {{3'd0}, MuxWrapper_0_Omuxes_0_2[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_0_i_mux_bus_0_2_rev_T_14 = {{1'd0}, _FDPE_0_i_mux_bus_0_2_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1804 = {{2'd0}, _FDPE_0_i_mux_bus_0_2_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_0_Omuxes_0_3 = MuxesWrapper_io_Omuxes_0_3; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_0_i_mux_bus_0_3_rev_T_2 = {MuxWrapper_0_Omuxes_0_3[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_0_i_mux_bus_0_3_rev_T_4 = {{1'd0}, MuxWrapper_0_Omuxes_0_3[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_1806 = {_FDPE_0_i_mux_bus_0_3_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_0_i_mux_bus_0_3_rev_T_6 = {{1'd0}, _GEN_1806}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_0_i_mux_bus_0_3_rev_T_7 = _FDPE_0_i_mux_bus_0_3_rev_T_2 | _FDPE_0_i_mux_bus_0_3_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_0_i_mux_bus_0_3_rev_T_8 = {{2'd0}, MuxWrapper_0_Omuxes_0_3[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_0_i_mux_bus_0_3_rev_T_10 = {_FDPE_0_i_mux_bus_0_3_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1808 = {{2'd0}, _FDPE_0_i_mux_bus_0_3_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_0_i_mux_bus_0_3_rev_T_11 = _FDPE_0_i_mux_bus_0_3_rev_T_7 | _GEN_1808; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_0_i_mux_bus_0_3_rev_T_12 = {{3'd0}, MuxWrapper_0_Omuxes_0_3[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_0_i_mux_bus_0_3_rev_T_14 = {{1'd0}, _FDPE_0_i_mux_bus_0_3_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1810 = {{2'd0}, _FDPE_0_i_mux_bus_0_3_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_0_Omuxes_1_0 = MuxesWrapper_io_Omuxes_1_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_0_i_mux_bus_1_0_rev_T_2 = {MuxWrapper_0_Omuxes_1_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_0_i_mux_bus_1_0_rev_T_4 = {{1'd0}, MuxWrapper_0_Omuxes_1_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_1812 = {_FDPE_0_i_mux_bus_1_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_0_i_mux_bus_1_0_rev_T_6 = {{1'd0}, _GEN_1812}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_0_i_mux_bus_1_0_rev_T_7 = _FDPE_0_i_mux_bus_1_0_rev_T_2 | _FDPE_0_i_mux_bus_1_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_0_i_mux_bus_1_0_rev_T_8 = {{2'd0}, MuxWrapper_0_Omuxes_1_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_0_i_mux_bus_1_0_rev_T_10 = {_FDPE_0_i_mux_bus_1_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1814 = {{2'd0}, _FDPE_0_i_mux_bus_1_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_0_i_mux_bus_1_0_rev_T_11 = _FDPE_0_i_mux_bus_1_0_rev_T_7 | _GEN_1814; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_0_i_mux_bus_1_0_rev_T_12 = {{3'd0}, MuxWrapper_0_Omuxes_1_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_0_i_mux_bus_1_0_rev_T_14 = {{1'd0}, _FDPE_0_i_mux_bus_1_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1816 = {{2'd0}, _FDPE_0_i_mux_bus_1_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_0_Omuxes_1_1 = MuxesWrapper_io_Omuxes_1_1; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_0_i_mux_bus_1_1_rev_T_2 = {MuxWrapper_0_Omuxes_1_1[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_0_i_mux_bus_1_1_rev_T_4 = {{1'd0}, MuxWrapper_0_Omuxes_1_1[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_1818 = {_FDPE_0_i_mux_bus_1_1_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_0_i_mux_bus_1_1_rev_T_6 = {{1'd0}, _GEN_1818}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_0_i_mux_bus_1_1_rev_T_7 = _FDPE_0_i_mux_bus_1_1_rev_T_2 | _FDPE_0_i_mux_bus_1_1_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_0_i_mux_bus_1_1_rev_T_8 = {{2'd0}, MuxWrapper_0_Omuxes_1_1[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_0_i_mux_bus_1_1_rev_T_10 = {_FDPE_0_i_mux_bus_1_1_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1820 = {{2'd0}, _FDPE_0_i_mux_bus_1_1_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_0_i_mux_bus_1_1_rev_T_11 = _FDPE_0_i_mux_bus_1_1_rev_T_7 | _GEN_1820; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_0_i_mux_bus_1_1_rev_T_12 = {{3'd0}, MuxWrapper_0_Omuxes_1_1[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_0_i_mux_bus_1_1_rev_T_14 = {{1'd0}, _FDPE_0_i_mux_bus_1_1_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1822 = {{2'd0}, _FDPE_0_i_mux_bus_1_1_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_0_Omuxes_1_2 = MuxesWrapper_io_Omuxes_1_2; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_0_i_mux_bus_1_2_rev_T_2 = {MuxWrapper_0_Omuxes_1_2[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_0_i_mux_bus_1_2_rev_T_4 = {{1'd0}, MuxWrapper_0_Omuxes_1_2[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_1824 = {_FDPE_0_i_mux_bus_1_2_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_0_i_mux_bus_1_2_rev_T_6 = {{1'd0}, _GEN_1824}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_0_i_mux_bus_1_2_rev_T_7 = _FDPE_0_i_mux_bus_1_2_rev_T_2 | _FDPE_0_i_mux_bus_1_2_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_0_i_mux_bus_1_2_rev_T_8 = {{2'd0}, MuxWrapper_0_Omuxes_1_2[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_0_i_mux_bus_1_2_rev_T_10 = {_FDPE_0_i_mux_bus_1_2_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1826 = {{2'd0}, _FDPE_0_i_mux_bus_1_2_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_0_i_mux_bus_1_2_rev_T_11 = _FDPE_0_i_mux_bus_1_2_rev_T_7 | _GEN_1826; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_0_i_mux_bus_1_2_rev_T_12 = {{3'd0}, MuxWrapper_0_Omuxes_1_2[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_0_i_mux_bus_1_2_rev_T_14 = {{1'd0}, _FDPE_0_i_mux_bus_1_2_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1828 = {{2'd0}, _FDPE_0_i_mux_bus_1_2_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_0_Omuxes_2_0 = MuxesWrapper_io_Omuxes_2_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_0_i_mux_bus_2_0_rev_T_2 = {MuxWrapper_0_Omuxes_2_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_0_i_mux_bus_2_0_rev_T_4 = {{1'd0}, MuxWrapper_0_Omuxes_2_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_1830 = {_FDPE_0_i_mux_bus_2_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_0_i_mux_bus_2_0_rev_T_6 = {{1'd0}, _GEN_1830}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_0_i_mux_bus_2_0_rev_T_7 = _FDPE_0_i_mux_bus_2_0_rev_T_2 | _FDPE_0_i_mux_bus_2_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_0_i_mux_bus_2_0_rev_T_8 = {{2'd0}, MuxWrapper_0_Omuxes_2_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_0_i_mux_bus_2_0_rev_T_10 = {_FDPE_0_i_mux_bus_2_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1832 = {{2'd0}, _FDPE_0_i_mux_bus_2_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_0_i_mux_bus_2_0_rev_T_11 = _FDPE_0_i_mux_bus_2_0_rev_T_7 | _GEN_1832; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_0_i_mux_bus_2_0_rev_T_12 = {{3'd0}, MuxWrapper_0_Omuxes_2_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_0_i_mux_bus_2_0_rev_T_14 = {{1'd0}, _FDPE_0_i_mux_bus_2_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1834 = {{2'd0}, _FDPE_0_i_mux_bus_2_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_0_Omuxes_2_1 = MuxesWrapper_io_Omuxes_2_1; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_0_i_mux_bus_2_1_rev_T_2 = {MuxWrapper_0_Omuxes_2_1[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_0_i_mux_bus_2_1_rev_T_4 = {{1'd0}, MuxWrapper_0_Omuxes_2_1[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_1836 = {_FDPE_0_i_mux_bus_2_1_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_0_i_mux_bus_2_1_rev_T_6 = {{1'd0}, _GEN_1836}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_0_i_mux_bus_2_1_rev_T_7 = _FDPE_0_i_mux_bus_2_1_rev_T_2 | _FDPE_0_i_mux_bus_2_1_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_0_i_mux_bus_2_1_rev_T_8 = {{2'd0}, MuxWrapper_0_Omuxes_2_1[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_0_i_mux_bus_2_1_rev_T_10 = {_FDPE_0_i_mux_bus_2_1_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1838 = {{2'd0}, _FDPE_0_i_mux_bus_2_1_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_0_i_mux_bus_2_1_rev_T_11 = _FDPE_0_i_mux_bus_2_1_rev_T_7 | _GEN_1838; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_0_i_mux_bus_2_1_rev_T_12 = {{3'd0}, MuxWrapper_0_Omuxes_2_1[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_0_i_mux_bus_2_1_rev_T_14 = {{1'd0}, _FDPE_0_i_mux_bus_2_1_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1840 = {{2'd0}, _FDPE_0_i_mux_bus_2_1_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_0_Omuxes_3_0 = MuxesWrapper_io_Omuxes_3_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_0_i_mux_bus_3_0_rev_T_2 = {MuxWrapper_0_Omuxes_3_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_0_i_mux_bus_3_0_rev_T_4 = {{1'd0}, MuxWrapper_0_Omuxes_3_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_1842 = {_FDPE_0_i_mux_bus_3_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_0_i_mux_bus_3_0_rev_T_6 = {{1'd0}, _GEN_1842}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_0_i_mux_bus_3_0_rev_T_7 = _FDPE_0_i_mux_bus_3_0_rev_T_2 | _FDPE_0_i_mux_bus_3_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_0_i_mux_bus_3_0_rev_T_8 = {{2'd0}, MuxWrapper_0_Omuxes_3_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_0_i_mux_bus_3_0_rev_T_10 = {_FDPE_0_i_mux_bus_3_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1844 = {{2'd0}, _FDPE_0_i_mux_bus_3_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_0_i_mux_bus_3_0_rev_T_11 = _FDPE_0_i_mux_bus_3_0_rev_T_7 | _GEN_1844; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_0_i_mux_bus_3_0_rev_T_12 = {{3'd0}, MuxWrapper_0_Omuxes_3_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_0_i_mux_bus_3_0_rev_T_14 = {{1'd0}, _FDPE_0_i_mux_bus_3_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1846 = {{2'd0}, _FDPE_0_i_mux_bus_3_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_1_Omuxes_0_0 = MuxesWrapper_1_io_Omuxes_0_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_1_i_mux_bus_0_0_rev_T_2 = {MuxWrapper_1_Omuxes_0_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_1_i_mux_bus_0_0_rev_T_4 = {{1'd0}, MuxWrapper_1_Omuxes_0_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_1848 = {_FDPE_1_i_mux_bus_0_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_1_i_mux_bus_0_0_rev_T_6 = {{1'd0}, _GEN_1848}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_1_i_mux_bus_0_0_rev_T_7 = _FDPE_1_i_mux_bus_0_0_rev_T_2 | _FDPE_1_i_mux_bus_0_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_1_i_mux_bus_0_0_rev_T_8 = {{2'd0}, MuxWrapper_1_Omuxes_0_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_1_i_mux_bus_0_0_rev_T_10 = {_FDPE_1_i_mux_bus_0_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1850 = {{2'd0}, _FDPE_1_i_mux_bus_0_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_1_i_mux_bus_0_0_rev_T_11 = _FDPE_1_i_mux_bus_0_0_rev_T_7 | _GEN_1850; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_1_i_mux_bus_0_0_rev_T_12 = {{3'd0}, MuxWrapper_1_Omuxes_0_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_1_i_mux_bus_0_0_rev_T_14 = {{1'd0}, _FDPE_1_i_mux_bus_0_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1852 = {{2'd0}, _FDPE_1_i_mux_bus_0_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_1_Omuxes_0_1 = MuxesWrapper_1_io_Omuxes_0_1; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_1_i_mux_bus_0_1_rev_T_2 = {MuxWrapper_1_Omuxes_0_1[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_1_i_mux_bus_0_1_rev_T_4 = {{1'd0}, MuxWrapper_1_Omuxes_0_1[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_1854 = {_FDPE_1_i_mux_bus_0_1_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_1_i_mux_bus_0_1_rev_T_6 = {{1'd0}, _GEN_1854}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_1_i_mux_bus_0_1_rev_T_7 = _FDPE_1_i_mux_bus_0_1_rev_T_2 | _FDPE_1_i_mux_bus_0_1_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_1_i_mux_bus_0_1_rev_T_8 = {{2'd0}, MuxWrapper_1_Omuxes_0_1[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_1_i_mux_bus_0_1_rev_T_10 = {_FDPE_1_i_mux_bus_0_1_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1856 = {{2'd0}, _FDPE_1_i_mux_bus_0_1_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_1_i_mux_bus_0_1_rev_T_11 = _FDPE_1_i_mux_bus_0_1_rev_T_7 | _GEN_1856; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_1_i_mux_bus_0_1_rev_T_12 = {{3'd0}, MuxWrapper_1_Omuxes_0_1[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_1_i_mux_bus_0_1_rev_T_14 = {{1'd0}, _FDPE_1_i_mux_bus_0_1_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1858 = {{2'd0}, _FDPE_1_i_mux_bus_0_1_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_1_Omuxes_0_2 = MuxesWrapper_1_io_Omuxes_0_2; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_1_i_mux_bus_0_2_rev_T_2 = {MuxWrapper_1_Omuxes_0_2[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_1_i_mux_bus_0_2_rev_T_4 = {{1'd0}, MuxWrapper_1_Omuxes_0_2[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_1860 = {_FDPE_1_i_mux_bus_0_2_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_1_i_mux_bus_0_2_rev_T_6 = {{1'd0}, _GEN_1860}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_1_i_mux_bus_0_2_rev_T_7 = _FDPE_1_i_mux_bus_0_2_rev_T_2 | _FDPE_1_i_mux_bus_0_2_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_1_i_mux_bus_0_2_rev_T_8 = {{2'd0}, MuxWrapper_1_Omuxes_0_2[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_1_i_mux_bus_0_2_rev_T_10 = {_FDPE_1_i_mux_bus_0_2_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1862 = {{2'd0}, _FDPE_1_i_mux_bus_0_2_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_1_i_mux_bus_0_2_rev_T_11 = _FDPE_1_i_mux_bus_0_2_rev_T_7 | _GEN_1862; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_1_i_mux_bus_0_2_rev_T_12 = {{3'd0}, MuxWrapper_1_Omuxes_0_2[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_1_i_mux_bus_0_2_rev_T_14 = {{1'd0}, _FDPE_1_i_mux_bus_0_2_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1864 = {{2'd0}, _FDPE_1_i_mux_bus_0_2_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_1_Omuxes_0_3 = MuxesWrapper_1_io_Omuxes_0_3; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_1_i_mux_bus_0_3_rev_T_2 = {MuxWrapper_1_Omuxes_0_3[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_1_i_mux_bus_0_3_rev_T_4 = {{1'd0}, MuxWrapper_1_Omuxes_0_3[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_1866 = {_FDPE_1_i_mux_bus_0_3_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_1_i_mux_bus_0_3_rev_T_6 = {{1'd0}, _GEN_1866}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_1_i_mux_bus_0_3_rev_T_7 = _FDPE_1_i_mux_bus_0_3_rev_T_2 | _FDPE_1_i_mux_bus_0_3_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_1_i_mux_bus_0_3_rev_T_8 = {{2'd0}, MuxWrapper_1_Omuxes_0_3[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_1_i_mux_bus_0_3_rev_T_10 = {_FDPE_1_i_mux_bus_0_3_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1868 = {{2'd0}, _FDPE_1_i_mux_bus_0_3_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_1_i_mux_bus_0_3_rev_T_11 = _FDPE_1_i_mux_bus_0_3_rev_T_7 | _GEN_1868; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_1_i_mux_bus_0_3_rev_T_12 = {{3'd0}, MuxWrapper_1_Omuxes_0_3[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_1_i_mux_bus_0_3_rev_T_14 = {{1'd0}, _FDPE_1_i_mux_bus_0_3_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1870 = {{2'd0}, _FDPE_1_i_mux_bus_0_3_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_1_Omuxes_1_0 = MuxesWrapper_1_io_Omuxes_1_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_1_i_mux_bus_1_0_rev_T_2 = {MuxWrapper_1_Omuxes_1_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_1_i_mux_bus_1_0_rev_T_4 = {{1'd0}, MuxWrapper_1_Omuxes_1_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_1872 = {_FDPE_1_i_mux_bus_1_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_1_i_mux_bus_1_0_rev_T_6 = {{1'd0}, _GEN_1872}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_1_i_mux_bus_1_0_rev_T_7 = _FDPE_1_i_mux_bus_1_0_rev_T_2 | _FDPE_1_i_mux_bus_1_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_1_i_mux_bus_1_0_rev_T_8 = {{2'd0}, MuxWrapper_1_Omuxes_1_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_1_i_mux_bus_1_0_rev_T_10 = {_FDPE_1_i_mux_bus_1_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1874 = {{2'd0}, _FDPE_1_i_mux_bus_1_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_1_i_mux_bus_1_0_rev_T_11 = _FDPE_1_i_mux_bus_1_0_rev_T_7 | _GEN_1874; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_1_i_mux_bus_1_0_rev_T_12 = {{3'd0}, MuxWrapper_1_Omuxes_1_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_1_i_mux_bus_1_0_rev_T_14 = {{1'd0}, _FDPE_1_i_mux_bus_1_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1876 = {{2'd0}, _FDPE_1_i_mux_bus_1_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_1_Omuxes_1_1 = MuxesWrapper_1_io_Omuxes_1_1; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_1_i_mux_bus_1_1_rev_T_2 = {MuxWrapper_1_Omuxes_1_1[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_1_i_mux_bus_1_1_rev_T_4 = {{1'd0}, MuxWrapper_1_Omuxes_1_1[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_1878 = {_FDPE_1_i_mux_bus_1_1_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_1_i_mux_bus_1_1_rev_T_6 = {{1'd0}, _GEN_1878}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_1_i_mux_bus_1_1_rev_T_7 = _FDPE_1_i_mux_bus_1_1_rev_T_2 | _FDPE_1_i_mux_bus_1_1_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_1_i_mux_bus_1_1_rev_T_8 = {{2'd0}, MuxWrapper_1_Omuxes_1_1[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_1_i_mux_bus_1_1_rev_T_10 = {_FDPE_1_i_mux_bus_1_1_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1880 = {{2'd0}, _FDPE_1_i_mux_bus_1_1_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_1_i_mux_bus_1_1_rev_T_11 = _FDPE_1_i_mux_bus_1_1_rev_T_7 | _GEN_1880; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_1_i_mux_bus_1_1_rev_T_12 = {{3'd0}, MuxWrapper_1_Omuxes_1_1[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_1_i_mux_bus_1_1_rev_T_14 = {{1'd0}, _FDPE_1_i_mux_bus_1_1_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1882 = {{2'd0}, _FDPE_1_i_mux_bus_1_1_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_1_Omuxes_1_2 = MuxesWrapper_1_io_Omuxes_1_2; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_1_i_mux_bus_1_2_rev_T_2 = {MuxWrapper_1_Omuxes_1_2[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_1_i_mux_bus_1_2_rev_T_4 = {{1'd0}, MuxWrapper_1_Omuxes_1_2[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_1884 = {_FDPE_1_i_mux_bus_1_2_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_1_i_mux_bus_1_2_rev_T_6 = {{1'd0}, _GEN_1884}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_1_i_mux_bus_1_2_rev_T_7 = _FDPE_1_i_mux_bus_1_2_rev_T_2 | _FDPE_1_i_mux_bus_1_2_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_1_i_mux_bus_1_2_rev_T_8 = {{2'd0}, MuxWrapper_1_Omuxes_1_2[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_1_i_mux_bus_1_2_rev_T_10 = {_FDPE_1_i_mux_bus_1_2_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1886 = {{2'd0}, _FDPE_1_i_mux_bus_1_2_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_1_i_mux_bus_1_2_rev_T_11 = _FDPE_1_i_mux_bus_1_2_rev_T_7 | _GEN_1886; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_1_i_mux_bus_1_2_rev_T_12 = {{3'd0}, MuxWrapper_1_Omuxes_1_2[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_1_i_mux_bus_1_2_rev_T_14 = {{1'd0}, _FDPE_1_i_mux_bus_1_2_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1888 = {{2'd0}, _FDPE_1_i_mux_bus_1_2_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_1_Omuxes_2_0 = MuxesWrapper_1_io_Omuxes_2_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_1_i_mux_bus_2_0_rev_T_2 = {MuxWrapper_1_Omuxes_2_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_1_i_mux_bus_2_0_rev_T_4 = {{1'd0}, MuxWrapper_1_Omuxes_2_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_1890 = {_FDPE_1_i_mux_bus_2_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_1_i_mux_bus_2_0_rev_T_6 = {{1'd0}, _GEN_1890}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_1_i_mux_bus_2_0_rev_T_7 = _FDPE_1_i_mux_bus_2_0_rev_T_2 | _FDPE_1_i_mux_bus_2_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_1_i_mux_bus_2_0_rev_T_8 = {{2'd0}, MuxWrapper_1_Omuxes_2_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_1_i_mux_bus_2_0_rev_T_10 = {_FDPE_1_i_mux_bus_2_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1892 = {{2'd0}, _FDPE_1_i_mux_bus_2_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_1_i_mux_bus_2_0_rev_T_11 = _FDPE_1_i_mux_bus_2_0_rev_T_7 | _GEN_1892; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_1_i_mux_bus_2_0_rev_T_12 = {{3'd0}, MuxWrapper_1_Omuxes_2_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_1_i_mux_bus_2_0_rev_T_14 = {{1'd0}, _FDPE_1_i_mux_bus_2_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1894 = {{2'd0}, _FDPE_1_i_mux_bus_2_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_1_Omuxes_2_1 = MuxesWrapper_1_io_Omuxes_2_1; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_1_i_mux_bus_2_1_rev_T_2 = {MuxWrapper_1_Omuxes_2_1[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_1_i_mux_bus_2_1_rev_T_4 = {{1'd0}, MuxWrapper_1_Omuxes_2_1[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_1896 = {_FDPE_1_i_mux_bus_2_1_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_1_i_mux_bus_2_1_rev_T_6 = {{1'd0}, _GEN_1896}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_1_i_mux_bus_2_1_rev_T_7 = _FDPE_1_i_mux_bus_2_1_rev_T_2 | _FDPE_1_i_mux_bus_2_1_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_1_i_mux_bus_2_1_rev_T_8 = {{2'd0}, MuxWrapper_1_Omuxes_2_1[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_1_i_mux_bus_2_1_rev_T_10 = {_FDPE_1_i_mux_bus_2_1_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1898 = {{2'd0}, _FDPE_1_i_mux_bus_2_1_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_1_i_mux_bus_2_1_rev_T_11 = _FDPE_1_i_mux_bus_2_1_rev_T_7 | _GEN_1898; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_1_i_mux_bus_2_1_rev_T_12 = {{3'd0}, MuxWrapper_1_Omuxes_2_1[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_1_i_mux_bus_2_1_rev_T_14 = {{1'd0}, _FDPE_1_i_mux_bus_2_1_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1900 = {{2'd0}, _FDPE_1_i_mux_bus_2_1_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_1_Omuxes_3_0 = MuxesWrapper_1_io_Omuxes_3_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_1_i_mux_bus_3_0_rev_T_2 = {MuxWrapper_1_Omuxes_3_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_1_i_mux_bus_3_0_rev_T_4 = {{1'd0}, MuxWrapper_1_Omuxes_3_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_1902 = {_FDPE_1_i_mux_bus_3_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_1_i_mux_bus_3_0_rev_T_6 = {{1'd0}, _GEN_1902}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_1_i_mux_bus_3_0_rev_T_7 = _FDPE_1_i_mux_bus_3_0_rev_T_2 | _FDPE_1_i_mux_bus_3_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_1_i_mux_bus_3_0_rev_T_8 = {{2'd0}, MuxWrapper_1_Omuxes_3_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_1_i_mux_bus_3_0_rev_T_10 = {_FDPE_1_i_mux_bus_3_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1904 = {{2'd0}, _FDPE_1_i_mux_bus_3_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_1_i_mux_bus_3_0_rev_T_11 = _FDPE_1_i_mux_bus_3_0_rev_T_7 | _GEN_1904; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_1_i_mux_bus_3_0_rev_T_12 = {{3'd0}, MuxWrapper_1_Omuxes_3_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_1_i_mux_bus_3_0_rev_T_14 = {{1'd0}, _FDPE_1_i_mux_bus_3_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1906 = {{2'd0}, _FDPE_1_i_mux_bus_3_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_2_Omuxes_0_0 = MuxesWrapper_2_io_Omuxes_0_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_2_i_mux_bus_0_0_rev_T_2 = {MuxWrapper_2_Omuxes_0_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_2_i_mux_bus_0_0_rev_T_4 = {{1'd0}, MuxWrapper_2_Omuxes_0_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_1908 = {_FDPE_2_i_mux_bus_0_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_2_i_mux_bus_0_0_rev_T_6 = {{1'd0}, _GEN_1908}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_2_i_mux_bus_0_0_rev_T_7 = _FDPE_2_i_mux_bus_0_0_rev_T_2 | _FDPE_2_i_mux_bus_0_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_2_i_mux_bus_0_0_rev_T_8 = {{2'd0}, MuxWrapper_2_Omuxes_0_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_2_i_mux_bus_0_0_rev_T_10 = {_FDPE_2_i_mux_bus_0_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1910 = {{2'd0}, _FDPE_2_i_mux_bus_0_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_2_i_mux_bus_0_0_rev_T_11 = _FDPE_2_i_mux_bus_0_0_rev_T_7 | _GEN_1910; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_2_i_mux_bus_0_0_rev_T_12 = {{3'd0}, MuxWrapper_2_Omuxes_0_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_2_i_mux_bus_0_0_rev_T_14 = {{1'd0}, _FDPE_2_i_mux_bus_0_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1912 = {{2'd0}, _FDPE_2_i_mux_bus_0_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_2_Omuxes_0_1 = MuxesWrapper_2_io_Omuxes_0_1; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_2_i_mux_bus_0_1_rev_T_2 = {MuxWrapper_2_Omuxes_0_1[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_2_i_mux_bus_0_1_rev_T_4 = {{1'd0}, MuxWrapper_2_Omuxes_0_1[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_1914 = {_FDPE_2_i_mux_bus_0_1_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_2_i_mux_bus_0_1_rev_T_6 = {{1'd0}, _GEN_1914}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_2_i_mux_bus_0_1_rev_T_7 = _FDPE_2_i_mux_bus_0_1_rev_T_2 | _FDPE_2_i_mux_bus_0_1_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_2_i_mux_bus_0_1_rev_T_8 = {{2'd0}, MuxWrapper_2_Omuxes_0_1[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_2_i_mux_bus_0_1_rev_T_10 = {_FDPE_2_i_mux_bus_0_1_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1916 = {{2'd0}, _FDPE_2_i_mux_bus_0_1_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_2_i_mux_bus_0_1_rev_T_11 = _FDPE_2_i_mux_bus_0_1_rev_T_7 | _GEN_1916; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_2_i_mux_bus_0_1_rev_T_12 = {{3'd0}, MuxWrapper_2_Omuxes_0_1[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_2_i_mux_bus_0_1_rev_T_14 = {{1'd0}, _FDPE_2_i_mux_bus_0_1_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1918 = {{2'd0}, _FDPE_2_i_mux_bus_0_1_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_2_Omuxes_0_2 = MuxesWrapper_2_io_Omuxes_0_2; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_2_i_mux_bus_0_2_rev_T_2 = {MuxWrapper_2_Omuxes_0_2[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_2_i_mux_bus_0_2_rev_T_4 = {{1'd0}, MuxWrapper_2_Omuxes_0_2[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_1920 = {_FDPE_2_i_mux_bus_0_2_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_2_i_mux_bus_0_2_rev_T_6 = {{1'd0}, _GEN_1920}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_2_i_mux_bus_0_2_rev_T_7 = _FDPE_2_i_mux_bus_0_2_rev_T_2 | _FDPE_2_i_mux_bus_0_2_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_2_i_mux_bus_0_2_rev_T_8 = {{2'd0}, MuxWrapper_2_Omuxes_0_2[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_2_i_mux_bus_0_2_rev_T_10 = {_FDPE_2_i_mux_bus_0_2_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1922 = {{2'd0}, _FDPE_2_i_mux_bus_0_2_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_2_i_mux_bus_0_2_rev_T_11 = _FDPE_2_i_mux_bus_0_2_rev_T_7 | _GEN_1922; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_2_i_mux_bus_0_2_rev_T_12 = {{3'd0}, MuxWrapper_2_Omuxes_0_2[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_2_i_mux_bus_0_2_rev_T_14 = {{1'd0}, _FDPE_2_i_mux_bus_0_2_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1924 = {{2'd0}, _FDPE_2_i_mux_bus_0_2_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_2_Omuxes_0_3 = MuxesWrapper_2_io_Omuxes_0_3; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_2_i_mux_bus_0_3_rev_T_2 = {MuxWrapper_2_Omuxes_0_3[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_2_i_mux_bus_0_3_rev_T_4 = {{1'd0}, MuxWrapper_2_Omuxes_0_3[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_1926 = {_FDPE_2_i_mux_bus_0_3_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_2_i_mux_bus_0_3_rev_T_6 = {{1'd0}, _GEN_1926}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_2_i_mux_bus_0_3_rev_T_7 = _FDPE_2_i_mux_bus_0_3_rev_T_2 | _FDPE_2_i_mux_bus_0_3_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_2_i_mux_bus_0_3_rev_T_8 = {{2'd0}, MuxWrapper_2_Omuxes_0_3[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_2_i_mux_bus_0_3_rev_T_10 = {_FDPE_2_i_mux_bus_0_3_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1928 = {{2'd0}, _FDPE_2_i_mux_bus_0_3_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_2_i_mux_bus_0_3_rev_T_11 = _FDPE_2_i_mux_bus_0_3_rev_T_7 | _GEN_1928; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_2_i_mux_bus_0_3_rev_T_12 = {{3'd0}, MuxWrapper_2_Omuxes_0_3[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_2_i_mux_bus_0_3_rev_T_14 = {{1'd0}, _FDPE_2_i_mux_bus_0_3_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1930 = {{2'd0}, _FDPE_2_i_mux_bus_0_3_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_2_Omuxes_1_0 = MuxesWrapper_2_io_Omuxes_1_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_2_i_mux_bus_1_0_rev_T_2 = {MuxWrapper_2_Omuxes_1_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_2_i_mux_bus_1_0_rev_T_4 = {{1'd0}, MuxWrapper_2_Omuxes_1_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_1932 = {_FDPE_2_i_mux_bus_1_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_2_i_mux_bus_1_0_rev_T_6 = {{1'd0}, _GEN_1932}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_2_i_mux_bus_1_0_rev_T_7 = _FDPE_2_i_mux_bus_1_0_rev_T_2 | _FDPE_2_i_mux_bus_1_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_2_i_mux_bus_1_0_rev_T_8 = {{2'd0}, MuxWrapper_2_Omuxes_1_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_2_i_mux_bus_1_0_rev_T_10 = {_FDPE_2_i_mux_bus_1_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1934 = {{2'd0}, _FDPE_2_i_mux_bus_1_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_2_i_mux_bus_1_0_rev_T_11 = _FDPE_2_i_mux_bus_1_0_rev_T_7 | _GEN_1934; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_2_i_mux_bus_1_0_rev_T_12 = {{3'd0}, MuxWrapper_2_Omuxes_1_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_2_i_mux_bus_1_0_rev_T_14 = {{1'd0}, _FDPE_2_i_mux_bus_1_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1936 = {{2'd0}, _FDPE_2_i_mux_bus_1_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_2_Omuxes_1_1 = MuxesWrapper_2_io_Omuxes_1_1; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_2_i_mux_bus_1_1_rev_T_2 = {MuxWrapper_2_Omuxes_1_1[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_2_i_mux_bus_1_1_rev_T_4 = {{1'd0}, MuxWrapper_2_Omuxes_1_1[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_1938 = {_FDPE_2_i_mux_bus_1_1_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_2_i_mux_bus_1_1_rev_T_6 = {{1'd0}, _GEN_1938}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_2_i_mux_bus_1_1_rev_T_7 = _FDPE_2_i_mux_bus_1_1_rev_T_2 | _FDPE_2_i_mux_bus_1_1_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_2_i_mux_bus_1_1_rev_T_8 = {{2'd0}, MuxWrapper_2_Omuxes_1_1[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_2_i_mux_bus_1_1_rev_T_10 = {_FDPE_2_i_mux_bus_1_1_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1940 = {{2'd0}, _FDPE_2_i_mux_bus_1_1_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_2_i_mux_bus_1_1_rev_T_11 = _FDPE_2_i_mux_bus_1_1_rev_T_7 | _GEN_1940; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_2_i_mux_bus_1_1_rev_T_12 = {{3'd0}, MuxWrapper_2_Omuxes_1_1[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_2_i_mux_bus_1_1_rev_T_14 = {{1'd0}, _FDPE_2_i_mux_bus_1_1_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1942 = {{2'd0}, _FDPE_2_i_mux_bus_1_1_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_2_Omuxes_1_2 = MuxesWrapper_2_io_Omuxes_1_2; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_2_i_mux_bus_1_2_rev_T_2 = {MuxWrapper_2_Omuxes_1_2[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_2_i_mux_bus_1_2_rev_T_4 = {{1'd0}, MuxWrapper_2_Omuxes_1_2[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_1944 = {_FDPE_2_i_mux_bus_1_2_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_2_i_mux_bus_1_2_rev_T_6 = {{1'd0}, _GEN_1944}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_2_i_mux_bus_1_2_rev_T_7 = _FDPE_2_i_mux_bus_1_2_rev_T_2 | _FDPE_2_i_mux_bus_1_2_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_2_i_mux_bus_1_2_rev_T_8 = {{2'd0}, MuxWrapper_2_Omuxes_1_2[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_2_i_mux_bus_1_2_rev_T_10 = {_FDPE_2_i_mux_bus_1_2_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1946 = {{2'd0}, _FDPE_2_i_mux_bus_1_2_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_2_i_mux_bus_1_2_rev_T_11 = _FDPE_2_i_mux_bus_1_2_rev_T_7 | _GEN_1946; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_2_i_mux_bus_1_2_rev_T_12 = {{3'd0}, MuxWrapper_2_Omuxes_1_2[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_2_i_mux_bus_1_2_rev_T_14 = {{1'd0}, _FDPE_2_i_mux_bus_1_2_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1948 = {{2'd0}, _FDPE_2_i_mux_bus_1_2_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_2_Omuxes_2_0 = MuxesWrapper_2_io_Omuxes_2_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_2_i_mux_bus_2_0_rev_T_2 = {MuxWrapper_2_Omuxes_2_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_2_i_mux_bus_2_0_rev_T_4 = {{1'd0}, MuxWrapper_2_Omuxes_2_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_1950 = {_FDPE_2_i_mux_bus_2_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_2_i_mux_bus_2_0_rev_T_6 = {{1'd0}, _GEN_1950}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_2_i_mux_bus_2_0_rev_T_7 = _FDPE_2_i_mux_bus_2_0_rev_T_2 | _FDPE_2_i_mux_bus_2_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_2_i_mux_bus_2_0_rev_T_8 = {{2'd0}, MuxWrapper_2_Omuxes_2_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_2_i_mux_bus_2_0_rev_T_10 = {_FDPE_2_i_mux_bus_2_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1952 = {{2'd0}, _FDPE_2_i_mux_bus_2_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_2_i_mux_bus_2_0_rev_T_11 = _FDPE_2_i_mux_bus_2_0_rev_T_7 | _GEN_1952; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_2_i_mux_bus_2_0_rev_T_12 = {{3'd0}, MuxWrapper_2_Omuxes_2_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_2_i_mux_bus_2_0_rev_T_14 = {{1'd0}, _FDPE_2_i_mux_bus_2_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1954 = {{2'd0}, _FDPE_2_i_mux_bus_2_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_2_Omuxes_2_1 = MuxesWrapper_2_io_Omuxes_2_1; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_2_i_mux_bus_2_1_rev_T_2 = {MuxWrapper_2_Omuxes_2_1[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_2_i_mux_bus_2_1_rev_T_4 = {{1'd0}, MuxWrapper_2_Omuxes_2_1[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_1956 = {_FDPE_2_i_mux_bus_2_1_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_2_i_mux_bus_2_1_rev_T_6 = {{1'd0}, _GEN_1956}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_2_i_mux_bus_2_1_rev_T_7 = _FDPE_2_i_mux_bus_2_1_rev_T_2 | _FDPE_2_i_mux_bus_2_1_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_2_i_mux_bus_2_1_rev_T_8 = {{2'd0}, MuxWrapper_2_Omuxes_2_1[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_2_i_mux_bus_2_1_rev_T_10 = {_FDPE_2_i_mux_bus_2_1_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1958 = {{2'd0}, _FDPE_2_i_mux_bus_2_1_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_2_i_mux_bus_2_1_rev_T_11 = _FDPE_2_i_mux_bus_2_1_rev_T_7 | _GEN_1958; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_2_i_mux_bus_2_1_rev_T_12 = {{3'd0}, MuxWrapper_2_Omuxes_2_1[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_2_i_mux_bus_2_1_rev_T_14 = {{1'd0}, _FDPE_2_i_mux_bus_2_1_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1960 = {{2'd0}, _FDPE_2_i_mux_bus_2_1_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_2_Omuxes_3_0 = MuxesWrapper_2_io_Omuxes_3_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_2_i_mux_bus_3_0_rev_T_2 = {MuxWrapper_2_Omuxes_3_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_2_i_mux_bus_3_0_rev_T_4 = {{1'd0}, MuxWrapper_2_Omuxes_3_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_1962 = {_FDPE_2_i_mux_bus_3_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_2_i_mux_bus_3_0_rev_T_6 = {{1'd0}, _GEN_1962}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_2_i_mux_bus_3_0_rev_T_7 = _FDPE_2_i_mux_bus_3_0_rev_T_2 | _FDPE_2_i_mux_bus_3_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_2_i_mux_bus_3_0_rev_T_8 = {{2'd0}, MuxWrapper_2_Omuxes_3_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_2_i_mux_bus_3_0_rev_T_10 = {_FDPE_2_i_mux_bus_3_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1964 = {{2'd0}, _FDPE_2_i_mux_bus_3_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_2_i_mux_bus_3_0_rev_T_11 = _FDPE_2_i_mux_bus_3_0_rev_T_7 | _GEN_1964; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_2_i_mux_bus_3_0_rev_T_12 = {{3'd0}, MuxWrapper_2_Omuxes_3_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_2_i_mux_bus_3_0_rev_T_14 = {{1'd0}, _FDPE_2_i_mux_bus_3_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1966 = {{2'd0}, _FDPE_2_i_mux_bus_3_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_3_Omuxes_0_0 = MuxesWrapper_3_io_Omuxes_0_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_3_i_mux_bus_0_0_rev_T_2 = {MuxWrapper_3_Omuxes_0_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_3_i_mux_bus_0_0_rev_T_4 = {{1'd0}, MuxWrapper_3_Omuxes_0_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_1968 = {_FDPE_3_i_mux_bus_0_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_3_i_mux_bus_0_0_rev_T_6 = {{1'd0}, _GEN_1968}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_3_i_mux_bus_0_0_rev_T_7 = _FDPE_3_i_mux_bus_0_0_rev_T_2 | _FDPE_3_i_mux_bus_0_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_3_i_mux_bus_0_0_rev_T_8 = {{2'd0}, MuxWrapper_3_Omuxes_0_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_3_i_mux_bus_0_0_rev_T_10 = {_FDPE_3_i_mux_bus_0_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1970 = {{2'd0}, _FDPE_3_i_mux_bus_0_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_3_i_mux_bus_0_0_rev_T_11 = _FDPE_3_i_mux_bus_0_0_rev_T_7 | _GEN_1970; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_3_i_mux_bus_0_0_rev_T_12 = {{3'd0}, MuxWrapper_3_Omuxes_0_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_3_i_mux_bus_0_0_rev_T_14 = {{1'd0}, _FDPE_3_i_mux_bus_0_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1972 = {{2'd0}, _FDPE_3_i_mux_bus_0_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_3_Omuxes_0_1 = MuxesWrapper_3_io_Omuxes_0_1; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_3_i_mux_bus_0_1_rev_T_2 = {MuxWrapper_3_Omuxes_0_1[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_3_i_mux_bus_0_1_rev_T_4 = {{1'd0}, MuxWrapper_3_Omuxes_0_1[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_1974 = {_FDPE_3_i_mux_bus_0_1_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_3_i_mux_bus_0_1_rev_T_6 = {{1'd0}, _GEN_1974}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_3_i_mux_bus_0_1_rev_T_7 = _FDPE_3_i_mux_bus_0_1_rev_T_2 | _FDPE_3_i_mux_bus_0_1_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_3_i_mux_bus_0_1_rev_T_8 = {{2'd0}, MuxWrapper_3_Omuxes_0_1[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_3_i_mux_bus_0_1_rev_T_10 = {_FDPE_3_i_mux_bus_0_1_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1976 = {{2'd0}, _FDPE_3_i_mux_bus_0_1_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_3_i_mux_bus_0_1_rev_T_11 = _FDPE_3_i_mux_bus_0_1_rev_T_7 | _GEN_1976; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_3_i_mux_bus_0_1_rev_T_12 = {{3'd0}, MuxWrapper_3_Omuxes_0_1[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_3_i_mux_bus_0_1_rev_T_14 = {{1'd0}, _FDPE_3_i_mux_bus_0_1_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1978 = {{2'd0}, _FDPE_3_i_mux_bus_0_1_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_3_Omuxes_0_2 = MuxesWrapper_3_io_Omuxes_0_2; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_3_i_mux_bus_0_2_rev_T_2 = {MuxWrapper_3_Omuxes_0_2[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_3_i_mux_bus_0_2_rev_T_4 = {{1'd0}, MuxWrapper_3_Omuxes_0_2[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_1980 = {_FDPE_3_i_mux_bus_0_2_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_3_i_mux_bus_0_2_rev_T_6 = {{1'd0}, _GEN_1980}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_3_i_mux_bus_0_2_rev_T_7 = _FDPE_3_i_mux_bus_0_2_rev_T_2 | _FDPE_3_i_mux_bus_0_2_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_3_i_mux_bus_0_2_rev_T_8 = {{2'd0}, MuxWrapper_3_Omuxes_0_2[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_3_i_mux_bus_0_2_rev_T_10 = {_FDPE_3_i_mux_bus_0_2_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1982 = {{2'd0}, _FDPE_3_i_mux_bus_0_2_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_3_i_mux_bus_0_2_rev_T_11 = _FDPE_3_i_mux_bus_0_2_rev_T_7 | _GEN_1982; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_3_i_mux_bus_0_2_rev_T_12 = {{3'd0}, MuxWrapper_3_Omuxes_0_2[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_3_i_mux_bus_0_2_rev_T_14 = {{1'd0}, _FDPE_3_i_mux_bus_0_2_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1984 = {{2'd0}, _FDPE_3_i_mux_bus_0_2_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_3_Omuxes_0_3 = MuxesWrapper_3_io_Omuxes_0_3; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_3_i_mux_bus_0_3_rev_T_2 = {MuxWrapper_3_Omuxes_0_3[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_3_i_mux_bus_0_3_rev_T_4 = {{1'd0}, MuxWrapper_3_Omuxes_0_3[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_1986 = {_FDPE_3_i_mux_bus_0_3_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_3_i_mux_bus_0_3_rev_T_6 = {{1'd0}, _GEN_1986}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_3_i_mux_bus_0_3_rev_T_7 = _FDPE_3_i_mux_bus_0_3_rev_T_2 | _FDPE_3_i_mux_bus_0_3_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_3_i_mux_bus_0_3_rev_T_8 = {{2'd0}, MuxWrapper_3_Omuxes_0_3[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_3_i_mux_bus_0_3_rev_T_10 = {_FDPE_3_i_mux_bus_0_3_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1988 = {{2'd0}, _FDPE_3_i_mux_bus_0_3_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_3_i_mux_bus_0_3_rev_T_11 = _FDPE_3_i_mux_bus_0_3_rev_T_7 | _GEN_1988; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_3_i_mux_bus_0_3_rev_T_12 = {{3'd0}, MuxWrapper_3_Omuxes_0_3[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_3_i_mux_bus_0_3_rev_T_14 = {{1'd0}, _FDPE_3_i_mux_bus_0_3_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1990 = {{2'd0}, _FDPE_3_i_mux_bus_0_3_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_3_Omuxes_1_0 = MuxesWrapper_3_io_Omuxes_1_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_3_i_mux_bus_1_0_rev_T_2 = {MuxWrapper_3_Omuxes_1_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_3_i_mux_bus_1_0_rev_T_4 = {{1'd0}, MuxWrapper_3_Omuxes_1_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_1992 = {_FDPE_3_i_mux_bus_1_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_3_i_mux_bus_1_0_rev_T_6 = {{1'd0}, _GEN_1992}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_3_i_mux_bus_1_0_rev_T_7 = _FDPE_3_i_mux_bus_1_0_rev_T_2 | _FDPE_3_i_mux_bus_1_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_3_i_mux_bus_1_0_rev_T_8 = {{2'd0}, MuxWrapper_3_Omuxes_1_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_3_i_mux_bus_1_0_rev_T_10 = {_FDPE_3_i_mux_bus_1_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1994 = {{2'd0}, _FDPE_3_i_mux_bus_1_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_3_i_mux_bus_1_0_rev_T_11 = _FDPE_3_i_mux_bus_1_0_rev_T_7 | _GEN_1994; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_3_i_mux_bus_1_0_rev_T_12 = {{3'd0}, MuxWrapper_3_Omuxes_1_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_3_i_mux_bus_1_0_rev_T_14 = {{1'd0}, _FDPE_3_i_mux_bus_1_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_1996 = {{2'd0}, _FDPE_3_i_mux_bus_1_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_3_Omuxes_1_1 = MuxesWrapper_3_io_Omuxes_1_1; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_3_i_mux_bus_1_1_rev_T_2 = {MuxWrapper_3_Omuxes_1_1[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_3_i_mux_bus_1_1_rev_T_4 = {{1'd0}, MuxWrapper_3_Omuxes_1_1[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_1998 = {_FDPE_3_i_mux_bus_1_1_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_3_i_mux_bus_1_1_rev_T_6 = {{1'd0}, _GEN_1998}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_3_i_mux_bus_1_1_rev_T_7 = _FDPE_3_i_mux_bus_1_1_rev_T_2 | _FDPE_3_i_mux_bus_1_1_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_3_i_mux_bus_1_1_rev_T_8 = {{2'd0}, MuxWrapper_3_Omuxes_1_1[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_3_i_mux_bus_1_1_rev_T_10 = {_FDPE_3_i_mux_bus_1_1_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2000 = {{2'd0}, _FDPE_3_i_mux_bus_1_1_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_3_i_mux_bus_1_1_rev_T_11 = _FDPE_3_i_mux_bus_1_1_rev_T_7 | _GEN_2000; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_3_i_mux_bus_1_1_rev_T_12 = {{3'd0}, MuxWrapper_3_Omuxes_1_1[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_3_i_mux_bus_1_1_rev_T_14 = {{1'd0}, _FDPE_3_i_mux_bus_1_1_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2002 = {{2'd0}, _FDPE_3_i_mux_bus_1_1_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_3_Omuxes_1_2 = MuxesWrapper_3_io_Omuxes_1_2; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_3_i_mux_bus_1_2_rev_T_2 = {MuxWrapper_3_Omuxes_1_2[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_3_i_mux_bus_1_2_rev_T_4 = {{1'd0}, MuxWrapper_3_Omuxes_1_2[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2004 = {_FDPE_3_i_mux_bus_1_2_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_3_i_mux_bus_1_2_rev_T_6 = {{1'd0}, _GEN_2004}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_3_i_mux_bus_1_2_rev_T_7 = _FDPE_3_i_mux_bus_1_2_rev_T_2 | _FDPE_3_i_mux_bus_1_2_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_3_i_mux_bus_1_2_rev_T_8 = {{2'd0}, MuxWrapper_3_Omuxes_1_2[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_3_i_mux_bus_1_2_rev_T_10 = {_FDPE_3_i_mux_bus_1_2_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2006 = {{2'd0}, _FDPE_3_i_mux_bus_1_2_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_3_i_mux_bus_1_2_rev_T_11 = _FDPE_3_i_mux_bus_1_2_rev_T_7 | _GEN_2006; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_3_i_mux_bus_1_2_rev_T_12 = {{3'd0}, MuxWrapper_3_Omuxes_1_2[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_3_i_mux_bus_1_2_rev_T_14 = {{1'd0}, _FDPE_3_i_mux_bus_1_2_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2008 = {{2'd0}, _FDPE_3_i_mux_bus_1_2_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_3_Omuxes_2_0 = MuxesWrapper_3_io_Omuxes_2_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_3_i_mux_bus_2_0_rev_T_2 = {MuxWrapper_3_Omuxes_2_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_3_i_mux_bus_2_0_rev_T_4 = {{1'd0}, MuxWrapper_3_Omuxes_2_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2010 = {_FDPE_3_i_mux_bus_2_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_3_i_mux_bus_2_0_rev_T_6 = {{1'd0}, _GEN_2010}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_3_i_mux_bus_2_0_rev_T_7 = _FDPE_3_i_mux_bus_2_0_rev_T_2 | _FDPE_3_i_mux_bus_2_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_3_i_mux_bus_2_0_rev_T_8 = {{2'd0}, MuxWrapper_3_Omuxes_2_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_3_i_mux_bus_2_0_rev_T_10 = {_FDPE_3_i_mux_bus_2_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2012 = {{2'd0}, _FDPE_3_i_mux_bus_2_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_3_i_mux_bus_2_0_rev_T_11 = _FDPE_3_i_mux_bus_2_0_rev_T_7 | _GEN_2012; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_3_i_mux_bus_2_0_rev_T_12 = {{3'd0}, MuxWrapper_3_Omuxes_2_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_3_i_mux_bus_2_0_rev_T_14 = {{1'd0}, _FDPE_3_i_mux_bus_2_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2014 = {{2'd0}, _FDPE_3_i_mux_bus_2_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_3_Omuxes_2_1 = MuxesWrapper_3_io_Omuxes_2_1; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_3_i_mux_bus_2_1_rev_T_2 = {MuxWrapper_3_Omuxes_2_1[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_3_i_mux_bus_2_1_rev_T_4 = {{1'd0}, MuxWrapper_3_Omuxes_2_1[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2016 = {_FDPE_3_i_mux_bus_2_1_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_3_i_mux_bus_2_1_rev_T_6 = {{1'd0}, _GEN_2016}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_3_i_mux_bus_2_1_rev_T_7 = _FDPE_3_i_mux_bus_2_1_rev_T_2 | _FDPE_3_i_mux_bus_2_1_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_3_i_mux_bus_2_1_rev_T_8 = {{2'd0}, MuxWrapper_3_Omuxes_2_1[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_3_i_mux_bus_2_1_rev_T_10 = {_FDPE_3_i_mux_bus_2_1_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2018 = {{2'd0}, _FDPE_3_i_mux_bus_2_1_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_3_i_mux_bus_2_1_rev_T_11 = _FDPE_3_i_mux_bus_2_1_rev_T_7 | _GEN_2018; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_3_i_mux_bus_2_1_rev_T_12 = {{3'd0}, MuxWrapper_3_Omuxes_2_1[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_3_i_mux_bus_2_1_rev_T_14 = {{1'd0}, _FDPE_3_i_mux_bus_2_1_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2020 = {{2'd0}, _FDPE_3_i_mux_bus_2_1_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_3_Omuxes_3_0 = MuxesWrapper_3_io_Omuxes_3_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_3_i_mux_bus_3_0_rev_T_2 = {MuxWrapper_3_Omuxes_3_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_3_i_mux_bus_3_0_rev_T_4 = {{1'd0}, MuxWrapper_3_Omuxes_3_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2022 = {_FDPE_3_i_mux_bus_3_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_3_i_mux_bus_3_0_rev_T_6 = {{1'd0}, _GEN_2022}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_3_i_mux_bus_3_0_rev_T_7 = _FDPE_3_i_mux_bus_3_0_rev_T_2 | _FDPE_3_i_mux_bus_3_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_3_i_mux_bus_3_0_rev_T_8 = {{2'd0}, MuxWrapper_3_Omuxes_3_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_3_i_mux_bus_3_0_rev_T_10 = {_FDPE_3_i_mux_bus_3_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2024 = {{2'd0}, _FDPE_3_i_mux_bus_3_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_3_i_mux_bus_3_0_rev_T_11 = _FDPE_3_i_mux_bus_3_0_rev_T_7 | _GEN_2024; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_3_i_mux_bus_3_0_rev_T_12 = {{3'd0}, MuxWrapper_3_Omuxes_3_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_3_i_mux_bus_3_0_rev_T_14 = {{1'd0}, _FDPE_3_i_mux_bus_3_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2026 = {{2'd0}, _FDPE_3_i_mux_bus_3_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_4_Omuxes_0_0 = MuxesWrapper_4_io_Omuxes_0_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_4_i_mux_bus_0_0_rev_T_2 = {MuxWrapper_4_Omuxes_0_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_4_i_mux_bus_0_0_rev_T_4 = {{1'd0}, MuxWrapper_4_Omuxes_0_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2028 = {_FDPE_4_i_mux_bus_0_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_4_i_mux_bus_0_0_rev_T_6 = {{1'd0}, _GEN_2028}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_4_i_mux_bus_0_0_rev_T_7 = _FDPE_4_i_mux_bus_0_0_rev_T_2 | _FDPE_4_i_mux_bus_0_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_4_i_mux_bus_0_0_rev_T_8 = {{2'd0}, MuxWrapper_4_Omuxes_0_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_4_i_mux_bus_0_0_rev_T_10 = {_FDPE_4_i_mux_bus_0_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2030 = {{2'd0}, _FDPE_4_i_mux_bus_0_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_4_i_mux_bus_0_0_rev_T_11 = _FDPE_4_i_mux_bus_0_0_rev_T_7 | _GEN_2030; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_4_i_mux_bus_0_0_rev_T_12 = {{3'd0}, MuxWrapper_4_Omuxes_0_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_4_i_mux_bus_0_0_rev_T_14 = {{1'd0}, _FDPE_4_i_mux_bus_0_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2032 = {{2'd0}, _FDPE_4_i_mux_bus_0_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_4_Omuxes_0_1 = MuxesWrapper_4_io_Omuxes_0_1; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_4_i_mux_bus_0_1_rev_T_2 = {MuxWrapper_4_Omuxes_0_1[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_4_i_mux_bus_0_1_rev_T_4 = {{1'd0}, MuxWrapper_4_Omuxes_0_1[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2034 = {_FDPE_4_i_mux_bus_0_1_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_4_i_mux_bus_0_1_rev_T_6 = {{1'd0}, _GEN_2034}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_4_i_mux_bus_0_1_rev_T_7 = _FDPE_4_i_mux_bus_0_1_rev_T_2 | _FDPE_4_i_mux_bus_0_1_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_4_i_mux_bus_0_1_rev_T_8 = {{2'd0}, MuxWrapper_4_Omuxes_0_1[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_4_i_mux_bus_0_1_rev_T_10 = {_FDPE_4_i_mux_bus_0_1_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2036 = {{2'd0}, _FDPE_4_i_mux_bus_0_1_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_4_i_mux_bus_0_1_rev_T_11 = _FDPE_4_i_mux_bus_0_1_rev_T_7 | _GEN_2036; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_4_i_mux_bus_0_1_rev_T_12 = {{3'd0}, MuxWrapper_4_Omuxes_0_1[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_4_i_mux_bus_0_1_rev_T_14 = {{1'd0}, _FDPE_4_i_mux_bus_0_1_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2038 = {{2'd0}, _FDPE_4_i_mux_bus_0_1_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_4_Omuxes_0_2 = MuxesWrapper_4_io_Omuxes_0_2; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_4_i_mux_bus_0_2_rev_T_2 = {MuxWrapper_4_Omuxes_0_2[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_4_i_mux_bus_0_2_rev_T_4 = {{1'd0}, MuxWrapper_4_Omuxes_0_2[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2040 = {_FDPE_4_i_mux_bus_0_2_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_4_i_mux_bus_0_2_rev_T_6 = {{1'd0}, _GEN_2040}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_4_i_mux_bus_0_2_rev_T_7 = _FDPE_4_i_mux_bus_0_2_rev_T_2 | _FDPE_4_i_mux_bus_0_2_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_4_i_mux_bus_0_2_rev_T_8 = {{2'd0}, MuxWrapper_4_Omuxes_0_2[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_4_i_mux_bus_0_2_rev_T_10 = {_FDPE_4_i_mux_bus_0_2_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2042 = {{2'd0}, _FDPE_4_i_mux_bus_0_2_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_4_i_mux_bus_0_2_rev_T_11 = _FDPE_4_i_mux_bus_0_2_rev_T_7 | _GEN_2042; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_4_i_mux_bus_0_2_rev_T_12 = {{3'd0}, MuxWrapper_4_Omuxes_0_2[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_4_i_mux_bus_0_2_rev_T_14 = {{1'd0}, _FDPE_4_i_mux_bus_0_2_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2044 = {{2'd0}, _FDPE_4_i_mux_bus_0_2_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_4_Omuxes_0_3 = MuxesWrapper_4_io_Omuxes_0_3; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_4_i_mux_bus_0_3_rev_T_2 = {MuxWrapper_4_Omuxes_0_3[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_4_i_mux_bus_0_3_rev_T_4 = {{1'd0}, MuxWrapper_4_Omuxes_0_3[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2046 = {_FDPE_4_i_mux_bus_0_3_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_4_i_mux_bus_0_3_rev_T_6 = {{1'd0}, _GEN_2046}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_4_i_mux_bus_0_3_rev_T_7 = _FDPE_4_i_mux_bus_0_3_rev_T_2 | _FDPE_4_i_mux_bus_0_3_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_4_i_mux_bus_0_3_rev_T_8 = {{2'd0}, MuxWrapper_4_Omuxes_0_3[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_4_i_mux_bus_0_3_rev_T_10 = {_FDPE_4_i_mux_bus_0_3_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2048 = {{2'd0}, _FDPE_4_i_mux_bus_0_3_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_4_i_mux_bus_0_3_rev_T_11 = _FDPE_4_i_mux_bus_0_3_rev_T_7 | _GEN_2048; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_4_i_mux_bus_0_3_rev_T_12 = {{3'd0}, MuxWrapper_4_Omuxes_0_3[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_4_i_mux_bus_0_3_rev_T_14 = {{1'd0}, _FDPE_4_i_mux_bus_0_3_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2050 = {{2'd0}, _FDPE_4_i_mux_bus_0_3_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_4_Omuxes_1_0 = MuxesWrapper_4_io_Omuxes_1_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_4_i_mux_bus_1_0_rev_T_2 = {MuxWrapper_4_Omuxes_1_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_4_i_mux_bus_1_0_rev_T_4 = {{1'd0}, MuxWrapper_4_Omuxes_1_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2052 = {_FDPE_4_i_mux_bus_1_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_4_i_mux_bus_1_0_rev_T_6 = {{1'd0}, _GEN_2052}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_4_i_mux_bus_1_0_rev_T_7 = _FDPE_4_i_mux_bus_1_0_rev_T_2 | _FDPE_4_i_mux_bus_1_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_4_i_mux_bus_1_0_rev_T_8 = {{2'd0}, MuxWrapper_4_Omuxes_1_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_4_i_mux_bus_1_0_rev_T_10 = {_FDPE_4_i_mux_bus_1_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2054 = {{2'd0}, _FDPE_4_i_mux_bus_1_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_4_i_mux_bus_1_0_rev_T_11 = _FDPE_4_i_mux_bus_1_0_rev_T_7 | _GEN_2054; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_4_i_mux_bus_1_0_rev_T_12 = {{3'd0}, MuxWrapper_4_Omuxes_1_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_4_i_mux_bus_1_0_rev_T_14 = {{1'd0}, _FDPE_4_i_mux_bus_1_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2056 = {{2'd0}, _FDPE_4_i_mux_bus_1_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_4_Omuxes_1_1 = MuxesWrapper_4_io_Omuxes_1_1; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_4_i_mux_bus_1_1_rev_T_2 = {MuxWrapper_4_Omuxes_1_1[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_4_i_mux_bus_1_1_rev_T_4 = {{1'd0}, MuxWrapper_4_Omuxes_1_1[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2058 = {_FDPE_4_i_mux_bus_1_1_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_4_i_mux_bus_1_1_rev_T_6 = {{1'd0}, _GEN_2058}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_4_i_mux_bus_1_1_rev_T_7 = _FDPE_4_i_mux_bus_1_1_rev_T_2 | _FDPE_4_i_mux_bus_1_1_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_4_i_mux_bus_1_1_rev_T_8 = {{2'd0}, MuxWrapper_4_Omuxes_1_1[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_4_i_mux_bus_1_1_rev_T_10 = {_FDPE_4_i_mux_bus_1_1_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2060 = {{2'd0}, _FDPE_4_i_mux_bus_1_1_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_4_i_mux_bus_1_1_rev_T_11 = _FDPE_4_i_mux_bus_1_1_rev_T_7 | _GEN_2060; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_4_i_mux_bus_1_1_rev_T_12 = {{3'd0}, MuxWrapper_4_Omuxes_1_1[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_4_i_mux_bus_1_1_rev_T_14 = {{1'd0}, _FDPE_4_i_mux_bus_1_1_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2062 = {{2'd0}, _FDPE_4_i_mux_bus_1_1_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_4_Omuxes_1_2 = MuxesWrapper_4_io_Omuxes_1_2; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_4_i_mux_bus_1_2_rev_T_2 = {MuxWrapper_4_Omuxes_1_2[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_4_i_mux_bus_1_2_rev_T_4 = {{1'd0}, MuxWrapper_4_Omuxes_1_2[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2064 = {_FDPE_4_i_mux_bus_1_2_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_4_i_mux_bus_1_2_rev_T_6 = {{1'd0}, _GEN_2064}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_4_i_mux_bus_1_2_rev_T_7 = _FDPE_4_i_mux_bus_1_2_rev_T_2 | _FDPE_4_i_mux_bus_1_2_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_4_i_mux_bus_1_2_rev_T_8 = {{2'd0}, MuxWrapper_4_Omuxes_1_2[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_4_i_mux_bus_1_2_rev_T_10 = {_FDPE_4_i_mux_bus_1_2_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2066 = {{2'd0}, _FDPE_4_i_mux_bus_1_2_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_4_i_mux_bus_1_2_rev_T_11 = _FDPE_4_i_mux_bus_1_2_rev_T_7 | _GEN_2066; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_4_i_mux_bus_1_2_rev_T_12 = {{3'd0}, MuxWrapper_4_Omuxes_1_2[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_4_i_mux_bus_1_2_rev_T_14 = {{1'd0}, _FDPE_4_i_mux_bus_1_2_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2068 = {{2'd0}, _FDPE_4_i_mux_bus_1_2_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_4_Omuxes_2_0 = MuxesWrapper_4_io_Omuxes_2_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_4_i_mux_bus_2_0_rev_T_2 = {MuxWrapper_4_Omuxes_2_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_4_i_mux_bus_2_0_rev_T_4 = {{1'd0}, MuxWrapper_4_Omuxes_2_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2070 = {_FDPE_4_i_mux_bus_2_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_4_i_mux_bus_2_0_rev_T_6 = {{1'd0}, _GEN_2070}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_4_i_mux_bus_2_0_rev_T_7 = _FDPE_4_i_mux_bus_2_0_rev_T_2 | _FDPE_4_i_mux_bus_2_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_4_i_mux_bus_2_0_rev_T_8 = {{2'd0}, MuxWrapper_4_Omuxes_2_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_4_i_mux_bus_2_0_rev_T_10 = {_FDPE_4_i_mux_bus_2_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2072 = {{2'd0}, _FDPE_4_i_mux_bus_2_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_4_i_mux_bus_2_0_rev_T_11 = _FDPE_4_i_mux_bus_2_0_rev_T_7 | _GEN_2072; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_4_i_mux_bus_2_0_rev_T_12 = {{3'd0}, MuxWrapper_4_Omuxes_2_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_4_i_mux_bus_2_0_rev_T_14 = {{1'd0}, _FDPE_4_i_mux_bus_2_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2074 = {{2'd0}, _FDPE_4_i_mux_bus_2_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_4_Omuxes_2_1 = MuxesWrapper_4_io_Omuxes_2_1; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_4_i_mux_bus_2_1_rev_T_2 = {MuxWrapper_4_Omuxes_2_1[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_4_i_mux_bus_2_1_rev_T_4 = {{1'd0}, MuxWrapper_4_Omuxes_2_1[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2076 = {_FDPE_4_i_mux_bus_2_1_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_4_i_mux_bus_2_1_rev_T_6 = {{1'd0}, _GEN_2076}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_4_i_mux_bus_2_1_rev_T_7 = _FDPE_4_i_mux_bus_2_1_rev_T_2 | _FDPE_4_i_mux_bus_2_1_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_4_i_mux_bus_2_1_rev_T_8 = {{2'd0}, MuxWrapper_4_Omuxes_2_1[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_4_i_mux_bus_2_1_rev_T_10 = {_FDPE_4_i_mux_bus_2_1_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2078 = {{2'd0}, _FDPE_4_i_mux_bus_2_1_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_4_i_mux_bus_2_1_rev_T_11 = _FDPE_4_i_mux_bus_2_1_rev_T_7 | _GEN_2078; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_4_i_mux_bus_2_1_rev_T_12 = {{3'd0}, MuxWrapper_4_Omuxes_2_1[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_4_i_mux_bus_2_1_rev_T_14 = {{1'd0}, _FDPE_4_i_mux_bus_2_1_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2080 = {{2'd0}, _FDPE_4_i_mux_bus_2_1_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_4_Omuxes_3_0 = MuxesWrapper_4_io_Omuxes_3_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_4_i_mux_bus_3_0_rev_T_2 = {MuxWrapper_4_Omuxes_3_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_4_i_mux_bus_3_0_rev_T_4 = {{1'd0}, MuxWrapper_4_Omuxes_3_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2082 = {_FDPE_4_i_mux_bus_3_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_4_i_mux_bus_3_0_rev_T_6 = {{1'd0}, _GEN_2082}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_4_i_mux_bus_3_0_rev_T_7 = _FDPE_4_i_mux_bus_3_0_rev_T_2 | _FDPE_4_i_mux_bus_3_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_4_i_mux_bus_3_0_rev_T_8 = {{2'd0}, MuxWrapper_4_Omuxes_3_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_4_i_mux_bus_3_0_rev_T_10 = {_FDPE_4_i_mux_bus_3_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2084 = {{2'd0}, _FDPE_4_i_mux_bus_3_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_4_i_mux_bus_3_0_rev_T_11 = _FDPE_4_i_mux_bus_3_0_rev_T_7 | _GEN_2084; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_4_i_mux_bus_3_0_rev_T_12 = {{3'd0}, MuxWrapper_4_Omuxes_3_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_4_i_mux_bus_3_0_rev_T_14 = {{1'd0}, _FDPE_4_i_mux_bus_3_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2086 = {{2'd0}, _FDPE_4_i_mux_bus_3_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_5_Omuxes_0_0 = MuxesWrapper_5_io_Omuxes_0_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_5_i_mux_bus_0_0_rev_T_2 = {MuxWrapper_5_Omuxes_0_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_5_i_mux_bus_0_0_rev_T_4 = {{1'd0}, MuxWrapper_5_Omuxes_0_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2088 = {_FDPE_5_i_mux_bus_0_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_5_i_mux_bus_0_0_rev_T_6 = {{1'd0}, _GEN_2088}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_5_i_mux_bus_0_0_rev_T_7 = _FDPE_5_i_mux_bus_0_0_rev_T_2 | _FDPE_5_i_mux_bus_0_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_5_i_mux_bus_0_0_rev_T_8 = {{2'd0}, MuxWrapper_5_Omuxes_0_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_5_i_mux_bus_0_0_rev_T_10 = {_FDPE_5_i_mux_bus_0_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2090 = {{2'd0}, _FDPE_5_i_mux_bus_0_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_5_i_mux_bus_0_0_rev_T_11 = _FDPE_5_i_mux_bus_0_0_rev_T_7 | _GEN_2090; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_5_i_mux_bus_0_0_rev_T_12 = {{3'd0}, MuxWrapper_5_Omuxes_0_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_5_i_mux_bus_0_0_rev_T_14 = {{1'd0}, _FDPE_5_i_mux_bus_0_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2092 = {{2'd0}, _FDPE_5_i_mux_bus_0_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_5_Omuxes_0_1 = MuxesWrapper_5_io_Omuxes_0_1; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_5_i_mux_bus_0_1_rev_T_2 = {MuxWrapper_5_Omuxes_0_1[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_5_i_mux_bus_0_1_rev_T_4 = {{1'd0}, MuxWrapper_5_Omuxes_0_1[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2094 = {_FDPE_5_i_mux_bus_0_1_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_5_i_mux_bus_0_1_rev_T_6 = {{1'd0}, _GEN_2094}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_5_i_mux_bus_0_1_rev_T_7 = _FDPE_5_i_mux_bus_0_1_rev_T_2 | _FDPE_5_i_mux_bus_0_1_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_5_i_mux_bus_0_1_rev_T_8 = {{2'd0}, MuxWrapper_5_Omuxes_0_1[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_5_i_mux_bus_0_1_rev_T_10 = {_FDPE_5_i_mux_bus_0_1_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2096 = {{2'd0}, _FDPE_5_i_mux_bus_0_1_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_5_i_mux_bus_0_1_rev_T_11 = _FDPE_5_i_mux_bus_0_1_rev_T_7 | _GEN_2096; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_5_i_mux_bus_0_1_rev_T_12 = {{3'd0}, MuxWrapper_5_Omuxes_0_1[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_5_i_mux_bus_0_1_rev_T_14 = {{1'd0}, _FDPE_5_i_mux_bus_0_1_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2098 = {{2'd0}, _FDPE_5_i_mux_bus_0_1_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_5_Omuxes_0_2 = MuxesWrapper_5_io_Omuxes_0_2; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_5_i_mux_bus_0_2_rev_T_2 = {MuxWrapper_5_Omuxes_0_2[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_5_i_mux_bus_0_2_rev_T_4 = {{1'd0}, MuxWrapper_5_Omuxes_0_2[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2100 = {_FDPE_5_i_mux_bus_0_2_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_5_i_mux_bus_0_2_rev_T_6 = {{1'd0}, _GEN_2100}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_5_i_mux_bus_0_2_rev_T_7 = _FDPE_5_i_mux_bus_0_2_rev_T_2 | _FDPE_5_i_mux_bus_0_2_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_5_i_mux_bus_0_2_rev_T_8 = {{2'd0}, MuxWrapper_5_Omuxes_0_2[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_5_i_mux_bus_0_2_rev_T_10 = {_FDPE_5_i_mux_bus_0_2_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2102 = {{2'd0}, _FDPE_5_i_mux_bus_0_2_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_5_i_mux_bus_0_2_rev_T_11 = _FDPE_5_i_mux_bus_0_2_rev_T_7 | _GEN_2102; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_5_i_mux_bus_0_2_rev_T_12 = {{3'd0}, MuxWrapper_5_Omuxes_0_2[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_5_i_mux_bus_0_2_rev_T_14 = {{1'd0}, _FDPE_5_i_mux_bus_0_2_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2104 = {{2'd0}, _FDPE_5_i_mux_bus_0_2_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_5_Omuxes_0_3 = MuxesWrapper_5_io_Omuxes_0_3; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_5_i_mux_bus_0_3_rev_T_2 = {MuxWrapper_5_Omuxes_0_3[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_5_i_mux_bus_0_3_rev_T_4 = {{1'd0}, MuxWrapper_5_Omuxes_0_3[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2106 = {_FDPE_5_i_mux_bus_0_3_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_5_i_mux_bus_0_3_rev_T_6 = {{1'd0}, _GEN_2106}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_5_i_mux_bus_0_3_rev_T_7 = _FDPE_5_i_mux_bus_0_3_rev_T_2 | _FDPE_5_i_mux_bus_0_3_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_5_i_mux_bus_0_3_rev_T_8 = {{2'd0}, MuxWrapper_5_Omuxes_0_3[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_5_i_mux_bus_0_3_rev_T_10 = {_FDPE_5_i_mux_bus_0_3_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2108 = {{2'd0}, _FDPE_5_i_mux_bus_0_3_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_5_i_mux_bus_0_3_rev_T_11 = _FDPE_5_i_mux_bus_0_3_rev_T_7 | _GEN_2108; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_5_i_mux_bus_0_3_rev_T_12 = {{3'd0}, MuxWrapper_5_Omuxes_0_3[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_5_i_mux_bus_0_3_rev_T_14 = {{1'd0}, _FDPE_5_i_mux_bus_0_3_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2110 = {{2'd0}, _FDPE_5_i_mux_bus_0_3_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_5_Omuxes_1_0 = MuxesWrapper_5_io_Omuxes_1_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_5_i_mux_bus_1_0_rev_T_2 = {MuxWrapper_5_Omuxes_1_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_5_i_mux_bus_1_0_rev_T_4 = {{1'd0}, MuxWrapper_5_Omuxes_1_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2112 = {_FDPE_5_i_mux_bus_1_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_5_i_mux_bus_1_0_rev_T_6 = {{1'd0}, _GEN_2112}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_5_i_mux_bus_1_0_rev_T_7 = _FDPE_5_i_mux_bus_1_0_rev_T_2 | _FDPE_5_i_mux_bus_1_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_5_i_mux_bus_1_0_rev_T_8 = {{2'd0}, MuxWrapper_5_Omuxes_1_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_5_i_mux_bus_1_0_rev_T_10 = {_FDPE_5_i_mux_bus_1_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2114 = {{2'd0}, _FDPE_5_i_mux_bus_1_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_5_i_mux_bus_1_0_rev_T_11 = _FDPE_5_i_mux_bus_1_0_rev_T_7 | _GEN_2114; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_5_i_mux_bus_1_0_rev_T_12 = {{3'd0}, MuxWrapper_5_Omuxes_1_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_5_i_mux_bus_1_0_rev_T_14 = {{1'd0}, _FDPE_5_i_mux_bus_1_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2116 = {{2'd0}, _FDPE_5_i_mux_bus_1_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_5_Omuxes_1_1 = MuxesWrapper_5_io_Omuxes_1_1; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_5_i_mux_bus_1_1_rev_T_2 = {MuxWrapper_5_Omuxes_1_1[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_5_i_mux_bus_1_1_rev_T_4 = {{1'd0}, MuxWrapper_5_Omuxes_1_1[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2118 = {_FDPE_5_i_mux_bus_1_1_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_5_i_mux_bus_1_1_rev_T_6 = {{1'd0}, _GEN_2118}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_5_i_mux_bus_1_1_rev_T_7 = _FDPE_5_i_mux_bus_1_1_rev_T_2 | _FDPE_5_i_mux_bus_1_1_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_5_i_mux_bus_1_1_rev_T_8 = {{2'd0}, MuxWrapper_5_Omuxes_1_1[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_5_i_mux_bus_1_1_rev_T_10 = {_FDPE_5_i_mux_bus_1_1_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2120 = {{2'd0}, _FDPE_5_i_mux_bus_1_1_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_5_i_mux_bus_1_1_rev_T_11 = _FDPE_5_i_mux_bus_1_1_rev_T_7 | _GEN_2120; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_5_i_mux_bus_1_1_rev_T_12 = {{3'd0}, MuxWrapper_5_Omuxes_1_1[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_5_i_mux_bus_1_1_rev_T_14 = {{1'd0}, _FDPE_5_i_mux_bus_1_1_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2122 = {{2'd0}, _FDPE_5_i_mux_bus_1_1_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_5_Omuxes_1_2 = MuxesWrapper_5_io_Omuxes_1_2; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_5_i_mux_bus_1_2_rev_T_2 = {MuxWrapper_5_Omuxes_1_2[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_5_i_mux_bus_1_2_rev_T_4 = {{1'd0}, MuxWrapper_5_Omuxes_1_2[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2124 = {_FDPE_5_i_mux_bus_1_2_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_5_i_mux_bus_1_2_rev_T_6 = {{1'd0}, _GEN_2124}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_5_i_mux_bus_1_2_rev_T_7 = _FDPE_5_i_mux_bus_1_2_rev_T_2 | _FDPE_5_i_mux_bus_1_2_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_5_i_mux_bus_1_2_rev_T_8 = {{2'd0}, MuxWrapper_5_Omuxes_1_2[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_5_i_mux_bus_1_2_rev_T_10 = {_FDPE_5_i_mux_bus_1_2_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2126 = {{2'd0}, _FDPE_5_i_mux_bus_1_2_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_5_i_mux_bus_1_2_rev_T_11 = _FDPE_5_i_mux_bus_1_2_rev_T_7 | _GEN_2126; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_5_i_mux_bus_1_2_rev_T_12 = {{3'd0}, MuxWrapper_5_Omuxes_1_2[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_5_i_mux_bus_1_2_rev_T_14 = {{1'd0}, _FDPE_5_i_mux_bus_1_2_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2128 = {{2'd0}, _FDPE_5_i_mux_bus_1_2_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_5_Omuxes_2_0 = MuxesWrapper_5_io_Omuxes_2_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_5_i_mux_bus_2_0_rev_T_2 = {MuxWrapper_5_Omuxes_2_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_5_i_mux_bus_2_0_rev_T_4 = {{1'd0}, MuxWrapper_5_Omuxes_2_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2130 = {_FDPE_5_i_mux_bus_2_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_5_i_mux_bus_2_0_rev_T_6 = {{1'd0}, _GEN_2130}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_5_i_mux_bus_2_0_rev_T_7 = _FDPE_5_i_mux_bus_2_0_rev_T_2 | _FDPE_5_i_mux_bus_2_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_5_i_mux_bus_2_0_rev_T_8 = {{2'd0}, MuxWrapper_5_Omuxes_2_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_5_i_mux_bus_2_0_rev_T_10 = {_FDPE_5_i_mux_bus_2_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2132 = {{2'd0}, _FDPE_5_i_mux_bus_2_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_5_i_mux_bus_2_0_rev_T_11 = _FDPE_5_i_mux_bus_2_0_rev_T_7 | _GEN_2132; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_5_i_mux_bus_2_0_rev_T_12 = {{3'd0}, MuxWrapper_5_Omuxes_2_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_5_i_mux_bus_2_0_rev_T_14 = {{1'd0}, _FDPE_5_i_mux_bus_2_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2134 = {{2'd0}, _FDPE_5_i_mux_bus_2_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_5_Omuxes_2_1 = MuxesWrapper_5_io_Omuxes_2_1; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_5_i_mux_bus_2_1_rev_T_2 = {MuxWrapper_5_Omuxes_2_1[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_5_i_mux_bus_2_1_rev_T_4 = {{1'd0}, MuxWrapper_5_Omuxes_2_1[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2136 = {_FDPE_5_i_mux_bus_2_1_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_5_i_mux_bus_2_1_rev_T_6 = {{1'd0}, _GEN_2136}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_5_i_mux_bus_2_1_rev_T_7 = _FDPE_5_i_mux_bus_2_1_rev_T_2 | _FDPE_5_i_mux_bus_2_1_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_5_i_mux_bus_2_1_rev_T_8 = {{2'd0}, MuxWrapper_5_Omuxes_2_1[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_5_i_mux_bus_2_1_rev_T_10 = {_FDPE_5_i_mux_bus_2_1_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2138 = {{2'd0}, _FDPE_5_i_mux_bus_2_1_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_5_i_mux_bus_2_1_rev_T_11 = _FDPE_5_i_mux_bus_2_1_rev_T_7 | _GEN_2138; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_5_i_mux_bus_2_1_rev_T_12 = {{3'd0}, MuxWrapper_5_Omuxes_2_1[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_5_i_mux_bus_2_1_rev_T_14 = {{1'd0}, _FDPE_5_i_mux_bus_2_1_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2140 = {{2'd0}, _FDPE_5_i_mux_bus_2_1_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_5_Omuxes_3_0 = MuxesWrapper_5_io_Omuxes_3_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_5_i_mux_bus_3_0_rev_T_2 = {MuxWrapper_5_Omuxes_3_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_5_i_mux_bus_3_0_rev_T_4 = {{1'd0}, MuxWrapper_5_Omuxes_3_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2142 = {_FDPE_5_i_mux_bus_3_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_5_i_mux_bus_3_0_rev_T_6 = {{1'd0}, _GEN_2142}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_5_i_mux_bus_3_0_rev_T_7 = _FDPE_5_i_mux_bus_3_0_rev_T_2 | _FDPE_5_i_mux_bus_3_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_5_i_mux_bus_3_0_rev_T_8 = {{2'd0}, MuxWrapper_5_Omuxes_3_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_5_i_mux_bus_3_0_rev_T_10 = {_FDPE_5_i_mux_bus_3_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2144 = {{2'd0}, _FDPE_5_i_mux_bus_3_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_5_i_mux_bus_3_0_rev_T_11 = _FDPE_5_i_mux_bus_3_0_rev_T_7 | _GEN_2144; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_5_i_mux_bus_3_0_rev_T_12 = {{3'd0}, MuxWrapper_5_Omuxes_3_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_5_i_mux_bus_3_0_rev_T_14 = {{1'd0}, _FDPE_5_i_mux_bus_3_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2146 = {{2'd0}, _FDPE_5_i_mux_bus_3_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_6_Omuxes_0_0 = MuxesWrapper_6_io_Omuxes_0_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_6_i_mux_bus_0_0_rev_T_2 = {MuxWrapper_6_Omuxes_0_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_6_i_mux_bus_0_0_rev_T_4 = {{1'd0}, MuxWrapper_6_Omuxes_0_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2148 = {_FDPE_6_i_mux_bus_0_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_6_i_mux_bus_0_0_rev_T_6 = {{1'd0}, _GEN_2148}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_6_i_mux_bus_0_0_rev_T_7 = _FDPE_6_i_mux_bus_0_0_rev_T_2 | _FDPE_6_i_mux_bus_0_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_6_i_mux_bus_0_0_rev_T_8 = {{2'd0}, MuxWrapper_6_Omuxes_0_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_6_i_mux_bus_0_0_rev_T_10 = {_FDPE_6_i_mux_bus_0_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2150 = {{2'd0}, _FDPE_6_i_mux_bus_0_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_6_i_mux_bus_0_0_rev_T_11 = _FDPE_6_i_mux_bus_0_0_rev_T_7 | _GEN_2150; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_6_i_mux_bus_0_0_rev_T_12 = {{3'd0}, MuxWrapper_6_Omuxes_0_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_6_i_mux_bus_0_0_rev_T_14 = {{1'd0}, _FDPE_6_i_mux_bus_0_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2152 = {{2'd0}, _FDPE_6_i_mux_bus_0_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_6_Omuxes_0_1 = MuxesWrapper_6_io_Omuxes_0_1; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_6_i_mux_bus_0_1_rev_T_2 = {MuxWrapper_6_Omuxes_0_1[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_6_i_mux_bus_0_1_rev_T_4 = {{1'd0}, MuxWrapper_6_Omuxes_0_1[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2154 = {_FDPE_6_i_mux_bus_0_1_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_6_i_mux_bus_0_1_rev_T_6 = {{1'd0}, _GEN_2154}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_6_i_mux_bus_0_1_rev_T_7 = _FDPE_6_i_mux_bus_0_1_rev_T_2 | _FDPE_6_i_mux_bus_0_1_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_6_i_mux_bus_0_1_rev_T_8 = {{2'd0}, MuxWrapper_6_Omuxes_0_1[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_6_i_mux_bus_0_1_rev_T_10 = {_FDPE_6_i_mux_bus_0_1_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2156 = {{2'd0}, _FDPE_6_i_mux_bus_0_1_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_6_i_mux_bus_0_1_rev_T_11 = _FDPE_6_i_mux_bus_0_1_rev_T_7 | _GEN_2156; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_6_i_mux_bus_0_1_rev_T_12 = {{3'd0}, MuxWrapper_6_Omuxes_0_1[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_6_i_mux_bus_0_1_rev_T_14 = {{1'd0}, _FDPE_6_i_mux_bus_0_1_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2158 = {{2'd0}, _FDPE_6_i_mux_bus_0_1_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_6_Omuxes_0_2 = MuxesWrapper_6_io_Omuxes_0_2; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_6_i_mux_bus_0_2_rev_T_2 = {MuxWrapper_6_Omuxes_0_2[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_6_i_mux_bus_0_2_rev_T_4 = {{1'd0}, MuxWrapper_6_Omuxes_0_2[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2160 = {_FDPE_6_i_mux_bus_0_2_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_6_i_mux_bus_0_2_rev_T_6 = {{1'd0}, _GEN_2160}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_6_i_mux_bus_0_2_rev_T_7 = _FDPE_6_i_mux_bus_0_2_rev_T_2 | _FDPE_6_i_mux_bus_0_2_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_6_i_mux_bus_0_2_rev_T_8 = {{2'd0}, MuxWrapper_6_Omuxes_0_2[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_6_i_mux_bus_0_2_rev_T_10 = {_FDPE_6_i_mux_bus_0_2_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2162 = {{2'd0}, _FDPE_6_i_mux_bus_0_2_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_6_i_mux_bus_0_2_rev_T_11 = _FDPE_6_i_mux_bus_0_2_rev_T_7 | _GEN_2162; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_6_i_mux_bus_0_2_rev_T_12 = {{3'd0}, MuxWrapper_6_Omuxes_0_2[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_6_i_mux_bus_0_2_rev_T_14 = {{1'd0}, _FDPE_6_i_mux_bus_0_2_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2164 = {{2'd0}, _FDPE_6_i_mux_bus_0_2_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_6_Omuxes_0_3 = MuxesWrapper_6_io_Omuxes_0_3; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_6_i_mux_bus_0_3_rev_T_2 = {MuxWrapper_6_Omuxes_0_3[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_6_i_mux_bus_0_3_rev_T_4 = {{1'd0}, MuxWrapper_6_Omuxes_0_3[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2166 = {_FDPE_6_i_mux_bus_0_3_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_6_i_mux_bus_0_3_rev_T_6 = {{1'd0}, _GEN_2166}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_6_i_mux_bus_0_3_rev_T_7 = _FDPE_6_i_mux_bus_0_3_rev_T_2 | _FDPE_6_i_mux_bus_0_3_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_6_i_mux_bus_0_3_rev_T_8 = {{2'd0}, MuxWrapper_6_Omuxes_0_3[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_6_i_mux_bus_0_3_rev_T_10 = {_FDPE_6_i_mux_bus_0_3_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2168 = {{2'd0}, _FDPE_6_i_mux_bus_0_3_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_6_i_mux_bus_0_3_rev_T_11 = _FDPE_6_i_mux_bus_0_3_rev_T_7 | _GEN_2168; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_6_i_mux_bus_0_3_rev_T_12 = {{3'd0}, MuxWrapper_6_Omuxes_0_3[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_6_i_mux_bus_0_3_rev_T_14 = {{1'd0}, _FDPE_6_i_mux_bus_0_3_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2170 = {{2'd0}, _FDPE_6_i_mux_bus_0_3_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_6_Omuxes_1_0 = MuxesWrapper_6_io_Omuxes_1_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_6_i_mux_bus_1_0_rev_T_2 = {MuxWrapper_6_Omuxes_1_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_6_i_mux_bus_1_0_rev_T_4 = {{1'd0}, MuxWrapper_6_Omuxes_1_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2172 = {_FDPE_6_i_mux_bus_1_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_6_i_mux_bus_1_0_rev_T_6 = {{1'd0}, _GEN_2172}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_6_i_mux_bus_1_0_rev_T_7 = _FDPE_6_i_mux_bus_1_0_rev_T_2 | _FDPE_6_i_mux_bus_1_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_6_i_mux_bus_1_0_rev_T_8 = {{2'd0}, MuxWrapper_6_Omuxes_1_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_6_i_mux_bus_1_0_rev_T_10 = {_FDPE_6_i_mux_bus_1_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2174 = {{2'd0}, _FDPE_6_i_mux_bus_1_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_6_i_mux_bus_1_0_rev_T_11 = _FDPE_6_i_mux_bus_1_0_rev_T_7 | _GEN_2174; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_6_i_mux_bus_1_0_rev_T_12 = {{3'd0}, MuxWrapper_6_Omuxes_1_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_6_i_mux_bus_1_0_rev_T_14 = {{1'd0}, _FDPE_6_i_mux_bus_1_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2176 = {{2'd0}, _FDPE_6_i_mux_bus_1_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_6_Omuxes_1_1 = MuxesWrapper_6_io_Omuxes_1_1; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_6_i_mux_bus_1_1_rev_T_2 = {MuxWrapper_6_Omuxes_1_1[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_6_i_mux_bus_1_1_rev_T_4 = {{1'd0}, MuxWrapper_6_Omuxes_1_1[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2178 = {_FDPE_6_i_mux_bus_1_1_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_6_i_mux_bus_1_1_rev_T_6 = {{1'd0}, _GEN_2178}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_6_i_mux_bus_1_1_rev_T_7 = _FDPE_6_i_mux_bus_1_1_rev_T_2 | _FDPE_6_i_mux_bus_1_1_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_6_i_mux_bus_1_1_rev_T_8 = {{2'd0}, MuxWrapper_6_Omuxes_1_1[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_6_i_mux_bus_1_1_rev_T_10 = {_FDPE_6_i_mux_bus_1_1_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2180 = {{2'd0}, _FDPE_6_i_mux_bus_1_1_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_6_i_mux_bus_1_1_rev_T_11 = _FDPE_6_i_mux_bus_1_1_rev_T_7 | _GEN_2180; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_6_i_mux_bus_1_1_rev_T_12 = {{3'd0}, MuxWrapper_6_Omuxes_1_1[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_6_i_mux_bus_1_1_rev_T_14 = {{1'd0}, _FDPE_6_i_mux_bus_1_1_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2182 = {{2'd0}, _FDPE_6_i_mux_bus_1_1_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_6_Omuxes_1_2 = MuxesWrapper_6_io_Omuxes_1_2; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_6_i_mux_bus_1_2_rev_T_2 = {MuxWrapper_6_Omuxes_1_2[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_6_i_mux_bus_1_2_rev_T_4 = {{1'd0}, MuxWrapper_6_Omuxes_1_2[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2184 = {_FDPE_6_i_mux_bus_1_2_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_6_i_mux_bus_1_2_rev_T_6 = {{1'd0}, _GEN_2184}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_6_i_mux_bus_1_2_rev_T_7 = _FDPE_6_i_mux_bus_1_2_rev_T_2 | _FDPE_6_i_mux_bus_1_2_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_6_i_mux_bus_1_2_rev_T_8 = {{2'd0}, MuxWrapper_6_Omuxes_1_2[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_6_i_mux_bus_1_2_rev_T_10 = {_FDPE_6_i_mux_bus_1_2_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2186 = {{2'd0}, _FDPE_6_i_mux_bus_1_2_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_6_i_mux_bus_1_2_rev_T_11 = _FDPE_6_i_mux_bus_1_2_rev_T_7 | _GEN_2186; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_6_i_mux_bus_1_2_rev_T_12 = {{3'd0}, MuxWrapper_6_Omuxes_1_2[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_6_i_mux_bus_1_2_rev_T_14 = {{1'd0}, _FDPE_6_i_mux_bus_1_2_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2188 = {{2'd0}, _FDPE_6_i_mux_bus_1_2_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_6_Omuxes_2_0 = MuxesWrapper_6_io_Omuxes_2_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_6_i_mux_bus_2_0_rev_T_2 = {MuxWrapper_6_Omuxes_2_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_6_i_mux_bus_2_0_rev_T_4 = {{1'd0}, MuxWrapper_6_Omuxes_2_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2190 = {_FDPE_6_i_mux_bus_2_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_6_i_mux_bus_2_0_rev_T_6 = {{1'd0}, _GEN_2190}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_6_i_mux_bus_2_0_rev_T_7 = _FDPE_6_i_mux_bus_2_0_rev_T_2 | _FDPE_6_i_mux_bus_2_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_6_i_mux_bus_2_0_rev_T_8 = {{2'd0}, MuxWrapper_6_Omuxes_2_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_6_i_mux_bus_2_0_rev_T_10 = {_FDPE_6_i_mux_bus_2_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2192 = {{2'd0}, _FDPE_6_i_mux_bus_2_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_6_i_mux_bus_2_0_rev_T_11 = _FDPE_6_i_mux_bus_2_0_rev_T_7 | _GEN_2192; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_6_i_mux_bus_2_0_rev_T_12 = {{3'd0}, MuxWrapper_6_Omuxes_2_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_6_i_mux_bus_2_0_rev_T_14 = {{1'd0}, _FDPE_6_i_mux_bus_2_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2194 = {{2'd0}, _FDPE_6_i_mux_bus_2_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_6_Omuxes_2_1 = MuxesWrapper_6_io_Omuxes_2_1; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_6_i_mux_bus_2_1_rev_T_2 = {MuxWrapper_6_Omuxes_2_1[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_6_i_mux_bus_2_1_rev_T_4 = {{1'd0}, MuxWrapper_6_Omuxes_2_1[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2196 = {_FDPE_6_i_mux_bus_2_1_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_6_i_mux_bus_2_1_rev_T_6 = {{1'd0}, _GEN_2196}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_6_i_mux_bus_2_1_rev_T_7 = _FDPE_6_i_mux_bus_2_1_rev_T_2 | _FDPE_6_i_mux_bus_2_1_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_6_i_mux_bus_2_1_rev_T_8 = {{2'd0}, MuxWrapper_6_Omuxes_2_1[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_6_i_mux_bus_2_1_rev_T_10 = {_FDPE_6_i_mux_bus_2_1_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2198 = {{2'd0}, _FDPE_6_i_mux_bus_2_1_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_6_i_mux_bus_2_1_rev_T_11 = _FDPE_6_i_mux_bus_2_1_rev_T_7 | _GEN_2198; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_6_i_mux_bus_2_1_rev_T_12 = {{3'd0}, MuxWrapper_6_Omuxes_2_1[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_6_i_mux_bus_2_1_rev_T_14 = {{1'd0}, _FDPE_6_i_mux_bus_2_1_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2200 = {{2'd0}, _FDPE_6_i_mux_bus_2_1_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_6_Omuxes_3_0 = MuxesWrapper_6_io_Omuxes_3_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_6_i_mux_bus_3_0_rev_T_2 = {MuxWrapper_6_Omuxes_3_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_6_i_mux_bus_3_0_rev_T_4 = {{1'd0}, MuxWrapper_6_Omuxes_3_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2202 = {_FDPE_6_i_mux_bus_3_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_6_i_mux_bus_3_0_rev_T_6 = {{1'd0}, _GEN_2202}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_6_i_mux_bus_3_0_rev_T_7 = _FDPE_6_i_mux_bus_3_0_rev_T_2 | _FDPE_6_i_mux_bus_3_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_6_i_mux_bus_3_0_rev_T_8 = {{2'd0}, MuxWrapper_6_Omuxes_3_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_6_i_mux_bus_3_0_rev_T_10 = {_FDPE_6_i_mux_bus_3_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2204 = {{2'd0}, _FDPE_6_i_mux_bus_3_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_6_i_mux_bus_3_0_rev_T_11 = _FDPE_6_i_mux_bus_3_0_rev_T_7 | _GEN_2204; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_6_i_mux_bus_3_0_rev_T_12 = {{3'd0}, MuxWrapper_6_Omuxes_3_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_6_i_mux_bus_3_0_rev_T_14 = {{1'd0}, _FDPE_6_i_mux_bus_3_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2206 = {{2'd0}, _FDPE_6_i_mux_bus_3_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_7_Omuxes_0_0 = MuxesWrapper_7_io_Omuxes_0_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_7_i_mux_bus_0_0_rev_T_2 = {MuxWrapper_7_Omuxes_0_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_7_i_mux_bus_0_0_rev_T_4 = {{1'd0}, MuxWrapper_7_Omuxes_0_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2208 = {_FDPE_7_i_mux_bus_0_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_7_i_mux_bus_0_0_rev_T_6 = {{1'd0}, _GEN_2208}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_7_i_mux_bus_0_0_rev_T_7 = _FDPE_7_i_mux_bus_0_0_rev_T_2 | _FDPE_7_i_mux_bus_0_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_7_i_mux_bus_0_0_rev_T_8 = {{2'd0}, MuxWrapper_7_Omuxes_0_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_7_i_mux_bus_0_0_rev_T_10 = {_FDPE_7_i_mux_bus_0_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2210 = {{2'd0}, _FDPE_7_i_mux_bus_0_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_7_i_mux_bus_0_0_rev_T_11 = _FDPE_7_i_mux_bus_0_0_rev_T_7 | _GEN_2210; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_7_i_mux_bus_0_0_rev_T_12 = {{3'd0}, MuxWrapper_7_Omuxes_0_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_7_i_mux_bus_0_0_rev_T_14 = {{1'd0}, _FDPE_7_i_mux_bus_0_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2212 = {{2'd0}, _FDPE_7_i_mux_bus_0_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_7_Omuxes_0_1 = MuxesWrapper_7_io_Omuxes_0_1; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_7_i_mux_bus_0_1_rev_T_2 = {MuxWrapper_7_Omuxes_0_1[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_7_i_mux_bus_0_1_rev_T_4 = {{1'd0}, MuxWrapper_7_Omuxes_0_1[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2214 = {_FDPE_7_i_mux_bus_0_1_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_7_i_mux_bus_0_1_rev_T_6 = {{1'd0}, _GEN_2214}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_7_i_mux_bus_0_1_rev_T_7 = _FDPE_7_i_mux_bus_0_1_rev_T_2 | _FDPE_7_i_mux_bus_0_1_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_7_i_mux_bus_0_1_rev_T_8 = {{2'd0}, MuxWrapper_7_Omuxes_0_1[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_7_i_mux_bus_0_1_rev_T_10 = {_FDPE_7_i_mux_bus_0_1_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2216 = {{2'd0}, _FDPE_7_i_mux_bus_0_1_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_7_i_mux_bus_0_1_rev_T_11 = _FDPE_7_i_mux_bus_0_1_rev_T_7 | _GEN_2216; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_7_i_mux_bus_0_1_rev_T_12 = {{3'd0}, MuxWrapper_7_Omuxes_0_1[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_7_i_mux_bus_0_1_rev_T_14 = {{1'd0}, _FDPE_7_i_mux_bus_0_1_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2218 = {{2'd0}, _FDPE_7_i_mux_bus_0_1_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_7_Omuxes_0_2 = MuxesWrapper_7_io_Omuxes_0_2; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_7_i_mux_bus_0_2_rev_T_2 = {MuxWrapper_7_Omuxes_0_2[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_7_i_mux_bus_0_2_rev_T_4 = {{1'd0}, MuxWrapper_7_Omuxes_0_2[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2220 = {_FDPE_7_i_mux_bus_0_2_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_7_i_mux_bus_0_2_rev_T_6 = {{1'd0}, _GEN_2220}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_7_i_mux_bus_0_2_rev_T_7 = _FDPE_7_i_mux_bus_0_2_rev_T_2 | _FDPE_7_i_mux_bus_0_2_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_7_i_mux_bus_0_2_rev_T_8 = {{2'd0}, MuxWrapper_7_Omuxes_0_2[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_7_i_mux_bus_0_2_rev_T_10 = {_FDPE_7_i_mux_bus_0_2_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2222 = {{2'd0}, _FDPE_7_i_mux_bus_0_2_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_7_i_mux_bus_0_2_rev_T_11 = _FDPE_7_i_mux_bus_0_2_rev_T_7 | _GEN_2222; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_7_i_mux_bus_0_2_rev_T_12 = {{3'd0}, MuxWrapper_7_Omuxes_0_2[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_7_i_mux_bus_0_2_rev_T_14 = {{1'd0}, _FDPE_7_i_mux_bus_0_2_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2224 = {{2'd0}, _FDPE_7_i_mux_bus_0_2_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_7_Omuxes_0_3 = MuxesWrapper_7_io_Omuxes_0_3; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_7_i_mux_bus_0_3_rev_T_2 = {MuxWrapper_7_Omuxes_0_3[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_7_i_mux_bus_0_3_rev_T_4 = {{1'd0}, MuxWrapper_7_Omuxes_0_3[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2226 = {_FDPE_7_i_mux_bus_0_3_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_7_i_mux_bus_0_3_rev_T_6 = {{1'd0}, _GEN_2226}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_7_i_mux_bus_0_3_rev_T_7 = _FDPE_7_i_mux_bus_0_3_rev_T_2 | _FDPE_7_i_mux_bus_0_3_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_7_i_mux_bus_0_3_rev_T_8 = {{2'd0}, MuxWrapper_7_Omuxes_0_3[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_7_i_mux_bus_0_3_rev_T_10 = {_FDPE_7_i_mux_bus_0_3_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2228 = {{2'd0}, _FDPE_7_i_mux_bus_0_3_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_7_i_mux_bus_0_3_rev_T_11 = _FDPE_7_i_mux_bus_0_3_rev_T_7 | _GEN_2228; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_7_i_mux_bus_0_3_rev_T_12 = {{3'd0}, MuxWrapper_7_Omuxes_0_3[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_7_i_mux_bus_0_3_rev_T_14 = {{1'd0}, _FDPE_7_i_mux_bus_0_3_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2230 = {{2'd0}, _FDPE_7_i_mux_bus_0_3_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_7_Omuxes_1_0 = MuxesWrapper_7_io_Omuxes_1_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_7_i_mux_bus_1_0_rev_T_2 = {MuxWrapper_7_Omuxes_1_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_7_i_mux_bus_1_0_rev_T_4 = {{1'd0}, MuxWrapper_7_Omuxes_1_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2232 = {_FDPE_7_i_mux_bus_1_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_7_i_mux_bus_1_0_rev_T_6 = {{1'd0}, _GEN_2232}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_7_i_mux_bus_1_0_rev_T_7 = _FDPE_7_i_mux_bus_1_0_rev_T_2 | _FDPE_7_i_mux_bus_1_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_7_i_mux_bus_1_0_rev_T_8 = {{2'd0}, MuxWrapper_7_Omuxes_1_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_7_i_mux_bus_1_0_rev_T_10 = {_FDPE_7_i_mux_bus_1_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2234 = {{2'd0}, _FDPE_7_i_mux_bus_1_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_7_i_mux_bus_1_0_rev_T_11 = _FDPE_7_i_mux_bus_1_0_rev_T_7 | _GEN_2234; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_7_i_mux_bus_1_0_rev_T_12 = {{3'd0}, MuxWrapper_7_Omuxes_1_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_7_i_mux_bus_1_0_rev_T_14 = {{1'd0}, _FDPE_7_i_mux_bus_1_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2236 = {{2'd0}, _FDPE_7_i_mux_bus_1_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_7_Omuxes_1_1 = MuxesWrapper_7_io_Omuxes_1_1; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_7_i_mux_bus_1_1_rev_T_2 = {MuxWrapper_7_Omuxes_1_1[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_7_i_mux_bus_1_1_rev_T_4 = {{1'd0}, MuxWrapper_7_Omuxes_1_1[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2238 = {_FDPE_7_i_mux_bus_1_1_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_7_i_mux_bus_1_1_rev_T_6 = {{1'd0}, _GEN_2238}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_7_i_mux_bus_1_1_rev_T_7 = _FDPE_7_i_mux_bus_1_1_rev_T_2 | _FDPE_7_i_mux_bus_1_1_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_7_i_mux_bus_1_1_rev_T_8 = {{2'd0}, MuxWrapper_7_Omuxes_1_1[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_7_i_mux_bus_1_1_rev_T_10 = {_FDPE_7_i_mux_bus_1_1_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2240 = {{2'd0}, _FDPE_7_i_mux_bus_1_1_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_7_i_mux_bus_1_1_rev_T_11 = _FDPE_7_i_mux_bus_1_1_rev_T_7 | _GEN_2240; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_7_i_mux_bus_1_1_rev_T_12 = {{3'd0}, MuxWrapper_7_Omuxes_1_1[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_7_i_mux_bus_1_1_rev_T_14 = {{1'd0}, _FDPE_7_i_mux_bus_1_1_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2242 = {{2'd0}, _FDPE_7_i_mux_bus_1_1_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_7_Omuxes_1_2 = MuxesWrapper_7_io_Omuxes_1_2; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_7_i_mux_bus_1_2_rev_T_2 = {MuxWrapper_7_Omuxes_1_2[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_7_i_mux_bus_1_2_rev_T_4 = {{1'd0}, MuxWrapper_7_Omuxes_1_2[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2244 = {_FDPE_7_i_mux_bus_1_2_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_7_i_mux_bus_1_2_rev_T_6 = {{1'd0}, _GEN_2244}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_7_i_mux_bus_1_2_rev_T_7 = _FDPE_7_i_mux_bus_1_2_rev_T_2 | _FDPE_7_i_mux_bus_1_2_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_7_i_mux_bus_1_2_rev_T_8 = {{2'd0}, MuxWrapper_7_Omuxes_1_2[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_7_i_mux_bus_1_2_rev_T_10 = {_FDPE_7_i_mux_bus_1_2_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2246 = {{2'd0}, _FDPE_7_i_mux_bus_1_2_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_7_i_mux_bus_1_2_rev_T_11 = _FDPE_7_i_mux_bus_1_2_rev_T_7 | _GEN_2246; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_7_i_mux_bus_1_2_rev_T_12 = {{3'd0}, MuxWrapper_7_Omuxes_1_2[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_7_i_mux_bus_1_2_rev_T_14 = {{1'd0}, _FDPE_7_i_mux_bus_1_2_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2248 = {{2'd0}, _FDPE_7_i_mux_bus_1_2_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_7_Omuxes_2_0 = MuxesWrapper_7_io_Omuxes_2_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_7_i_mux_bus_2_0_rev_T_2 = {MuxWrapper_7_Omuxes_2_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_7_i_mux_bus_2_0_rev_T_4 = {{1'd0}, MuxWrapper_7_Omuxes_2_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2250 = {_FDPE_7_i_mux_bus_2_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_7_i_mux_bus_2_0_rev_T_6 = {{1'd0}, _GEN_2250}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_7_i_mux_bus_2_0_rev_T_7 = _FDPE_7_i_mux_bus_2_0_rev_T_2 | _FDPE_7_i_mux_bus_2_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_7_i_mux_bus_2_0_rev_T_8 = {{2'd0}, MuxWrapper_7_Omuxes_2_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_7_i_mux_bus_2_0_rev_T_10 = {_FDPE_7_i_mux_bus_2_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2252 = {{2'd0}, _FDPE_7_i_mux_bus_2_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_7_i_mux_bus_2_0_rev_T_11 = _FDPE_7_i_mux_bus_2_0_rev_T_7 | _GEN_2252; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_7_i_mux_bus_2_0_rev_T_12 = {{3'd0}, MuxWrapper_7_Omuxes_2_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_7_i_mux_bus_2_0_rev_T_14 = {{1'd0}, _FDPE_7_i_mux_bus_2_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2254 = {{2'd0}, _FDPE_7_i_mux_bus_2_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_7_Omuxes_2_1 = MuxesWrapper_7_io_Omuxes_2_1; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_7_i_mux_bus_2_1_rev_T_2 = {MuxWrapper_7_Omuxes_2_1[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_7_i_mux_bus_2_1_rev_T_4 = {{1'd0}, MuxWrapper_7_Omuxes_2_1[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2256 = {_FDPE_7_i_mux_bus_2_1_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_7_i_mux_bus_2_1_rev_T_6 = {{1'd0}, _GEN_2256}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_7_i_mux_bus_2_1_rev_T_7 = _FDPE_7_i_mux_bus_2_1_rev_T_2 | _FDPE_7_i_mux_bus_2_1_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_7_i_mux_bus_2_1_rev_T_8 = {{2'd0}, MuxWrapper_7_Omuxes_2_1[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_7_i_mux_bus_2_1_rev_T_10 = {_FDPE_7_i_mux_bus_2_1_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2258 = {{2'd0}, _FDPE_7_i_mux_bus_2_1_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_7_i_mux_bus_2_1_rev_T_11 = _FDPE_7_i_mux_bus_2_1_rev_T_7 | _GEN_2258; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_7_i_mux_bus_2_1_rev_T_12 = {{3'd0}, MuxWrapper_7_Omuxes_2_1[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_7_i_mux_bus_2_1_rev_T_14 = {{1'd0}, _FDPE_7_i_mux_bus_2_1_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2260 = {{2'd0}, _FDPE_7_i_mux_bus_2_1_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_7_Omuxes_3_0 = MuxesWrapper_7_io_Omuxes_3_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_7_i_mux_bus_3_0_rev_T_2 = {MuxWrapper_7_Omuxes_3_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_7_i_mux_bus_3_0_rev_T_4 = {{1'd0}, MuxWrapper_7_Omuxes_3_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2262 = {_FDPE_7_i_mux_bus_3_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_7_i_mux_bus_3_0_rev_T_6 = {{1'd0}, _GEN_2262}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_7_i_mux_bus_3_0_rev_T_7 = _FDPE_7_i_mux_bus_3_0_rev_T_2 | _FDPE_7_i_mux_bus_3_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_7_i_mux_bus_3_0_rev_T_8 = {{2'd0}, MuxWrapper_7_Omuxes_3_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_7_i_mux_bus_3_0_rev_T_10 = {_FDPE_7_i_mux_bus_3_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2264 = {{2'd0}, _FDPE_7_i_mux_bus_3_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_7_i_mux_bus_3_0_rev_T_11 = _FDPE_7_i_mux_bus_3_0_rev_T_7 | _GEN_2264; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_7_i_mux_bus_3_0_rev_T_12 = {{3'd0}, MuxWrapper_7_Omuxes_3_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_7_i_mux_bus_3_0_rev_T_14 = {{1'd0}, _FDPE_7_i_mux_bus_3_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2266 = {{2'd0}, _FDPE_7_i_mux_bus_3_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_8_Omuxes_0_0 = MuxesWrapper_8_io_Omuxes_0_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_8_i_mux_bus_0_0_rev_T_2 = {MuxWrapper_8_Omuxes_0_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_8_i_mux_bus_0_0_rev_T_4 = {{1'd0}, MuxWrapper_8_Omuxes_0_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2268 = {_FDPE_8_i_mux_bus_0_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_8_i_mux_bus_0_0_rev_T_6 = {{1'd0}, _GEN_2268}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_8_i_mux_bus_0_0_rev_T_7 = _FDPE_8_i_mux_bus_0_0_rev_T_2 | _FDPE_8_i_mux_bus_0_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_8_i_mux_bus_0_0_rev_T_8 = {{2'd0}, MuxWrapper_8_Omuxes_0_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_8_i_mux_bus_0_0_rev_T_10 = {_FDPE_8_i_mux_bus_0_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2270 = {{2'd0}, _FDPE_8_i_mux_bus_0_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_8_i_mux_bus_0_0_rev_T_11 = _FDPE_8_i_mux_bus_0_0_rev_T_7 | _GEN_2270; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_8_i_mux_bus_0_0_rev_T_12 = {{3'd0}, MuxWrapper_8_Omuxes_0_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_8_i_mux_bus_0_0_rev_T_14 = {{1'd0}, _FDPE_8_i_mux_bus_0_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2272 = {{2'd0}, _FDPE_8_i_mux_bus_0_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_8_Omuxes_0_1 = MuxesWrapper_8_io_Omuxes_0_1; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_8_i_mux_bus_0_1_rev_T_2 = {MuxWrapper_8_Omuxes_0_1[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_8_i_mux_bus_0_1_rev_T_4 = {{1'd0}, MuxWrapper_8_Omuxes_0_1[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2274 = {_FDPE_8_i_mux_bus_0_1_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_8_i_mux_bus_0_1_rev_T_6 = {{1'd0}, _GEN_2274}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_8_i_mux_bus_0_1_rev_T_7 = _FDPE_8_i_mux_bus_0_1_rev_T_2 | _FDPE_8_i_mux_bus_0_1_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_8_i_mux_bus_0_1_rev_T_8 = {{2'd0}, MuxWrapper_8_Omuxes_0_1[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_8_i_mux_bus_0_1_rev_T_10 = {_FDPE_8_i_mux_bus_0_1_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2276 = {{2'd0}, _FDPE_8_i_mux_bus_0_1_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_8_i_mux_bus_0_1_rev_T_11 = _FDPE_8_i_mux_bus_0_1_rev_T_7 | _GEN_2276; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_8_i_mux_bus_0_1_rev_T_12 = {{3'd0}, MuxWrapper_8_Omuxes_0_1[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_8_i_mux_bus_0_1_rev_T_14 = {{1'd0}, _FDPE_8_i_mux_bus_0_1_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2278 = {{2'd0}, _FDPE_8_i_mux_bus_0_1_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_8_Omuxes_0_2 = MuxesWrapper_8_io_Omuxes_0_2; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_8_i_mux_bus_0_2_rev_T_2 = {MuxWrapper_8_Omuxes_0_2[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_8_i_mux_bus_0_2_rev_T_4 = {{1'd0}, MuxWrapper_8_Omuxes_0_2[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2280 = {_FDPE_8_i_mux_bus_0_2_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_8_i_mux_bus_0_2_rev_T_6 = {{1'd0}, _GEN_2280}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_8_i_mux_bus_0_2_rev_T_7 = _FDPE_8_i_mux_bus_0_2_rev_T_2 | _FDPE_8_i_mux_bus_0_2_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_8_i_mux_bus_0_2_rev_T_8 = {{2'd0}, MuxWrapper_8_Omuxes_0_2[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_8_i_mux_bus_0_2_rev_T_10 = {_FDPE_8_i_mux_bus_0_2_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2282 = {{2'd0}, _FDPE_8_i_mux_bus_0_2_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_8_i_mux_bus_0_2_rev_T_11 = _FDPE_8_i_mux_bus_0_2_rev_T_7 | _GEN_2282; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_8_i_mux_bus_0_2_rev_T_12 = {{3'd0}, MuxWrapper_8_Omuxes_0_2[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_8_i_mux_bus_0_2_rev_T_14 = {{1'd0}, _FDPE_8_i_mux_bus_0_2_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2284 = {{2'd0}, _FDPE_8_i_mux_bus_0_2_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_8_Omuxes_0_3 = MuxesWrapper_8_io_Omuxes_0_3; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_8_i_mux_bus_0_3_rev_T_2 = {MuxWrapper_8_Omuxes_0_3[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_8_i_mux_bus_0_3_rev_T_4 = {{1'd0}, MuxWrapper_8_Omuxes_0_3[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2286 = {_FDPE_8_i_mux_bus_0_3_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_8_i_mux_bus_0_3_rev_T_6 = {{1'd0}, _GEN_2286}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_8_i_mux_bus_0_3_rev_T_7 = _FDPE_8_i_mux_bus_0_3_rev_T_2 | _FDPE_8_i_mux_bus_0_3_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_8_i_mux_bus_0_3_rev_T_8 = {{2'd0}, MuxWrapper_8_Omuxes_0_3[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_8_i_mux_bus_0_3_rev_T_10 = {_FDPE_8_i_mux_bus_0_3_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2288 = {{2'd0}, _FDPE_8_i_mux_bus_0_3_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_8_i_mux_bus_0_3_rev_T_11 = _FDPE_8_i_mux_bus_0_3_rev_T_7 | _GEN_2288; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_8_i_mux_bus_0_3_rev_T_12 = {{3'd0}, MuxWrapper_8_Omuxes_0_3[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_8_i_mux_bus_0_3_rev_T_14 = {{1'd0}, _FDPE_8_i_mux_bus_0_3_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2290 = {{2'd0}, _FDPE_8_i_mux_bus_0_3_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_8_Omuxes_1_0 = MuxesWrapper_8_io_Omuxes_1_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_8_i_mux_bus_1_0_rev_T_2 = {MuxWrapper_8_Omuxes_1_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_8_i_mux_bus_1_0_rev_T_4 = {{1'd0}, MuxWrapper_8_Omuxes_1_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2292 = {_FDPE_8_i_mux_bus_1_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_8_i_mux_bus_1_0_rev_T_6 = {{1'd0}, _GEN_2292}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_8_i_mux_bus_1_0_rev_T_7 = _FDPE_8_i_mux_bus_1_0_rev_T_2 | _FDPE_8_i_mux_bus_1_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_8_i_mux_bus_1_0_rev_T_8 = {{2'd0}, MuxWrapper_8_Omuxes_1_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_8_i_mux_bus_1_0_rev_T_10 = {_FDPE_8_i_mux_bus_1_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2294 = {{2'd0}, _FDPE_8_i_mux_bus_1_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_8_i_mux_bus_1_0_rev_T_11 = _FDPE_8_i_mux_bus_1_0_rev_T_7 | _GEN_2294; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_8_i_mux_bus_1_0_rev_T_12 = {{3'd0}, MuxWrapper_8_Omuxes_1_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_8_i_mux_bus_1_0_rev_T_14 = {{1'd0}, _FDPE_8_i_mux_bus_1_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2296 = {{2'd0}, _FDPE_8_i_mux_bus_1_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_8_Omuxes_1_1 = MuxesWrapper_8_io_Omuxes_1_1; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_8_i_mux_bus_1_1_rev_T_2 = {MuxWrapper_8_Omuxes_1_1[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_8_i_mux_bus_1_1_rev_T_4 = {{1'd0}, MuxWrapper_8_Omuxes_1_1[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2298 = {_FDPE_8_i_mux_bus_1_1_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_8_i_mux_bus_1_1_rev_T_6 = {{1'd0}, _GEN_2298}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_8_i_mux_bus_1_1_rev_T_7 = _FDPE_8_i_mux_bus_1_1_rev_T_2 | _FDPE_8_i_mux_bus_1_1_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_8_i_mux_bus_1_1_rev_T_8 = {{2'd0}, MuxWrapper_8_Omuxes_1_1[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_8_i_mux_bus_1_1_rev_T_10 = {_FDPE_8_i_mux_bus_1_1_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2300 = {{2'd0}, _FDPE_8_i_mux_bus_1_1_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_8_i_mux_bus_1_1_rev_T_11 = _FDPE_8_i_mux_bus_1_1_rev_T_7 | _GEN_2300; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_8_i_mux_bus_1_1_rev_T_12 = {{3'd0}, MuxWrapper_8_Omuxes_1_1[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_8_i_mux_bus_1_1_rev_T_14 = {{1'd0}, _FDPE_8_i_mux_bus_1_1_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2302 = {{2'd0}, _FDPE_8_i_mux_bus_1_1_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_8_Omuxes_1_2 = MuxesWrapper_8_io_Omuxes_1_2; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_8_i_mux_bus_1_2_rev_T_2 = {MuxWrapper_8_Omuxes_1_2[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_8_i_mux_bus_1_2_rev_T_4 = {{1'd0}, MuxWrapper_8_Omuxes_1_2[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2304 = {_FDPE_8_i_mux_bus_1_2_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_8_i_mux_bus_1_2_rev_T_6 = {{1'd0}, _GEN_2304}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_8_i_mux_bus_1_2_rev_T_7 = _FDPE_8_i_mux_bus_1_2_rev_T_2 | _FDPE_8_i_mux_bus_1_2_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_8_i_mux_bus_1_2_rev_T_8 = {{2'd0}, MuxWrapper_8_Omuxes_1_2[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_8_i_mux_bus_1_2_rev_T_10 = {_FDPE_8_i_mux_bus_1_2_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2306 = {{2'd0}, _FDPE_8_i_mux_bus_1_2_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_8_i_mux_bus_1_2_rev_T_11 = _FDPE_8_i_mux_bus_1_2_rev_T_7 | _GEN_2306; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_8_i_mux_bus_1_2_rev_T_12 = {{3'd0}, MuxWrapper_8_Omuxes_1_2[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_8_i_mux_bus_1_2_rev_T_14 = {{1'd0}, _FDPE_8_i_mux_bus_1_2_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2308 = {{2'd0}, _FDPE_8_i_mux_bus_1_2_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_8_Omuxes_2_0 = MuxesWrapper_8_io_Omuxes_2_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_8_i_mux_bus_2_0_rev_T_2 = {MuxWrapper_8_Omuxes_2_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_8_i_mux_bus_2_0_rev_T_4 = {{1'd0}, MuxWrapper_8_Omuxes_2_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2310 = {_FDPE_8_i_mux_bus_2_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_8_i_mux_bus_2_0_rev_T_6 = {{1'd0}, _GEN_2310}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_8_i_mux_bus_2_0_rev_T_7 = _FDPE_8_i_mux_bus_2_0_rev_T_2 | _FDPE_8_i_mux_bus_2_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_8_i_mux_bus_2_0_rev_T_8 = {{2'd0}, MuxWrapper_8_Omuxes_2_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_8_i_mux_bus_2_0_rev_T_10 = {_FDPE_8_i_mux_bus_2_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2312 = {{2'd0}, _FDPE_8_i_mux_bus_2_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_8_i_mux_bus_2_0_rev_T_11 = _FDPE_8_i_mux_bus_2_0_rev_T_7 | _GEN_2312; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_8_i_mux_bus_2_0_rev_T_12 = {{3'd0}, MuxWrapper_8_Omuxes_2_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_8_i_mux_bus_2_0_rev_T_14 = {{1'd0}, _FDPE_8_i_mux_bus_2_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2314 = {{2'd0}, _FDPE_8_i_mux_bus_2_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_8_Omuxes_2_1 = MuxesWrapper_8_io_Omuxes_2_1; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_8_i_mux_bus_2_1_rev_T_2 = {MuxWrapper_8_Omuxes_2_1[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_8_i_mux_bus_2_1_rev_T_4 = {{1'd0}, MuxWrapper_8_Omuxes_2_1[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2316 = {_FDPE_8_i_mux_bus_2_1_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_8_i_mux_bus_2_1_rev_T_6 = {{1'd0}, _GEN_2316}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_8_i_mux_bus_2_1_rev_T_7 = _FDPE_8_i_mux_bus_2_1_rev_T_2 | _FDPE_8_i_mux_bus_2_1_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_8_i_mux_bus_2_1_rev_T_8 = {{2'd0}, MuxWrapper_8_Omuxes_2_1[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_8_i_mux_bus_2_1_rev_T_10 = {_FDPE_8_i_mux_bus_2_1_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2318 = {{2'd0}, _FDPE_8_i_mux_bus_2_1_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_8_i_mux_bus_2_1_rev_T_11 = _FDPE_8_i_mux_bus_2_1_rev_T_7 | _GEN_2318; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_8_i_mux_bus_2_1_rev_T_12 = {{3'd0}, MuxWrapper_8_Omuxes_2_1[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_8_i_mux_bus_2_1_rev_T_14 = {{1'd0}, _FDPE_8_i_mux_bus_2_1_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2320 = {{2'd0}, _FDPE_8_i_mux_bus_2_1_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_8_Omuxes_3_0 = MuxesWrapper_8_io_Omuxes_3_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_8_i_mux_bus_3_0_rev_T_2 = {MuxWrapper_8_Omuxes_3_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_8_i_mux_bus_3_0_rev_T_4 = {{1'd0}, MuxWrapper_8_Omuxes_3_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2322 = {_FDPE_8_i_mux_bus_3_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_8_i_mux_bus_3_0_rev_T_6 = {{1'd0}, _GEN_2322}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_8_i_mux_bus_3_0_rev_T_7 = _FDPE_8_i_mux_bus_3_0_rev_T_2 | _FDPE_8_i_mux_bus_3_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_8_i_mux_bus_3_0_rev_T_8 = {{2'd0}, MuxWrapper_8_Omuxes_3_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_8_i_mux_bus_3_0_rev_T_10 = {_FDPE_8_i_mux_bus_3_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2324 = {{2'd0}, _FDPE_8_i_mux_bus_3_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_8_i_mux_bus_3_0_rev_T_11 = _FDPE_8_i_mux_bus_3_0_rev_T_7 | _GEN_2324; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_8_i_mux_bus_3_0_rev_T_12 = {{3'd0}, MuxWrapper_8_Omuxes_3_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_8_i_mux_bus_3_0_rev_T_14 = {{1'd0}, _FDPE_8_i_mux_bus_3_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2326 = {{2'd0}, _FDPE_8_i_mux_bus_3_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_9_Omuxes_0_0 = MuxesWrapper_9_io_Omuxes_0_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_9_i_mux_bus_0_0_rev_T_2 = {MuxWrapper_9_Omuxes_0_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_9_i_mux_bus_0_0_rev_T_4 = {{1'd0}, MuxWrapper_9_Omuxes_0_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2328 = {_FDPE_9_i_mux_bus_0_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_9_i_mux_bus_0_0_rev_T_6 = {{1'd0}, _GEN_2328}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_9_i_mux_bus_0_0_rev_T_7 = _FDPE_9_i_mux_bus_0_0_rev_T_2 | _FDPE_9_i_mux_bus_0_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_9_i_mux_bus_0_0_rev_T_8 = {{2'd0}, MuxWrapper_9_Omuxes_0_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_9_i_mux_bus_0_0_rev_T_10 = {_FDPE_9_i_mux_bus_0_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2330 = {{2'd0}, _FDPE_9_i_mux_bus_0_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_9_i_mux_bus_0_0_rev_T_11 = _FDPE_9_i_mux_bus_0_0_rev_T_7 | _GEN_2330; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_9_i_mux_bus_0_0_rev_T_12 = {{3'd0}, MuxWrapper_9_Omuxes_0_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_9_i_mux_bus_0_0_rev_T_14 = {{1'd0}, _FDPE_9_i_mux_bus_0_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2332 = {{2'd0}, _FDPE_9_i_mux_bus_0_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_9_Omuxes_0_1 = MuxesWrapper_9_io_Omuxes_0_1; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_9_i_mux_bus_0_1_rev_T_2 = {MuxWrapper_9_Omuxes_0_1[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_9_i_mux_bus_0_1_rev_T_4 = {{1'd0}, MuxWrapper_9_Omuxes_0_1[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2334 = {_FDPE_9_i_mux_bus_0_1_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_9_i_mux_bus_0_1_rev_T_6 = {{1'd0}, _GEN_2334}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_9_i_mux_bus_0_1_rev_T_7 = _FDPE_9_i_mux_bus_0_1_rev_T_2 | _FDPE_9_i_mux_bus_0_1_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_9_i_mux_bus_0_1_rev_T_8 = {{2'd0}, MuxWrapper_9_Omuxes_0_1[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_9_i_mux_bus_0_1_rev_T_10 = {_FDPE_9_i_mux_bus_0_1_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2336 = {{2'd0}, _FDPE_9_i_mux_bus_0_1_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_9_i_mux_bus_0_1_rev_T_11 = _FDPE_9_i_mux_bus_0_1_rev_T_7 | _GEN_2336; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_9_i_mux_bus_0_1_rev_T_12 = {{3'd0}, MuxWrapper_9_Omuxes_0_1[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_9_i_mux_bus_0_1_rev_T_14 = {{1'd0}, _FDPE_9_i_mux_bus_0_1_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2338 = {{2'd0}, _FDPE_9_i_mux_bus_0_1_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_9_Omuxes_0_2 = MuxesWrapper_9_io_Omuxes_0_2; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_9_i_mux_bus_0_2_rev_T_2 = {MuxWrapper_9_Omuxes_0_2[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_9_i_mux_bus_0_2_rev_T_4 = {{1'd0}, MuxWrapper_9_Omuxes_0_2[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2340 = {_FDPE_9_i_mux_bus_0_2_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_9_i_mux_bus_0_2_rev_T_6 = {{1'd0}, _GEN_2340}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_9_i_mux_bus_0_2_rev_T_7 = _FDPE_9_i_mux_bus_0_2_rev_T_2 | _FDPE_9_i_mux_bus_0_2_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_9_i_mux_bus_0_2_rev_T_8 = {{2'd0}, MuxWrapper_9_Omuxes_0_2[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_9_i_mux_bus_0_2_rev_T_10 = {_FDPE_9_i_mux_bus_0_2_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2342 = {{2'd0}, _FDPE_9_i_mux_bus_0_2_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_9_i_mux_bus_0_2_rev_T_11 = _FDPE_9_i_mux_bus_0_2_rev_T_7 | _GEN_2342; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_9_i_mux_bus_0_2_rev_T_12 = {{3'd0}, MuxWrapper_9_Omuxes_0_2[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_9_i_mux_bus_0_2_rev_T_14 = {{1'd0}, _FDPE_9_i_mux_bus_0_2_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2344 = {{2'd0}, _FDPE_9_i_mux_bus_0_2_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_9_Omuxes_0_3 = MuxesWrapper_9_io_Omuxes_0_3; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_9_i_mux_bus_0_3_rev_T_2 = {MuxWrapper_9_Omuxes_0_3[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_9_i_mux_bus_0_3_rev_T_4 = {{1'd0}, MuxWrapper_9_Omuxes_0_3[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2346 = {_FDPE_9_i_mux_bus_0_3_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_9_i_mux_bus_0_3_rev_T_6 = {{1'd0}, _GEN_2346}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_9_i_mux_bus_0_3_rev_T_7 = _FDPE_9_i_mux_bus_0_3_rev_T_2 | _FDPE_9_i_mux_bus_0_3_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_9_i_mux_bus_0_3_rev_T_8 = {{2'd0}, MuxWrapper_9_Omuxes_0_3[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_9_i_mux_bus_0_3_rev_T_10 = {_FDPE_9_i_mux_bus_0_3_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2348 = {{2'd0}, _FDPE_9_i_mux_bus_0_3_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_9_i_mux_bus_0_3_rev_T_11 = _FDPE_9_i_mux_bus_0_3_rev_T_7 | _GEN_2348; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_9_i_mux_bus_0_3_rev_T_12 = {{3'd0}, MuxWrapper_9_Omuxes_0_3[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_9_i_mux_bus_0_3_rev_T_14 = {{1'd0}, _FDPE_9_i_mux_bus_0_3_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2350 = {{2'd0}, _FDPE_9_i_mux_bus_0_3_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_9_Omuxes_1_0 = MuxesWrapper_9_io_Omuxes_1_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_9_i_mux_bus_1_0_rev_T_2 = {MuxWrapper_9_Omuxes_1_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_9_i_mux_bus_1_0_rev_T_4 = {{1'd0}, MuxWrapper_9_Omuxes_1_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2352 = {_FDPE_9_i_mux_bus_1_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_9_i_mux_bus_1_0_rev_T_6 = {{1'd0}, _GEN_2352}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_9_i_mux_bus_1_0_rev_T_7 = _FDPE_9_i_mux_bus_1_0_rev_T_2 | _FDPE_9_i_mux_bus_1_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_9_i_mux_bus_1_0_rev_T_8 = {{2'd0}, MuxWrapper_9_Omuxes_1_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_9_i_mux_bus_1_0_rev_T_10 = {_FDPE_9_i_mux_bus_1_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2354 = {{2'd0}, _FDPE_9_i_mux_bus_1_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_9_i_mux_bus_1_0_rev_T_11 = _FDPE_9_i_mux_bus_1_0_rev_T_7 | _GEN_2354; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_9_i_mux_bus_1_0_rev_T_12 = {{3'd0}, MuxWrapper_9_Omuxes_1_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_9_i_mux_bus_1_0_rev_T_14 = {{1'd0}, _FDPE_9_i_mux_bus_1_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2356 = {{2'd0}, _FDPE_9_i_mux_bus_1_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_9_Omuxes_1_1 = MuxesWrapper_9_io_Omuxes_1_1; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_9_i_mux_bus_1_1_rev_T_2 = {MuxWrapper_9_Omuxes_1_1[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_9_i_mux_bus_1_1_rev_T_4 = {{1'd0}, MuxWrapper_9_Omuxes_1_1[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2358 = {_FDPE_9_i_mux_bus_1_1_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_9_i_mux_bus_1_1_rev_T_6 = {{1'd0}, _GEN_2358}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_9_i_mux_bus_1_1_rev_T_7 = _FDPE_9_i_mux_bus_1_1_rev_T_2 | _FDPE_9_i_mux_bus_1_1_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_9_i_mux_bus_1_1_rev_T_8 = {{2'd0}, MuxWrapper_9_Omuxes_1_1[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_9_i_mux_bus_1_1_rev_T_10 = {_FDPE_9_i_mux_bus_1_1_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2360 = {{2'd0}, _FDPE_9_i_mux_bus_1_1_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_9_i_mux_bus_1_1_rev_T_11 = _FDPE_9_i_mux_bus_1_1_rev_T_7 | _GEN_2360; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_9_i_mux_bus_1_1_rev_T_12 = {{3'd0}, MuxWrapper_9_Omuxes_1_1[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_9_i_mux_bus_1_1_rev_T_14 = {{1'd0}, _FDPE_9_i_mux_bus_1_1_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2362 = {{2'd0}, _FDPE_9_i_mux_bus_1_1_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_9_Omuxes_1_2 = MuxesWrapper_9_io_Omuxes_1_2; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_9_i_mux_bus_1_2_rev_T_2 = {MuxWrapper_9_Omuxes_1_2[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_9_i_mux_bus_1_2_rev_T_4 = {{1'd0}, MuxWrapper_9_Omuxes_1_2[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2364 = {_FDPE_9_i_mux_bus_1_2_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_9_i_mux_bus_1_2_rev_T_6 = {{1'd0}, _GEN_2364}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_9_i_mux_bus_1_2_rev_T_7 = _FDPE_9_i_mux_bus_1_2_rev_T_2 | _FDPE_9_i_mux_bus_1_2_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_9_i_mux_bus_1_2_rev_T_8 = {{2'd0}, MuxWrapper_9_Omuxes_1_2[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_9_i_mux_bus_1_2_rev_T_10 = {_FDPE_9_i_mux_bus_1_2_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2366 = {{2'd0}, _FDPE_9_i_mux_bus_1_2_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_9_i_mux_bus_1_2_rev_T_11 = _FDPE_9_i_mux_bus_1_2_rev_T_7 | _GEN_2366; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_9_i_mux_bus_1_2_rev_T_12 = {{3'd0}, MuxWrapper_9_Omuxes_1_2[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_9_i_mux_bus_1_2_rev_T_14 = {{1'd0}, _FDPE_9_i_mux_bus_1_2_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2368 = {{2'd0}, _FDPE_9_i_mux_bus_1_2_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_9_Omuxes_2_0 = MuxesWrapper_9_io_Omuxes_2_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_9_i_mux_bus_2_0_rev_T_2 = {MuxWrapper_9_Omuxes_2_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_9_i_mux_bus_2_0_rev_T_4 = {{1'd0}, MuxWrapper_9_Omuxes_2_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2370 = {_FDPE_9_i_mux_bus_2_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_9_i_mux_bus_2_0_rev_T_6 = {{1'd0}, _GEN_2370}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_9_i_mux_bus_2_0_rev_T_7 = _FDPE_9_i_mux_bus_2_0_rev_T_2 | _FDPE_9_i_mux_bus_2_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_9_i_mux_bus_2_0_rev_T_8 = {{2'd0}, MuxWrapper_9_Omuxes_2_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_9_i_mux_bus_2_0_rev_T_10 = {_FDPE_9_i_mux_bus_2_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2372 = {{2'd0}, _FDPE_9_i_mux_bus_2_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_9_i_mux_bus_2_0_rev_T_11 = _FDPE_9_i_mux_bus_2_0_rev_T_7 | _GEN_2372; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_9_i_mux_bus_2_0_rev_T_12 = {{3'd0}, MuxWrapper_9_Omuxes_2_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_9_i_mux_bus_2_0_rev_T_14 = {{1'd0}, _FDPE_9_i_mux_bus_2_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2374 = {{2'd0}, _FDPE_9_i_mux_bus_2_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_9_Omuxes_2_1 = MuxesWrapper_9_io_Omuxes_2_1; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_9_i_mux_bus_2_1_rev_T_2 = {MuxWrapper_9_Omuxes_2_1[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_9_i_mux_bus_2_1_rev_T_4 = {{1'd0}, MuxWrapper_9_Omuxes_2_1[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2376 = {_FDPE_9_i_mux_bus_2_1_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_9_i_mux_bus_2_1_rev_T_6 = {{1'd0}, _GEN_2376}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_9_i_mux_bus_2_1_rev_T_7 = _FDPE_9_i_mux_bus_2_1_rev_T_2 | _FDPE_9_i_mux_bus_2_1_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_9_i_mux_bus_2_1_rev_T_8 = {{2'd0}, MuxWrapper_9_Omuxes_2_1[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_9_i_mux_bus_2_1_rev_T_10 = {_FDPE_9_i_mux_bus_2_1_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2378 = {{2'd0}, _FDPE_9_i_mux_bus_2_1_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_9_i_mux_bus_2_1_rev_T_11 = _FDPE_9_i_mux_bus_2_1_rev_T_7 | _GEN_2378; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_9_i_mux_bus_2_1_rev_T_12 = {{3'd0}, MuxWrapper_9_Omuxes_2_1[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_9_i_mux_bus_2_1_rev_T_14 = {{1'd0}, _FDPE_9_i_mux_bus_2_1_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2380 = {{2'd0}, _FDPE_9_i_mux_bus_2_1_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_9_Omuxes_3_0 = MuxesWrapper_9_io_Omuxes_3_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_9_i_mux_bus_3_0_rev_T_2 = {MuxWrapper_9_Omuxes_3_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_9_i_mux_bus_3_0_rev_T_4 = {{1'd0}, MuxWrapper_9_Omuxes_3_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2382 = {_FDPE_9_i_mux_bus_3_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_9_i_mux_bus_3_0_rev_T_6 = {{1'd0}, _GEN_2382}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_9_i_mux_bus_3_0_rev_T_7 = _FDPE_9_i_mux_bus_3_0_rev_T_2 | _FDPE_9_i_mux_bus_3_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_9_i_mux_bus_3_0_rev_T_8 = {{2'd0}, MuxWrapper_9_Omuxes_3_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_9_i_mux_bus_3_0_rev_T_10 = {_FDPE_9_i_mux_bus_3_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2384 = {{2'd0}, _FDPE_9_i_mux_bus_3_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_9_i_mux_bus_3_0_rev_T_11 = _FDPE_9_i_mux_bus_3_0_rev_T_7 | _GEN_2384; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_9_i_mux_bus_3_0_rev_T_12 = {{3'd0}, MuxWrapper_9_Omuxes_3_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_9_i_mux_bus_3_0_rev_T_14 = {{1'd0}, _FDPE_9_i_mux_bus_3_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2386 = {{2'd0}, _FDPE_9_i_mux_bus_3_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_10_Omuxes_0_0 = MuxesWrapper_10_io_Omuxes_0_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_10_i_mux_bus_0_0_rev_T_2 = {MuxWrapper_10_Omuxes_0_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_10_i_mux_bus_0_0_rev_T_4 = {{1'd0}, MuxWrapper_10_Omuxes_0_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2388 = {_FDPE_10_i_mux_bus_0_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_10_i_mux_bus_0_0_rev_T_6 = {{1'd0}, _GEN_2388}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_10_i_mux_bus_0_0_rev_T_7 = _FDPE_10_i_mux_bus_0_0_rev_T_2 | _FDPE_10_i_mux_bus_0_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_10_i_mux_bus_0_0_rev_T_8 = {{2'd0}, MuxWrapper_10_Omuxes_0_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_10_i_mux_bus_0_0_rev_T_10 = {_FDPE_10_i_mux_bus_0_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2390 = {{2'd0}, _FDPE_10_i_mux_bus_0_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_10_i_mux_bus_0_0_rev_T_11 = _FDPE_10_i_mux_bus_0_0_rev_T_7 | _GEN_2390; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_10_i_mux_bus_0_0_rev_T_12 = {{3'd0}, MuxWrapper_10_Omuxes_0_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_10_i_mux_bus_0_0_rev_T_14 = {{1'd0}, _FDPE_10_i_mux_bus_0_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2392 = {{2'd0}, _FDPE_10_i_mux_bus_0_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_10_Omuxes_0_1 = MuxesWrapper_10_io_Omuxes_0_1; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_10_i_mux_bus_0_1_rev_T_2 = {MuxWrapper_10_Omuxes_0_1[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_10_i_mux_bus_0_1_rev_T_4 = {{1'd0}, MuxWrapper_10_Omuxes_0_1[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2394 = {_FDPE_10_i_mux_bus_0_1_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_10_i_mux_bus_0_1_rev_T_6 = {{1'd0}, _GEN_2394}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_10_i_mux_bus_0_1_rev_T_7 = _FDPE_10_i_mux_bus_0_1_rev_T_2 | _FDPE_10_i_mux_bus_0_1_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_10_i_mux_bus_0_1_rev_T_8 = {{2'd0}, MuxWrapper_10_Omuxes_0_1[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_10_i_mux_bus_0_1_rev_T_10 = {_FDPE_10_i_mux_bus_0_1_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2396 = {{2'd0}, _FDPE_10_i_mux_bus_0_1_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_10_i_mux_bus_0_1_rev_T_11 = _FDPE_10_i_mux_bus_0_1_rev_T_7 | _GEN_2396; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_10_i_mux_bus_0_1_rev_T_12 = {{3'd0}, MuxWrapper_10_Omuxes_0_1[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_10_i_mux_bus_0_1_rev_T_14 = {{1'd0}, _FDPE_10_i_mux_bus_0_1_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2398 = {{2'd0}, _FDPE_10_i_mux_bus_0_1_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_10_Omuxes_0_2 = MuxesWrapper_10_io_Omuxes_0_2; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_10_i_mux_bus_0_2_rev_T_2 = {MuxWrapper_10_Omuxes_0_2[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_10_i_mux_bus_0_2_rev_T_4 = {{1'd0}, MuxWrapper_10_Omuxes_0_2[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2400 = {_FDPE_10_i_mux_bus_0_2_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_10_i_mux_bus_0_2_rev_T_6 = {{1'd0}, _GEN_2400}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_10_i_mux_bus_0_2_rev_T_7 = _FDPE_10_i_mux_bus_0_2_rev_T_2 | _FDPE_10_i_mux_bus_0_2_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_10_i_mux_bus_0_2_rev_T_8 = {{2'd0}, MuxWrapper_10_Omuxes_0_2[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_10_i_mux_bus_0_2_rev_T_10 = {_FDPE_10_i_mux_bus_0_2_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2402 = {{2'd0}, _FDPE_10_i_mux_bus_0_2_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_10_i_mux_bus_0_2_rev_T_11 = _FDPE_10_i_mux_bus_0_2_rev_T_7 | _GEN_2402; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_10_i_mux_bus_0_2_rev_T_12 = {{3'd0}, MuxWrapper_10_Omuxes_0_2[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_10_i_mux_bus_0_2_rev_T_14 = {{1'd0}, _FDPE_10_i_mux_bus_0_2_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2404 = {{2'd0}, _FDPE_10_i_mux_bus_0_2_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_10_Omuxes_0_3 = MuxesWrapper_10_io_Omuxes_0_3; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_10_i_mux_bus_0_3_rev_T_2 = {MuxWrapper_10_Omuxes_0_3[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_10_i_mux_bus_0_3_rev_T_4 = {{1'd0}, MuxWrapper_10_Omuxes_0_3[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2406 = {_FDPE_10_i_mux_bus_0_3_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_10_i_mux_bus_0_3_rev_T_6 = {{1'd0}, _GEN_2406}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_10_i_mux_bus_0_3_rev_T_7 = _FDPE_10_i_mux_bus_0_3_rev_T_2 | _FDPE_10_i_mux_bus_0_3_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_10_i_mux_bus_0_3_rev_T_8 = {{2'd0}, MuxWrapper_10_Omuxes_0_3[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_10_i_mux_bus_0_3_rev_T_10 = {_FDPE_10_i_mux_bus_0_3_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2408 = {{2'd0}, _FDPE_10_i_mux_bus_0_3_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_10_i_mux_bus_0_3_rev_T_11 = _FDPE_10_i_mux_bus_0_3_rev_T_7 | _GEN_2408; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_10_i_mux_bus_0_3_rev_T_12 = {{3'd0}, MuxWrapper_10_Omuxes_0_3[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_10_i_mux_bus_0_3_rev_T_14 = {{1'd0}, _FDPE_10_i_mux_bus_0_3_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2410 = {{2'd0}, _FDPE_10_i_mux_bus_0_3_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_10_Omuxes_1_0 = MuxesWrapper_10_io_Omuxes_1_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_10_i_mux_bus_1_0_rev_T_2 = {MuxWrapper_10_Omuxes_1_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_10_i_mux_bus_1_0_rev_T_4 = {{1'd0}, MuxWrapper_10_Omuxes_1_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2412 = {_FDPE_10_i_mux_bus_1_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_10_i_mux_bus_1_0_rev_T_6 = {{1'd0}, _GEN_2412}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_10_i_mux_bus_1_0_rev_T_7 = _FDPE_10_i_mux_bus_1_0_rev_T_2 | _FDPE_10_i_mux_bus_1_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_10_i_mux_bus_1_0_rev_T_8 = {{2'd0}, MuxWrapper_10_Omuxes_1_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_10_i_mux_bus_1_0_rev_T_10 = {_FDPE_10_i_mux_bus_1_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2414 = {{2'd0}, _FDPE_10_i_mux_bus_1_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_10_i_mux_bus_1_0_rev_T_11 = _FDPE_10_i_mux_bus_1_0_rev_T_7 | _GEN_2414; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_10_i_mux_bus_1_0_rev_T_12 = {{3'd0}, MuxWrapper_10_Omuxes_1_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_10_i_mux_bus_1_0_rev_T_14 = {{1'd0}, _FDPE_10_i_mux_bus_1_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2416 = {{2'd0}, _FDPE_10_i_mux_bus_1_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_10_Omuxes_1_1 = MuxesWrapper_10_io_Omuxes_1_1; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_10_i_mux_bus_1_1_rev_T_2 = {MuxWrapper_10_Omuxes_1_1[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_10_i_mux_bus_1_1_rev_T_4 = {{1'd0}, MuxWrapper_10_Omuxes_1_1[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2418 = {_FDPE_10_i_mux_bus_1_1_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_10_i_mux_bus_1_1_rev_T_6 = {{1'd0}, _GEN_2418}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_10_i_mux_bus_1_1_rev_T_7 = _FDPE_10_i_mux_bus_1_1_rev_T_2 | _FDPE_10_i_mux_bus_1_1_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_10_i_mux_bus_1_1_rev_T_8 = {{2'd0}, MuxWrapper_10_Omuxes_1_1[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_10_i_mux_bus_1_1_rev_T_10 = {_FDPE_10_i_mux_bus_1_1_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2420 = {{2'd0}, _FDPE_10_i_mux_bus_1_1_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_10_i_mux_bus_1_1_rev_T_11 = _FDPE_10_i_mux_bus_1_1_rev_T_7 | _GEN_2420; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_10_i_mux_bus_1_1_rev_T_12 = {{3'd0}, MuxWrapper_10_Omuxes_1_1[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_10_i_mux_bus_1_1_rev_T_14 = {{1'd0}, _FDPE_10_i_mux_bus_1_1_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2422 = {{2'd0}, _FDPE_10_i_mux_bus_1_1_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_10_Omuxes_1_2 = MuxesWrapper_10_io_Omuxes_1_2; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_10_i_mux_bus_1_2_rev_T_2 = {MuxWrapper_10_Omuxes_1_2[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_10_i_mux_bus_1_2_rev_T_4 = {{1'd0}, MuxWrapper_10_Omuxes_1_2[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2424 = {_FDPE_10_i_mux_bus_1_2_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_10_i_mux_bus_1_2_rev_T_6 = {{1'd0}, _GEN_2424}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_10_i_mux_bus_1_2_rev_T_7 = _FDPE_10_i_mux_bus_1_2_rev_T_2 | _FDPE_10_i_mux_bus_1_2_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_10_i_mux_bus_1_2_rev_T_8 = {{2'd0}, MuxWrapper_10_Omuxes_1_2[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_10_i_mux_bus_1_2_rev_T_10 = {_FDPE_10_i_mux_bus_1_2_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2426 = {{2'd0}, _FDPE_10_i_mux_bus_1_2_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_10_i_mux_bus_1_2_rev_T_11 = _FDPE_10_i_mux_bus_1_2_rev_T_7 | _GEN_2426; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_10_i_mux_bus_1_2_rev_T_12 = {{3'd0}, MuxWrapper_10_Omuxes_1_2[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_10_i_mux_bus_1_2_rev_T_14 = {{1'd0}, _FDPE_10_i_mux_bus_1_2_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2428 = {{2'd0}, _FDPE_10_i_mux_bus_1_2_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_10_Omuxes_2_0 = MuxesWrapper_10_io_Omuxes_2_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_10_i_mux_bus_2_0_rev_T_2 = {MuxWrapper_10_Omuxes_2_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_10_i_mux_bus_2_0_rev_T_4 = {{1'd0}, MuxWrapper_10_Omuxes_2_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2430 = {_FDPE_10_i_mux_bus_2_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_10_i_mux_bus_2_0_rev_T_6 = {{1'd0}, _GEN_2430}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_10_i_mux_bus_2_0_rev_T_7 = _FDPE_10_i_mux_bus_2_0_rev_T_2 | _FDPE_10_i_mux_bus_2_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_10_i_mux_bus_2_0_rev_T_8 = {{2'd0}, MuxWrapper_10_Omuxes_2_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_10_i_mux_bus_2_0_rev_T_10 = {_FDPE_10_i_mux_bus_2_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2432 = {{2'd0}, _FDPE_10_i_mux_bus_2_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_10_i_mux_bus_2_0_rev_T_11 = _FDPE_10_i_mux_bus_2_0_rev_T_7 | _GEN_2432; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_10_i_mux_bus_2_0_rev_T_12 = {{3'd0}, MuxWrapper_10_Omuxes_2_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_10_i_mux_bus_2_0_rev_T_14 = {{1'd0}, _FDPE_10_i_mux_bus_2_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2434 = {{2'd0}, _FDPE_10_i_mux_bus_2_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_10_Omuxes_2_1 = MuxesWrapper_10_io_Omuxes_2_1; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_10_i_mux_bus_2_1_rev_T_2 = {MuxWrapper_10_Omuxes_2_1[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_10_i_mux_bus_2_1_rev_T_4 = {{1'd0}, MuxWrapper_10_Omuxes_2_1[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2436 = {_FDPE_10_i_mux_bus_2_1_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_10_i_mux_bus_2_1_rev_T_6 = {{1'd0}, _GEN_2436}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_10_i_mux_bus_2_1_rev_T_7 = _FDPE_10_i_mux_bus_2_1_rev_T_2 | _FDPE_10_i_mux_bus_2_1_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_10_i_mux_bus_2_1_rev_T_8 = {{2'd0}, MuxWrapper_10_Omuxes_2_1[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_10_i_mux_bus_2_1_rev_T_10 = {_FDPE_10_i_mux_bus_2_1_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2438 = {{2'd0}, _FDPE_10_i_mux_bus_2_1_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_10_i_mux_bus_2_1_rev_T_11 = _FDPE_10_i_mux_bus_2_1_rev_T_7 | _GEN_2438; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_10_i_mux_bus_2_1_rev_T_12 = {{3'd0}, MuxWrapper_10_Omuxes_2_1[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_10_i_mux_bus_2_1_rev_T_14 = {{1'd0}, _FDPE_10_i_mux_bus_2_1_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2440 = {{2'd0}, _FDPE_10_i_mux_bus_2_1_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_10_Omuxes_3_0 = MuxesWrapper_10_io_Omuxes_3_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_10_i_mux_bus_3_0_rev_T_2 = {MuxWrapper_10_Omuxes_3_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_10_i_mux_bus_3_0_rev_T_4 = {{1'd0}, MuxWrapper_10_Omuxes_3_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2442 = {_FDPE_10_i_mux_bus_3_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_10_i_mux_bus_3_0_rev_T_6 = {{1'd0}, _GEN_2442}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_10_i_mux_bus_3_0_rev_T_7 = _FDPE_10_i_mux_bus_3_0_rev_T_2 | _FDPE_10_i_mux_bus_3_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_10_i_mux_bus_3_0_rev_T_8 = {{2'd0}, MuxWrapper_10_Omuxes_3_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_10_i_mux_bus_3_0_rev_T_10 = {_FDPE_10_i_mux_bus_3_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2444 = {{2'd0}, _FDPE_10_i_mux_bus_3_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_10_i_mux_bus_3_0_rev_T_11 = _FDPE_10_i_mux_bus_3_0_rev_T_7 | _GEN_2444; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_10_i_mux_bus_3_0_rev_T_12 = {{3'd0}, MuxWrapper_10_Omuxes_3_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_10_i_mux_bus_3_0_rev_T_14 = {{1'd0}, _FDPE_10_i_mux_bus_3_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2446 = {{2'd0}, _FDPE_10_i_mux_bus_3_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_11_Omuxes_0_0 = MuxesWrapper_11_io_Omuxes_0_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_11_i_mux_bus_0_0_rev_T_2 = {MuxWrapper_11_Omuxes_0_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_11_i_mux_bus_0_0_rev_T_4 = {{1'd0}, MuxWrapper_11_Omuxes_0_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2448 = {_FDPE_11_i_mux_bus_0_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_11_i_mux_bus_0_0_rev_T_6 = {{1'd0}, _GEN_2448}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_11_i_mux_bus_0_0_rev_T_7 = _FDPE_11_i_mux_bus_0_0_rev_T_2 | _FDPE_11_i_mux_bus_0_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_11_i_mux_bus_0_0_rev_T_8 = {{2'd0}, MuxWrapper_11_Omuxes_0_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_11_i_mux_bus_0_0_rev_T_10 = {_FDPE_11_i_mux_bus_0_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2450 = {{2'd0}, _FDPE_11_i_mux_bus_0_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_11_i_mux_bus_0_0_rev_T_11 = _FDPE_11_i_mux_bus_0_0_rev_T_7 | _GEN_2450; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_11_i_mux_bus_0_0_rev_T_12 = {{3'd0}, MuxWrapper_11_Omuxes_0_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_11_i_mux_bus_0_0_rev_T_14 = {{1'd0}, _FDPE_11_i_mux_bus_0_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2452 = {{2'd0}, _FDPE_11_i_mux_bus_0_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_11_Omuxes_0_1 = MuxesWrapper_11_io_Omuxes_0_1; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_11_i_mux_bus_0_1_rev_T_2 = {MuxWrapper_11_Omuxes_0_1[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_11_i_mux_bus_0_1_rev_T_4 = {{1'd0}, MuxWrapper_11_Omuxes_0_1[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2454 = {_FDPE_11_i_mux_bus_0_1_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_11_i_mux_bus_0_1_rev_T_6 = {{1'd0}, _GEN_2454}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_11_i_mux_bus_0_1_rev_T_7 = _FDPE_11_i_mux_bus_0_1_rev_T_2 | _FDPE_11_i_mux_bus_0_1_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_11_i_mux_bus_0_1_rev_T_8 = {{2'd0}, MuxWrapper_11_Omuxes_0_1[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_11_i_mux_bus_0_1_rev_T_10 = {_FDPE_11_i_mux_bus_0_1_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2456 = {{2'd0}, _FDPE_11_i_mux_bus_0_1_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_11_i_mux_bus_0_1_rev_T_11 = _FDPE_11_i_mux_bus_0_1_rev_T_7 | _GEN_2456; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_11_i_mux_bus_0_1_rev_T_12 = {{3'd0}, MuxWrapper_11_Omuxes_0_1[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_11_i_mux_bus_0_1_rev_T_14 = {{1'd0}, _FDPE_11_i_mux_bus_0_1_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2458 = {{2'd0}, _FDPE_11_i_mux_bus_0_1_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_11_Omuxes_0_2 = MuxesWrapper_11_io_Omuxes_0_2; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_11_i_mux_bus_0_2_rev_T_2 = {MuxWrapper_11_Omuxes_0_2[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_11_i_mux_bus_0_2_rev_T_4 = {{1'd0}, MuxWrapper_11_Omuxes_0_2[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2460 = {_FDPE_11_i_mux_bus_0_2_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_11_i_mux_bus_0_2_rev_T_6 = {{1'd0}, _GEN_2460}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_11_i_mux_bus_0_2_rev_T_7 = _FDPE_11_i_mux_bus_0_2_rev_T_2 | _FDPE_11_i_mux_bus_0_2_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_11_i_mux_bus_0_2_rev_T_8 = {{2'd0}, MuxWrapper_11_Omuxes_0_2[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_11_i_mux_bus_0_2_rev_T_10 = {_FDPE_11_i_mux_bus_0_2_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2462 = {{2'd0}, _FDPE_11_i_mux_bus_0_2_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_11_i_mux_bus_0_2_rev_T_11 = _FDPE_11_i_mux_bus_0_2_rev_T_7 | _GEN_2462; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_11_i_mux_bus_0_2_rev_T_12 = {{3'd0}, MuxWrapper_11_Omuxes_0_2[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_11_i_mux_bus_0_2_rev_T_14 = {{1'd0}, _FDPE_11_i_mux_bus_0_2_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2464 = {{2'd0}, _FDPE_11_i_mux_bus_0_2_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_11_Omuxes_0_3 = MuxesWrapper_11_io_Omuxes_0_3; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_11_i_mux_bus_0_3_rev_T_2 = {MuxWrapper_11_Omuxes_0_3[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_11_i_mux_bus_0_3_rev_T_4 = {{1'd0}, MuxWrapper_11_Omuxes_0_3[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2466 = {_FDPE_11_i_mux_bus_0_3_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_11_i_mux_bus_0_3_rev_T_6 = {{1'd0}, _GEN_2466}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_11_i_mux_bus_0_3_rev_T_7 = _FDPE_11_i_mux_bus_0_3_rev_T_2 | _FDPE_11_i_mux_bus_0_3_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_11_i_mux_bus_0_3_rev_T_8 = {{2'd0}, MuxWrapper_11_Omuxes_0_3[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_11_i_mux_bus_0_3_rev_T_10 = {_FDPE_11_i_mux_bus_0_3_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2468 = {{2'd0}, _FDPE_11_i_mux_bus_0_3_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_11_i_mux_bus_0_3_rev_T_11 = _FDPE_11_i_mux_bus_0_3_rev_T_7 | _GEN_2468; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_11_i_mux_bus_0_3_rev_T_12 = {{3'd0}, MuxWrapper_11_Omuxes_0_3[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_11_i_mux_bus_0_3_rev_T_14 = {{1'd0}, _FDPE_11_i_mux_bus_0_3_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2470 = {{2'd0}, _FDPE_11_i_mux_bus_0_3_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_11_Omuxes_1_0 = MuxesWrapper_11_io_Omuxes_1_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_11_i_mux_bus_1_0_rev_T_2 = {MuxWrapper_11_Omuxes_1_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_11_i_mux_bus_1_0_rev_T_4 = {{1'd0}, MuxWrapper_11_Omuxes_1_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2472 = {_FDPE_11_i_mux_bus_1_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_11_i_mux_bus_1_0_rev_T_6 = {{1'd0}, _GEN_2472}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_11_i_mux_bus_1_0_rev_T_7 = _FDPE_11_i_mux_bus_1_0_rev_T_2 | _FDPE_11_i_mux_bus_1_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_11_i_mux_bus_1_0_rev_T_8 = {{2'd0}, MuxWrapper_11_Omuxes_1_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_11_i_mux_bus_1_0_rev_T_10 = {_FDPE_11_i_mux_bus_1_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2474 = {{2'd0}, _FDPE_11_i_mux_bus_1_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_11_i_mux_bus_1_0_rev_T_11 = _FDPE_11_i_mux_bus_1_0_rev_T_7 | _GEN_2474; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_11_i_mux_bus_1_0_rev_T_12 = {{3'd0}, MuxWrapper_11_Omuxes_1_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_11_i_mux_bus_1_0_rev_T_14 = {{1'd0}, _FDPE_11_i_mux_bus_1_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2476 = {{2'd0}, _FDPE_11_i_mux_bus_1_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_11_Omuxes_1_1 = MuxesWrapper_11_io_Omuxes_1_1; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_11_i_mux_bus_1_1_rev_T_2 = {MuxWrapper_11_Omuxes_1_1[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_11_i_mux_bus_1_1_rev_T_4 = {{1'd0}, MuxWrapper_11_Omuxes_1_1[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2478 = {_FDPE_11_i_mux_bus_1_1_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_11_i_mux_bus_1_1_rev_T_6 = {{1'd0}, _GEN_2478}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_11_i_mux_bus_1_1_rev_T_7 = _FDPE_11_i_mux_bus_1_1_rev_T_2 | _FDPE_11_i_mux_bus_1_1_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_11_i_mux_bus_1_1_rev_T_8 = {{2'd0}, MuxWrapper_11_Omuxes_1_1[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_11_i_mux_bus_1_1_rev_T_10 = {_FDPE_11_i_mux_bus_1_1_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2480 = {{2'd0}, _FDPE_11_i_mux_bus_1_1_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_11_i_mux_bus_1_1_rev_T_11 = _FDPE_11_i_mux_bus_1_1_rev_T_7 | _GEN_2480; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_11_i_mux_bus_1_1_rev_T_12 = {{3'd0}, MuxWrapper_11_Omuxes_1_1[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_11_i_mux_bus_1_1_rev_T_14 = {{1'd0}, _FDPE_11_i_mux_bus_1_1_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2482 = {{2'd0}, _FDPE_11_i_mux_bus_1_1_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_11_Omuxes_1_2 = MuxesWrapper_11_io_Omuxes_1_2; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_11_i_mux_bus_1_2_rev_T_2 = {MuxWrapper_11_Omuxes_1_2[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_11_i_mux_bus_1_2_rev_T_4 = {{1'd0}, MuxWrapper_11_Omuxes_1_2[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2484 = {_FDPE_11_i_mux_bus_1_2_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_11_i_mux_bus_1_2_rev_T_6 = {{1'd0}, _GEN_2484}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_11_i_mux_bus_1_2_rev_T_7 = _FDPE_11_i_mux_bus_1_2_rev_T_2 | _FDPE_11_i_mux_bus_1_2_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_11_i_mux_bus_1_2_rev_T_8 = {{2'd0}, MuxWrapper_11_Omuxes_1_2[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_11_i_mux_bus_1_2_rev_T_10 = {_FDPE_11_i_mux_bus_1_2_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2486 = {{2'd0}, _FDPE_11_i_mux_bus_1_2_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_11_i_mux_bus_1_2_rev_T_11 = _FDPE_11_i_mux_bus_1_2_rev_T_7 | _GEN_2486; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_11_i_mux_bus_1_2_rev_T_12 = {{3'd0}, MuxWrapper_11_Omuxes_1_2[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_11_i_mux_bus_1_2_rev_T_14 = {{1'd0}, _FDPE_11_i_mux_bus_1_2_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2488 = {{2'd0}, _FDPE_11_i_mux_bus_1_2_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_11_Omuxes_2_0 = MuxesWrapper_11_io_Omuxes_2_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_11_i_mux_bus_2_0_rev_T_2 = {MuxWrapper_11_Omuxes_2_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_11_i_mux_bus_2_0_rev_T_4 = {{1'd0}, MuxWrapper_11_Omuxes_2_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2490 = {_FDPE_11_i_mux_bus_2_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_11_i_mux_bus_2_0_rev_T_6 = {{1'd0}, _GEN_2490}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_11_i_mux_bus_2_0_rev_T_7 = _FDPE_11_i_mux_bus_2_0_rev_T_2 | _FDPE_11_i_mux_bus_2_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_11_i_mux_bus_2_0_rev_T_8 = {{2'd0}, MuxWrapper_11_Omuxes_2_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_11_i_mux_bus_2_0_rev_T_10 = {_FDPE_11_i_mux_bus_2_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2492 = {{2'd0}, _FDPE_11_i_mux_bus_2_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_11_i_mux_bus_2_0_rev_T_11 = _FDPE_11_i_mux_bus_2_0_rev_T_7 | _GEN_2492; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_11_i_mux_bus_2_0_rev_T_12 = {{3'd0}, MuxWrapper_11_Omuxes_2_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_11_i_mux_bus_2_0_rev_T_14 = {{1'd0}, _FDPE_11_i_mux_bus_2_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2494 = {{2'd0}, _FDPE_11_i_mux_bus_2_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_11_Omuxes_2_1 = MuxesWrapper_11_io_Omuxes_2_1; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_11_i_mux_bus_2_1_rev_T_2 = {MuxWrapper_11_Omuxes_2_1[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_11_i_mux_bus_2_1_rev_T_4 = {{1'd0}, MuxWrapper_11_Omuxes_2_1[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2496 = {_FDPE_11_i_mux_bus_2_1_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_11_i_mux_bus_2_1_rev_T_6 = {{1'd0}, _GEN_2496}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_11_i_mux_bus_2_1_rev_T_7 = _FDPE_11_i_mux_bus_2_1_rev_T_2 | _FDPE_11_i_mux_bus_2_1_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_11_i_mux_bus_2_1_rev_T_8 = {{2'd0}, MuxWrapper_11_Omuxes_2_1[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_11_i_mux_bus_2_1_rev_T_10 = {_FDPE_11_i_mux_bus_2_1_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2498 = {{2'd0}, _FDPE_11_i_mux_bus_2_1_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_11_i_mux_bus_2_1_rev_T_11 = _FDPE_11_i_mux_bus_2_1_rev_T_7 | _GEN_2498; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_11_i_mux_bus_2_1_rev_T_12 = {{3'd0}, MuxWrapper_11_Omuxes_2_1[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_11_i_mux_bus_2_1_rev_T_14 = {{1'd0}, _FDPE_11_i_mux_bus_2_1_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2500 = {{2'd0}, _FDPE_11_i_mux_bus_2_1_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_11_Omuxes_3_0 = MuxesWrapper_11_io_Omuxes_3_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_11_i_mux_bus_3_0_rev_T_2 = {MuxWrapper_11_Omuxes_3_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_11_i_mux_bus_3_0_rev_T_4 = {{1'd0}, MuxWrapper_11_Omuxes_3_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2502 = {_FDPE_11_i_mux_bus_3_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_11_i_mux_bus_3_0_rev_T_6 = {{1'd0}, _GEN_2502}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_11_i_mux_bus_3_0_rev_T_7 = _FDPE_11_i_mux_bus_3_0_rev_T_2 | _FDPE_11_i_mux_bus_3_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_11_i_mux_bus_3_0_rev_T_8 = {{2'd0}, MuxWrapper_11_Omuxes_3_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_11_i_mux_bus_3_0_rev_T_10 = {_FDPE_11_i_mux_bus_3_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2504 = {{2'd0}, _FDPE_11_i_mux_bus_3_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_11_i_mux_bus_3_0_rev_T_11 = _FDPE_11_i_mux_bus_3_0_rev_T_7 | _GEN_2504; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_11_i_mux_bus_3_0_rev_T_12 = {{3'd0}, MuxWrapper_11_Omuxes_3_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_11_i_mux_bus_3_0_rev_T_14 = {{1'd0}, _FDPE_11_i_mux_bus_3_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2506 = {{2'd0}, _FDPE_11_i_mux_bus_3_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_12_Omuxes_0_0 = MuxesWrapper_12_io_Omuxes_0_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_12_i_mux_bus_0_0_rev_T_2 = {MuxWrapper_12_Omuxes_0_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_12_i_mux_bus_0_0_rev_T_4 = {{1'd0}, MuxWrapper_12_Omuxes_0_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2508 = {_FDPE_12_i_mux_bus_0_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_12_i_mux_bus_0_0_rev_T_6 = {{1'd0}, _GEN_2508}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_12_i_mux_bus_0_0_rev_T_7 = _FDPE_12_i_mux_bus_0_0_rev_T_2 | _FDPE_12_i_mux_bus_0_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_12_i_mux_bus_0_0_rev_T_8 = {{2'd0}, MuxWrapper_12_Omuxes_0_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_12_i_mux_bus_0_0_rev_T_10 = {_FDPE_12_i_mux_bus_0_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2510 = {{2'd0}, _FDPE_12_i_mux_bus_0_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_12_i_mux_bus_0_0_rev_T_11 = _FDPE_12_i_mux_bus_0_0_rev_T_7 | _GEN_2510; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_12_i_mux_bus_0_0_rev_T_12 = {{3'd0}, MuxWrapper_12_Omuxes_0_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_12_i_mux_bus_0_0_rev_T_14 = {{1'd0}, _FDPE_12_i_mux_bus_0_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2512 = {{2'd0}, _FDPE_12_i_mux_bus_0_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_12_Omuxes_0_1 = MuxesWrapper_12_io_Omuxes_0_1; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_12_i_mux_bus_0_1_rev_T_2 = {MuxWrapper_12_Omuxes_0_1[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_12_i_mux_bus_0_1_rev_T_4 = {{1'd0}, MuxWrapper_12_Omuxes_0_1[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2514 = {_FDPE_12_i_mux_bus_0_1_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_12_i_mux_bus_0_1_rev_T_6 = {{1'd0}, _GEN_2514}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_12_i_mux_bus_0_1_rev_T_7 = _FDPE_12_i_mux_bus_0_1_rev_T_2 | _FDPE_12_i_mux_bus_0_1_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_12_i_mux_bus_0_1_rev_T_8 = {{2'd0}, MuxWrapper_12_Omuxes_0_1[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_12_i_mux_bus_0_1_rev_T_10 = {_FDPE_12_i_mux_bus_0_1_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2516 = {{2'd0}, _FDPE_12_i_mux_bus_0_1_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_12_i_mux_bus_0_1_rev_T_11 = _FDPE_12_i_mux_bus_0_1_rev_T_7 | _GEN_2516; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_12_i_mux_bus_0_1_rev_T_12 = {{3'd0}, MuxWrapper_12_Omuxes_0_1[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_12_i_mux_bus_0_1_rev_T_14 = {{1'd0}, _FDPE_12_i_mux_bus_0_1_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2518 = {{2'd0}, _FDPE_12_i_mux_bus_0_1_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_12_Omuxes_0_2 = MuxesWrapper_12_io_Omuxes_0_2; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_12_i_mux_bus_0_2_rev_T_2 = {MuxWrapper_12_Omuxes_0_2[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_12_i_mux_bus_0_2_rev_T_4 = {{1'd0}, MuxWrapper_12_Omuxes_0_2[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2520 = {_FDPE_12_i_mux_bus_0_2_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_12_i_mux_bus_0_2_rev_T_6 = {{1'd0}, _GEN_2520}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_12_i_mux_bus_0_2_rev_T_7 = _FDPE_12_i_mux_bus_0_2_rev_T_2 | _FDPE_12_i_mux_bus_0_2_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_12_i_mux_bus_0_2_rev_T_8 = {{2'd0}, MuxWrapper_12_Omuxes_0_2[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_12_i_mux_bus_0_2_rev_T_10 = {_FDPE_12_i_mux_bus_0_2_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2522 = {{2'd0}, _FDPE_12_i_mux_bus_0_2_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_12_i_mux_bus_0_2_rev_T_11 = _FDPE_12_i_mux_bus_0_2_rev_T_7 | _GEN_2522; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_12_i_mux_bus_0_2_rev_T_12 = {{3'd0}, MuxWrapper_12_Omuxes_0_2[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_12_i_mux_bus_0_2_rev_T_14 = {{1'd0}, _FDPE_12_i_mux_bus_0_2_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2524 = {{2'd0}, _FDPE_12_i_mux_bus_0_2_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_12_Omuxes_0_3 = MuxesWrapper_12_io_Omuxes_0_3; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_12_i_mux_bus_0_3_rev_T_2 = {MuxWrapper_12_Omuxes_0_3[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_12_i_mux_bus_0_3_rev_T_4 = {{1'd0}, MuxWrapper_12_Omuxes_0_3[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2526 = {_FDPE_12_i_mux_bus_0_3_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_12_i_mux_bus_0_3_rev_T_6 = {{1'd0}, _GEN_2526}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_12_i_mux_bus_0_3_rev_T_7 = _FDPE_12_i_mux_bus_0_3_rev_T_2 | _FDPE_12_i_mux_bus_0_3_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_12_i_mux_bus_0_3_rev_T_8 = {{2'd0}, MuxWrapper_12_Omuxes_0_3[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_12_i_mux_bus_0_3_rev_T_10 = {_FDPE_12_i_mux_bus_0_3_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2528 = {{2'd0}, _FDPE_12_i_mux_bus_0_3_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_12_i_mux_bus_0_3_rev_T_11 = _FDPE_12_i_mux_bus_0_3_rev_T_7 | _GEN_2528; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_12_i_mux_bus_0_3_rev_T_12 = {{3'd0}, MuxWrapper_12_Omuxes_0_3[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_12_i_mux_bus_0_3_rev_T_14 = {{1'd0}, _FDPE_12_i_mux_bus_0_3_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2530 = {{2'd0}, _FDPE_12_i_mux_bus_0_3_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_12_Omuxes_1_0 = MuxesWrapper_12_io_Omuxes_1_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_12_i_mux_bus_1_0_rev_T_2 = {MuxWrapper_12_Omuxes_1_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_12_i_mux_bus_1_0_rev_T_4 = {{1'd0}, MuxWrapper_12_Omuxes_1_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2532 = {_FDPE_12_i_mux_bus_1_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_12_i_mux_bus_1_0_rev_T_6 = {{1'd0}, _GEN_2532}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_12_i_mux_bus_1_0_rev_T_7 = _FDPE_12_i_mux_bus_1_0_rev_T_2 | _FDPE_12_i_mux_bus_1_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_12_i_mux_bus_1_0_rev_T_8 = {{2'd0}, MuxWrapper_12_Omuxes_1_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_12_i_mux_bus_1_0_rev_T_10 = {_FDPE_12_i_mux_bus_1_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2534 = {{2'd0}, _FDPE_12_i_mux_bus_1_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_12_i_mux_bus_1_0_rev_T_11 = _FDPE_12_i_mux_bus_1_0_rev_T_7 | _GEN_2534; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_12_i_mux_bus_1_0_rev_T_12 = {{3'd0}, MuxWrapper_12_Omuxes_1_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_12_i_mux_bus_1_0_rev_T_14 = {{1'd0}, _FDPE_12_i_mux_bus_1_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2536 = {{2'd0}, _FDPE_12_i_mux_bus_1_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_12_Omuxes_1_1 = MuxesWrapper_12_io_Omuxes_1_1; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_12_i_mux_bus_1_1_rev_T_2 = {MuxWrapper_12_Omuxes_1_1[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_12_i_mux_bus_1_1_rev_T_4 = {{1'd0}, MuxWrapper_12_Omuxes_1_1[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2538 = {_FDPE_12_i_mux_bus_1_1_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_12_i_mux_bus_1_1_rev_T_6 = {{1'd0}, _GEN_2538}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_12_i_mux_bus_1_1_rev_T_7 = _FDPE_12_i_mux_bus_1_1_rev_T_2 | _FDPE_12_i_mux_bus_1_1_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_12_i_mux_bus_1_1_rev_T_8 = {{2'd0}, MuxWrapper_12_Omuxes_1_1[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_12_i_mux_bus_1_1_rev_T_10 = {_FDPE_12_i_mux_bus_1_1_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2540 = {{2'd0}, _FDPE_12_i_mux_bus_1_1_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_12_i_mux_bus_1_1_rev_T_11 = _FDPE_12_i_mux_bus_1_1_rev_T_7 | _GEN_2540; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_12_i_mux_bus_1_1_rev_T_12 = {{3'd0}, MuxWrapper_12_Omuxes_1_1[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_12_i_mux_bus_1_1_rev_T_14 = {{1'd0}, _FDPE_12_i_mux_bus_1_1_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2542 = {{2'd0}, _FDPE_12_i_mux_bus_1_1_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_12_Omuxes_1_2 = MuxesWrapper_12_io_Omuxes_1_2; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_12_i_mux_bus_1_2_rev_T_2 = {MuxWrapper_12_Omuxes_1_2[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_12_i_mux_bus_1_2_rev_T_4 = {{1'd0}, MuxWrapper_12_Omuxes_1_2[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2544 = {_FDPE_12_i_mux_bus_1_2_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_12_i_mux_bus_1_2_rev_T_6 = {{1'd0}, _GEN_2544}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_12_i_mux_bus_1_2_rev_T_7 = _FDPE_12_i_mux_bus_1_2_rev_T_2 | _FDPE_12_i_mux_bus_1_2_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_12_i_mux_bus_1_2_rev_T_8 = {{2'd0}, MuxWrapper_12_Omuxes_1_2[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_12_i_mux_bus_1_2_rev_T_10 = {_FDPE_12_i_mux_bus_1_2_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2546 = {{2'd0}, _FDPE_12_i_mux_bus_1_2_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_12_i_mux_bus_1_2_rev_T_11 = _FDPE_12_i_mux_bus_1_2_rev_T_7 | _GEN_2546; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_12_i_mux_bus_1_2_rev_T_12 = {{3'd0}, MuxWrapper_12_Omuxes_1_2[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_12_i_mux_bus_1_2_rev_T_14 = {{1'd0}, _FDPE_12_i_mux_bus_1_2_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2548 = {{2'd0}, _FDPE_12_i_mux_bus_1_2_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_12_Omuxes_2_0 = MuxesWrapper_12_io_Omuxes_2_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_12_i_mux_bus_2_0_rev_T_2 = {MuxWrapper_12_Omuxes_2_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_12_i_mux_bus_2_0_rev_T_4 = {{1'd0}, MuxWrapper_12_Omuxes_2_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2550 = {_FDPE_12_i_mux_bus_2_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_12_i_mux_bus_2_0_rev_T_6 = {{1'd0}, _GEN_2550}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_12_i_mux_bus_2_0_rev_T_7 = _FDPE_12_i_mux_bus_2_0_rev_T_2 | _FDPE_12_i_mux_bus_2_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_12_i_mux_bus_2_0_rev_T_8 = {{2'd0}, MuxWrapper_12_Omuxes_2_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_12_i_mux_bus_2_0_rev_T_10 = {_FDPE_12_i_mux_bus_2_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2552 = {{2'd0}, _FDPE_12_i_mux_bus_2_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_12_i_mux_bus_2_0_rev_T_11 = _FDPE_12_i_mux_bus_2_0_rev_T_7 | _GEN_2552; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_12_i_mux_bus_2_0_rev_T_12 = {{3'd0}, MuxWrapper_12_Omuxes_2_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_12_i_mux_bus_2_0_rev_T_14 = {{1'd0}, _FDPE_12_i_mux_bus_2_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2554 = {{2'd0}, _FDPE_12_i_mux_bus_2_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_12_Omuxes_2_1 = MuxesWrapper_12_io_Omuxes_2_1; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_12_i_mux_bus_2_1_rev_T_2 = {MuxWrapper_12_Omuxes_2_1[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_12_i_mux_bus_2_1_rev_T_4 = {{1'd0}, MuxWrapper_12_Omuxes_2_1[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2556 = {_FDPE_12_i_mux_bus_2_1_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_12_i_mux_bus_2_1_rev_T_6 = {{1'd0}, _GEN_2556}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_12_i_mux_bus_2_1_rev_T_7 = _FDPE_12_i_mux_bus_2_1_rev_T_2 | _FDPE_12_i_mux_bus_2_1_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_12_i_mux_bus_2_1_rev_T_8 = {{2'd0}, MuxWrapper_12_Omuxes_2_1[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_12_i_mux_bus_2_1_rev_T_10 = {_FDPE_12_i_mux_bus_2_1_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2558 = {{2'd0}, _FDPE_12_i_mux_bus_2_1_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_12_i_mux_bus_2_1_rev_T_11 = _FDPE_12_i_mux_bus_2_1_rev_T_7 | _GEN_2558; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_12_i_mux_bus_2_1_rev_T_12 = {{3'd0}, MuxWrapper_12_Omuxes_2_1[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_12_i_mux_bus_2_1_rev_T_14 = {{1'd0}, _FDPE_12_i_mux_bus_2_1_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2560 = {{2'd0}, _FDPE_12_i_mux_bus_2_1_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_12_Omuxes_3_0 = MuxesWrapper_12_io_Omuxes_3_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_12_i_mux_bus_3_0_rev_T_2 = {MuxWrapper_12_Omuxes_3_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_12_i_mux_bus_3_0_rev_T_4 = {{1'd0}, MuxWrapper_12_Omuxes_3_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2562 = {_FDPE_12_i_mux_bus_3_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_12_i_mux_bus_3_0_rev_T_6 = {{1'd0}, _GEN_2562}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_12_i_mux_bus_3_0_rev_T_7 = _FDPE_12_i_mux_bus_3_0_rev_T_2 | _FDPE_12_i_mux_bus_3_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_12_i_mux_bus_3_0_rev_T_8 = {{2'd0}, MuxWrapper_12_Omuxes_3_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_12_i_mux_bus_3_0_rev_T_10 = {_FDPE_12_i_mux_bus_3_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2564 = {{2'd0}, _FDPE_12_i_mux_bus_3_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_12_i_mux_bus_3_0_rev_T_11 = _FDPE_12_i_mux_bus_3_0_rev_T_7 | _GEN_2564; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_12_i_mux_bus_3_0_rev_T_12 = {{3'd0}, MuxWrapper_12_Omuxes_3_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_12_i_mux_bus_3_0_rev_T_14 = {{1'd0}, _FDPE_12_i_mux_bus_3_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2566 = {{2'd0}, _FDPE_12_i_mux_bus_3_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_13_Omuxes_0_0 = MuxesWrapper_13_io_Omuxes_0_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_13_i_mux_bus_0_0_rev_T_2 = {MuxWrapper_13_Omuxes_0_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_13_i_mux_bus_0_0_rev_T_4 = {{1'd0}, MuxWrapper_13_Omuxes_0_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2568 = {_FDPE_13_i_mux_bus_0_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_13_i_mux_bus_0_0_rev_T_6 = {{1'd0}, _GEN_2568}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_13_i_mux_bus_0_0_rev_T_7 = _FDPE_13_i_mux_bus_0_0_rev_T_2 | _FDPE_13_i_mux_bus_0_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_13_i_mux_bus_0_0_rev_T_8 = {{2'd0}, MuxWrapper_13_Omuxes_0_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_13_i_mux_bus_0_0_rev_T_10 = {_FDPE_13_i_mux_bus_0_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2570 = {{2'd0}, _FDPE_13_i_mux_bus_0_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_13_i_mux_bus_0_0_rev_T_11 = _FDPE_13_i_mux_bus_0_0_rev_T_7 | _GEN_2570; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_13_i_mux_bus_0_0_rev_T_12 = {{3'd0}, MuxWrapper_13_Omuxes_0_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_13_i_mux_bus_0_0_rev_T_14 = {{1'd0}, _FDPE_13_i_mux_bus_0_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2572 = {{2'd0}, _FDPE_13_i_mux_bus_0_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_13_Omuxes_0_1 = MuxesWrapper_13_io_Omuxes_0_1; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_13_i_mux_bus_0_1_rev_T_2 = {MuxWrapper_13_Omuxes_0_1[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_13_i_mux_bus_0_1_rev_T_4 = {{1'd0}, MuxWrapper_13_Omuxes_0_1[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2574 = {_FDPE_13_i_mux_bus_0_1_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_13_i_mux_bus_0_1_rev_T_6 = {{1'd0}, _GEN_2574}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_13_i_mux_bus_0_1_rev_T_7 = _FDPE_13_i_mux_bus_0_1_rev_T_2 | _FDPE_13_i_mux_bus_0_1_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_13_i_mux_bus_0_1_rev_T_8 = {{2'd0}, MuxWrapper_13_Omuxes_0_1[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_13_i_mux_bus_0_1_rev_T_10 = {_FDPE_13_i_mux_bus_0_1_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2576 = {{2'd0}, _FDPE_13_i_mux_bus_0_1_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_13_i_mux_bus_0_1_rev_T_11 = _FDPE_13_i_mux_bus_0_1_rev_T_7 | _GEN_2576; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_13_i_mux_bus_0_1_rev_T_12 = {{3'd0}, MuxWrapper_13_Omuxes_0_1[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_13_i_mux_bus_0_1_rev_T_14 = {{1'd0}, _FDPE_13_i_mux_bus_0_1_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2578 = {{2'd0}, _FDPE_13_i_mux_bus_0_1_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_13_Omuxes_0_2 = MuxesWrapper_13_io_Omuxes_0_2; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_13_i_mux_bus_0_2_rev_T_2 = {MuxWrapper_13_Omuxes_0_2[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_13_i_mux_bus_0_2_rev_T_4 = {{1'd0}, MuxWrapper_13_Omuxes_0_2[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2580 = {_FDPE_13_i_mux_bus_0_2_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_13_i_mux_bus_0_2_rev_T_6 = {{1'd0}, _GEN_2580}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_13_i_mux_bus_0_2_rev_T_7 = _FDPE_13_i_mux_bus_0_2_rev_T_2 | _FDPE_13_i_mux_bus_0_2_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_13_i_mux_bus_0_2_rev_T_8 = {{2'd0}, MuxWrapper_13_Omuxes_0_2[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_13_i_mux_bus_0_2_rev_T_10 = {_FDPE_13_i_mux_bus_0_2_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2582 = {{2'd0}, _FDPE_13_i_mux_bus_0_2_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_13_i_mux_bus_0_2_rev_T_11 = _FDPE_13_i_mux_bus_0_2_rev_T_7 | _GEN_2582; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_13_i_mux_bus_0_2_rev_T_12 = {{3'd0}, MuxWrapper_13_Omuxes_0_2[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_13_i_mux_bus_0_2_rev_T_14 = {{1'd0}, _FDPE_13_i_mux_bus_0_2_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2584 = {{2'd0}, _FDPE_13_i_mux_bus_0_2_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_13_Omuxes_0_3 = MuxesWrapper_13_io_Omuxes_0_3; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_13_i_mux_bus_0_3_rev_T_2 = {MuxWrapper_13_Omuxes_0_3[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_13_i_mux_bus_0_3_rev_T_4 = {{1'd0}, MuxWrapper_13_Omuxes_0_3[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2586 = {_FDPE_13_i_mux_bus_0_3_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_13_i_mux_bus_0_3_rev_T_6 = {{1'd0}, _GEN_2586}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_13_i_mux_bus_0_3_rev_T_7 = _FDPE_13_i_mux_bus_0_3_rev_T_2 | _FDPE_13_i_mux_bus_0_3_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_13_i_mux_bus_0_3_rev_T_8 = {{2'd0}, MuxWrapper_13_Omuxes_0_3[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_13_i_mux_bus_0_3_rev_T_10 = {_FDPE_13_i_mux_bus_0_3_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2588 = {{2'd0}, _FDPE_13_i_mux_bus_0_3_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_13_i_mux_bus_0_3_rev_T_11 = _FDPE_13_i_mux_bus_0_3_rev_T_7 | _GEN_2588; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_13_i_mux_bus_0_3_rev_T_12 = {{3'd0}, MuxWrapper_13_Omuxes_0_3[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_13_i_mux_bus_0_3_rev_T_14 = {{1'd0}, _FDPE_13_i_mux_bus_0_3_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2590 = {{2'd0}, _FDPE_13_i_mux_bus_0_3_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_13_Omuxes_1_0 = MuxesWrapper_13_io_Omuxes_1_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_13_i_mux_bus_1_0_rev_T_2 = {MuxWrapper_13_Omuxes_1_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_13_i_mux_bus_1_0_rev_T_4 = {{1'd0}, MuxWrapper_13_Omuxes_1_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2592 = {_FDPE_13_i_mux_bus_1_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_13_i_mux_bus_1_0_rev_T_6 = {{1'd0}, _GEN_2592}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_13_i_mux_bus_1_0_rev_T_7 = _FDPE_13_i_mux_bus_1_0_rev_T_2 | _FDPE_13_i_mux_bus_1_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_13_i_mux_bus_1_0_rev_T_8 = {{2'd0}, MuxWrapper_13_Omuxes_1_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_13_i_mux_bus_1_0_rev_T_10 = {_FDPE_13_i_mux_bus_1_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2594 = {{2'd0}, _FDPE_13_i_mux_bus_1_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_13_i_mux_bus_1_0_rev_T_11 = _FDPE_13_i_mux_bus_1_0_rev_T_7 | _GEN_2594; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_13_i_mux_bus_1_0_rev_T_12 = {{3'd0}, MuxWrapper_13_Omuxes_1_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_13_i_mux_bus_1_0_rev_T_14 = {{1'd0}, _FDPE_13_i_mux_bus_1_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2596 = {{2'd0}, _FDPE_13_i_mux_bus_1_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_13_Omuxes_1_1 = MuxesWrapper_13_io_Omuxes_1_1; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_13_i_mux_bus_1_1_rev_T_2 = {MuxWrapper_13_Omuxes_1_1[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_13_i_mux_bus_1_1_rev_T_4 = {{1'd0}, MuxWrapper_13_Omuxes_1_1[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2598 = {_FDPE_13_i_mux_bus_1_1_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_13_i_mux_bus_1_1_rev_T_6 = {{1'd0}, _GEN_2598}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_13_i_mux_bus_1_1_rev_T_7 = _FDPE_13_i_mux_bus_1_1_rev_T_2 | _FDPE_13_i_mux_bus_1_1_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_13_i_mux_bus_1_1_rev_T_8 = {{2'd0}, MuxWrapper_13_Omuxes_1_1[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_13_i_mux_bus_1_1_rev_T_10 = {_FDPE_13_i_mux_bus_1_1_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2600 = {{2'd0}, _FDPE_13_i_mux_bus_1_1_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_13_i_mux_bus_1_1_rev_T_11 = _FDPE_13_i_mux_bus_1_1_rev_T_7 | _GEN_2600; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_13_i_mux_bus_1_1_rev_T_12 = {{3'd0}, MuxWrapper_13_Omuxes_1_1[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_13_i_mux_bus_1_1_rev_T_14 = {{1'd0}, _FDPE_13_i_mux_bus_1_1_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2602 = {{2'd0}, _FDPE_13_i_mux_bus_1_1_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_13_Omuxes_1_2 = MuxesWrapper_13_io_Omuxes_1_2; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_13_i_mux_bus_1_2_rev_T_2 = {MuxWrapper_13_Omuxes_1_2[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_13_i_mux_bus_1_2_rev_T_4 = {{1'd0}, MuxWrapper_13_Omuxes_1_2[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2604 = {_FDPE_13_i_mux_bus_1_2_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_13_i_mux_bus_1_2_rev_T_6 = {{1'd0}, _GEN_2604}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_13_i_mux_bus_1_2_rev_T_7 = _FDPE_13_i_mux_bus_1_2_rev_T_2 | _FDPE_13_i_mux_bus_1_2_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_13_i_mux_bus_1_2_rev_T_8 = {{2'd0}, MuxWrapper_13_Omuxes_1_2[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_13_i_mux_bus_1_2_rev_T_10 = {_FDPE_13_i_mux_bus_1_2_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2606 = {{2'd0}, _FDPE_13_i_mux_bus_1_2_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_13_i_mux_bus_1_2_rev_T_11 = _FDPE_13_i_mux_bus_1_2_rev_T_7 | _GEN_2606; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_13_i_mux_bus_1_2_rev_T_12 = {{3'd0}, MuxWrapper_13_Omuxes_1_2[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_13_i_mux_bus_1_2_rev_T_14 = {{1'd0}, _FDPE_13_i_mux_bus_1_2_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2608 = {{2'd0}, _FDPE_13_i_mux_bus_1_2_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_13_Omuxes_2_0 = MuxesWrapper_13_io_Omuxes_2_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_13_i_mux_bus_2_0_rev_T_2 = {MuxWrapper_13_Omuxes_2_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_13_i_mux_bus_2_0_rev_T_4 = {{1'd0}, MuxWrapper_13_Omuxes_2_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2610 = {_FDPE_13_i_mux_bus_2_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_13_i_mux_bus_2_0_rev_T_6 = {{1'd0}, _GEN_2610}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_13_i_mux_bus_2_0_rev_T_7 = _FDPE_13_i_mux_bus_2_0_rev_T_2 | _FDPE_13_i_mux_bus_2_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_13_i_mux_bus_2_0_rev_T_8 = {{2'd0}, MuxWrapper_13_Omuxes_2_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_13_i_mux_bus_2_0_rev_T_10 = {_FDPE_13_i_mux_bus_2_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2612 = {{2'd0}, _FDPE_13_i_mux_bus_2_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_13_i_mux_bus_2_0_rev_T_11 = _FDPE_13_i_mux_bus_2_0_rev_T_7 | _GEN_2612; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_13_i_mux_bus_2_0_rev_T_12 = {{3'd0}, MuxWrapper_13_Omuxes_2_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_13_i_mux_bus_2_0_rev_T_14 = {{1'd0}, _FDPE_13_i_mux_bus_2_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2614 = {{2'd0}, _FDPE_13_i_mux_bus_2_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_13_Omuxes_2_1 = MuxesWrapper_13_io_Omuxes_2_1; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_13_i_mux_bus_2_1_rev_T_2 = {MuxWrapper_13_Omuxes_2_1[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_13_i_mux_bus_2_1_rev_T_4 = {{1'd0}, MuxWrapper_13_Omuxes_2_1[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2616 = {_FDPE_13_i_mux_bus_2_1_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_13_i_mux_bus_2_1_rev_T_6 = {{1'd0}, _GEN_2616}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_13_i_mux_bus_2_1_rev_T_7 = _FDPE_13_i_mux_bus_2_1_rev_T_2 | _FDPE_13_i_mux_bus_2_1_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_13_i_mux_bus_2_1_rev_T_8 = {{2'd0}, MuxWrapper_13_Omuxes_2_1[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_13_i_mux_bus_2_1_rev_T_10 = {_FDPE_13_i_mux_bus_2_1_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2618 = {{2'd0}, _FDPE_13_i_mux_bus_2_1_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_13_i_mux_bus_2_1_rev_T_11 = _FDPE_13_i_mux_bus_2_1_rev_T_7 | _GEN_2618; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_13_i_mux_bus_2_1_rev_T_12 = {{3'd0}, MuxWrapper_13_Omuxes_2_1[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_13_i_mux_bus_2_1_rev_T_14 = {{1'd0}, _FDPE_13_i_mux_bus_2_1_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2620 = {{2'd0}, _FDPE_13_i_mux_bus_2_1_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_13_Omuxes_3_0 = MuxesWrapper_13_io_Omuxes_3_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_13_i_mux_bus_3_0_rev_T_2 = {MuxWrapper_13_Omuxes_3_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_13_i_mux_bus_3_0_rev_T_4 = {{1'd0}, MuxWrapper_13_Omuxes_3_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2622 = {_FDPE_13_i_mux_bus_3_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_13_i_mux_bus_3_0_rev_T_6 = {{1'd0}, _GEN_2622}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_13_i_mux_bus_3_0_rev_T_7 = _FDPE_13_i_mux_bus_3_0_rev_T_2 | _FDPE_13_i_mux_bus_3_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_13_i_mux_bus_3_0_rev_T_8 = {{2'd0}, MuxWrapper_13_Omuxes_3_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_13_i_mux_bus_3_0_rev_T_10 = {_FDPE_13_i_mux_bus_3_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2624 = {{2'd0}, _FDPE_13_i_mux_bus_3_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_13_i_mux_bus_3_0_rev_T_11 = _FDPE_13_i_mux_bus_3_0_rev_T_7 | _GEN_2624; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_13_i_mux_bus_3_0_rev_T_12 = {{3'd0}, MuxWrapper_13_Omuxes_3_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_13_i_mux_bus_3_0_rev_T_14 = {{1'd0}, _FDPE_13_i_mux_bus_3_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2626 = {{2'd0}, _FDPE_13_i_mux_bus_3_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_14_Omuxes_0_0 = MuxesWrapper_14_io_Omuxes_0_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_14_i_mux_bus_0_0_rev_T_2 = {MuxWrapper_14_Omuxes_0_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_14_i_mux_bus_0_0_rev_T_4 = {{1'd0}, MuxWrapper_14_Omuxes_0_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2628 = {_FDPE_14_i_mux_bus_0_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_14_i_mux_bus_0_0_rev_T_6 = {{1'd0}, _GEN_2628}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_14_i_mux_bus_0_0_rev_T_7 = _FDPE_14_i_mux_bus_0_0_rev_T_2 | _FDPE_14_i_mux_bus_0_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_14_i_mux_bus_0_0_rev_T_8 = {{2'd0}, MuxWrapper_14_Omuxes_0_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_14_i_mux_bus_0_0_rev_T_10 = {_FDPE_14_i_mux_bus_0_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2630 = {{2'd0}, _FDPE_14_i_mux_bus_0_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_14_i_mux_bus_0_0_rev_T_11 = _FDPE_14_i_mux_bus_0_0_rev_T_7 | _GEN_2630; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_14_i_mux_bus_0_0_rev_T_12 = {{3'd0}, MuxWrapper_14_Omuxes_0_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_14_i_mux_bus_0_0_rev_T_14 = {{1'd0}, _FDPE_14_i_mux_bus_0_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2632 = {{2'd0}, _FDPE_14_i_mux_bus_0_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_14_Omuxes_0_1 = MuxesWrapper_14_io_Omuxes_0_1; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_14_i_mux_bus_0_1_rev_T_2 = {MuxWrapper_14_Omuxes_0_1[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_14_i_mux_bus_0_1_rev_T_4 = {{1'd0}, MuxWrapper_14_Omuxes_0_1[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2634 = {_FDPE_14_i_mux_bus_0_1_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_14_i_mux_bus_0_1_rev_T_6 = {{1'd0}, _GEN_2634}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_14_i_mux_bus_0_1_rev_T_7 = _FDPE_14_i_mux_bus_0_1_rev_T_2 | _FDPE_14_i_mux_bus_0_1_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_14_i_mux_bus_0_1_rev_T_8 = {{2'd0}, MuxWrapper_14_Omuxes_0_1[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_14_i_mux_bus_0_1_rev_T_10 = {_FDPE_14_i_mux_bus_0_1_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2636 = {{2'd0}, _FDPE_14_i_mux_bus_0_1_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_14_i_mux_bus_0_1_rev_T_11 = _FDPE_14_i_mux_bus_0_1_rev_T_7 | _GEN_2636; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_14_i_mux_bus_0_1_rev_T_12 = {{3'd0}, MuxWrapper_14_Omuxes_0_1[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_14_i_mux_bus_0_1_rev_T_14 = {{1'd0}, _FDPE_14_i_mux_bus_0_1_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2638 = {{2'd0}, _FDPE_14_i_mux_bus_0_1_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_14_Omuxes_0_2 = MuxesWrapper_14_io_Omuxes_0_2; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_14_i_mux_bus_0_2_rev_T_2 = {MuxWrapper_14_Omuxes_0_2[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_14_i_mux_bus_0_2_rev_T_4 = {{1'd0}, MuxWrapper_14_Omuxes_0_2[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2640 = {_FDPE_14_i_mux_bus_0_2_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_14_i_mux_bus_0_2_rev_T_6 = {{1'd0}, _GEN_2640}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_14_i_mux_bus_0_2_rev_T_7 = _FDPE_14_i_mux_bus_0_2_rev_T_2 | _FDPE_14_i_mux_bus_0_2_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_14_i_mux_bus_0_2_rev_T_8 = {{2'd0}, MuxWrapper_14_Omuxes_0_2[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_14_i_mux_bus_0_2_rev_T_10 = {_FDPE_14_i_mux_bus_0_2_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2642 = {{2'd0}, _FDPE_14_i_mux_bus_0_2_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_14_i_mux_bus_0_2_rev_T_11 = _FDPE_14_i_mux_bus_0_2_rev_T_7 | _GEN_2642; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_14_i_mux_bus_0_2_rev_T_12 = {{3'd0}, MuxWrapper_14_Omuxes_0_2[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_14_i_mux_bus_0_2_rev_T_14 = {{1'd0}, _FDPE_14_i_mux_bus_0_2_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2644 = {{2'd0}, _FDPE_14_i_mux_bus_0_2_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_14_Omuxes_0_3 = MuxesWrapper_14_io_Omuxes_0_3; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_14_i_mux_bus_0_3_rev_T_2 = {MuxWrapper_14_Omuxes_0_3[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_14_i_mux_bus_0_3_rev_T_4 = {{1'd0}, MuxWrapper_14_Omuxes_0_3[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2646 = {_FDPE_14_i_mux_bus_0_3_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_14_i_mux_bus_0_3_rev_T_6 = {{1'd0}, _GEN_2646}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_14_i_mux_bus_0_3_rev_T_7 = _FDPE_14_i_mux_bus_0_3_rev_T_2 | _FDPE_14_i_mux_bus_0_3_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_14_i_mux_bus_0_3_rev_T_8 = {{2'd0}, MuxWrapper_14_Omuxes_0_3[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_14_i_mux_bus_0_3_rev_T_10 = {_FDPE_14_i_mux_bus_0_3_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2648 = {{2'd0}, _FDPE_14_i_mux_bus_0_3_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_14_i_mux_bus_0_3_rev_T_11 = _FDPE_14_i_mux_bus_0_3_rev_T_7 | _GEN_2648; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_14_i_mux_bus_0_3_rev_T_12 = {{3'd0}, MuxWrapper_14_Omuxes_0_3[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_14_i_mux_bus_0_3_rev_T_14 = {{1'd0}, _FDPE_14_i_mux_bus_0_3_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2650 = {{2'd0}, _FDPE_14_i_mux_bus_0_3_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_14_Omuxes_1_0 = MuxesWrapper_14_io_Omuxes_1_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_14_i_mux_bus_1_0_rev_T_2 = {MuxWrapper_14_Omuxes_1_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_14_i_mux_bus_1_0_rev_T_4 = {{1'd0}, MuxWrapper_14_Omuxes_1_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2652 = {_FDPE_14_i_mux_bus_1_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_14_i_mux_bus_1_0_rev_T_6 = {{1'd0}, _GEN_2652}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_14_i_mux_bus_1_0_rev_T_7 = _FDPE_14_i_mux_bus_1_0_rev_T_2 | _FDPE_14_i_mux_bus_1_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_14_i_mux_bus_1_0_rev_T_8 = {{2'd0}, MuxWrapper_14_Omuxes_1_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_14_i_mux_bus_1_0_rev_T_10 = {_FDPE_14_i_mux_bus_1_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2654 = {{2'd0}, _FDPE_14_i_mux_bus_1_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_14_i_mux_bus_1_0_rev_T_11 = _FDPE_14_i_mux_bus_1_0_rev_T_7 | _GEN_2654; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_14_i_mux_bus_1_0_rev_T_12 = {{3'd0}, MuxWrapper_14_Omuxes_1_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_14_i_mux_bus_1_0_rev_T_14 = {{1'd0}, _FDPE_14_i_mux_bus_1_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2656 = {{2'd0}, _FDPE_14_i_mux_bus_1_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_14_Omuxes_1_1 = MuxesWrapper_14_io_Omuxes_1_1; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_14_i_mux_bus_1_1_rev_T_2 = {MuxWrapper_14_Omuxes_1_1[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_14_i_mux_bus_1_1_rev_T_4 = {{1'd0}, MuxWrapper_14_Omuxes_1_1[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2658 = {_FDPE_14_i_mux_bus_1_1_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_14_i_mux_bus_1_1_rev_T_6 = {{1'd0}, _GEN_2658}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_14_i_mux_bus_1_1_rev_T_7 = _FDPE_14_i_mux_bus_1_1_rev_T_2 | _FDPE_14_i_mux_bus_1_1_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_14_i_mux_bus_1_1_rev_T_8 = {{2'd0}, MuxWrapper_14_Omuxes_1_1[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_14_i_mux_bus_1_1_rev_T_10 = {_FDPE_14_i_mux_bus_1_1_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2660 = {{2'd0}, _FDPE_14_i_mux_bus_1_1_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_14_i_mux_bus_1_1_rev_T_11 = _FDPE_14_i_mux_bus_1_1_rev_T_7 | _GEN_2660; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_14_i_mux_bus_1_1_rev_T_12 = {{3'd0}, MuxWrapper_14_Omuxes_1_1[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_14_i_mux_bus_1_1_rev_T_14 = {{1'd0}, _FDPE_14_i_mux_bus_1_1_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2662 = {{2'd0}, _FDPE_14_i_mux_bus_1_1_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_14_Omuxes_1_2 = MuxesWrapper_14_io_Omuxes_1_2; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_14_i_mux_bus_1_2_rev_T_2 = {MuxWrapper_14_Omuxes_1_2[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_14_i_mux_bus_1_2_rev_T_4 = {{1'd0}, MuxWrapper_14_Omuxes_1_2[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2664 = {_FDPE_14_i_mux_bus_1_2_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_14_i_mux_bus_1_2_rev_T_6 = {{1'd0}, _GEN_2664}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_14_i_mux_bus_1_2_rev_T_7 = _FDPE_14_i_mux_bus_1_2_rev_T_2 | _FDPE_14_i_mux_bus_1_2_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_14_i_mux_bus_1_2_rev_T_8 = {{2'd0}, MuxWrapper_14_Omuxes_1_2[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_14_i_mux_bus_1_2_rev_T_10 = {_FDPE_14_i_mux_bus_1_2_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2666 = {{2'd0}, _FDPE_14_i_mux_bus_1_2_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_14_i_mux_bus_1_2_rev_T_11 = _FDPE_14_i_mux_bus_1_2_rev_T_7 | _GEN_2666; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_14_i_mux_bus_1_2_rev_T_12 = {{3'd0}, MuxWrapper_14_Omuxes_1_2[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_14_i_mux_bus_1_2_rev_T_14 = {{1'd0}, _FDPE_14_i_mux_bus_1_2_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2668 = {{2'd0}, _FDPE_14_i_mux_bus_1_2_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_14_Omuxes_2_0 = MuxesWrapper_14_io_Omuxes_2_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_14_i_mux_bus_2_0_rev_T_2 = {MuxWrapper_14_Omuxes_2_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_14_i_mux_bus_2_0_rev_T_4 = {{1'd0}, MuxWrapper_14_Omuxes_2_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2670 = {_FDPE_14_i_mux_bus_2_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_14_i_mux_bus_2_0_rev_T_6 = {{1'd0}, _GEN_2670}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_14_i_mux_bus_2_0_rev_T_7 = _FDPE_14_i_mux_bus_2_0_rev_T_2 | _FDPE_14_i_mux_bus_2_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_14_i_mux_bus_2_0_rev_T_8 = {{2'd0}, MuxWrapper_14_Omuxes_2_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_14_i_mux_bus_2_0_rev_T_10 = {_FDPE_14_i_mux_bus_2_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2672 = {{2'd0}, _FDPE_14_i_mux_bus_2_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_14_i_mux_bus_2_0_rev_T_11 = _FDPE_14_i_mux_bus_2_0_rev_T_7 | _GEN_2672; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_14_i_mux_bus_2_0_rev_T_12 = {{3'd0}, MuxWrapper_14_Omuxes_2_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_14_i_mux_bus_2_0_rev_T_14 = {{1'd0}, _FDPE_14_i_mux_bus_2_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2674 = {{2'd0}, _FDPE_14_i_mux_bus_2_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_14_Omuxes_2_1 = MuxesWrapper_14_io_Omuxes_2_1; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_14_i_mux_bus_2_1_rev_T_2 = {MuxWrapper_14_Omuxes_2_1[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_14_i_mux_bus_2_1_rev_T_4 = {{1'd0}, MuxWrapper_14_Omuxes_2_1[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2676 = {_FDPE_14_i_mux_bus_2_1_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_14_i_mux_bus_2_1_rev_T_6 = {{1'd0}, _GEN_2676}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_14_i_mux_bus_2_1_rev_T_7 = _FDPE_14_i_mux_bus_2_1_rev_T_2 | _FDPE_14_i_mux_bus_2_1_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_14_i_mux_bus_2_1_rev_T_8 = {{2'd0}, MuxWrapper_14_Omuxes_2_1[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_14_i_mux_bus_2_1_rev_T_10 = {_FDPE_14_i_mux_bus_2_1_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2678 = {{2'd0}, _FDPE_14_i_mux_bus_2_1_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_14_i_mux_bus_2_1_rev_T_11 = _FDPE_14_i_mux_bus_2_1_rev_T_7 | _GEN_2678; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_14_i_mux_bus_2_1_rev_T_12 = {{3'd0}, MuxWrapper_14_Omuxes_2_1[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_14_i_mux_bus_2_1_rev_T_14 = {{1'd0}, _FDPE_14_i_mux_bus_2_1_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2680 = {{2'd0}, _FDPE_14_i_mux_bus_2_1_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_14_Omuxes_3_0 = MuxesWrapper_14_io_Omuxes_3_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_14_i_mux_bus_3_0_rev_T_2 = {MuxWrapper_14_Omuxes_3_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_14_i_mux_bus_3_0_rev_T_4 = {{1'd0}, MuxWrapper_14_Omuxes_3_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2682 = {_FDPE_14_i_mux_bus_3_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_14_i_mux_bus_3_0_rev_T_6 = {{1'd0}, _GEN_2682}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_14_i_mux_bus_3_0_rev_T_7 = _FDPE_14_i_mux_bus_3_0_rev_T_2 | _FDPE_14_i_mux_bus_3_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_14_i_mux_bus_3_0_rev_T_8 = {{2'd0}, MuxWrapper_14_Omuxes_3_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_14_i_mux_bus_3_0_rev_T_10 = {_FDPE_14_i_mux_bus_3_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2684 = {{2'd0}, _FDPE_14_i_mux_bus_3_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_14_i_mux_bus_3_0_rev_T_11 = _FDPE_14_i_mux_bus_3_0_rev_T_7 | _GEN_2684; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_14_i_mux_bus_3_0_rev_T_12 = {{3'd0}, MuxWrapper_14_Omuxes_3_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_14_i_mux_bus_3_0_rev_T_14 = {{1'd0}, _FDPE_14_i_mux_bus_3_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2686 = {{2'd0}, _FDPE_14_i_mux_bus_3_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_15_Omuxes_0_0 = MuxesWrapper_15_io_Omuxes_0_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_15_i_mux_bus_0_0_rev_T_2 = {MuxWrapper_15_Omuxes_0_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_15_i_mux_bus_0_0_rev_T_4 = {{1'd0}, MuxWrapper_15_Omuxes_0_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2688 = {_FDPE_15_i_mux_bus_0_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_15_i_mux_bus_0_0_rev_T_6 = {{1'd0}, _GEN_2688}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_15_i_mux_bus_0_0_rev_T_7 = _FDPE_15_i_mux_bus_0_0_rev_T_2 | _FDPE_15_i_mux_bus_0_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_15_i_mux_bus_0_0_rev_T_8 = {{2'd0}, MuxWrapper_15_Omuxes_0_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_15_i_mux_bus_0_0_rev_T_10 = {_FDPE_15_i_mux_bus_0_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2690 = {{2'd0}, _FDPE_15_i_mux_bus_0_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_15_i_mux_bus_0_0_rev_T_11 = _FDPE_15_i_mux_bus_0_0_rev_T_7 | _GEN_2690; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_15_i_mux_bus_0_0_rev_T_12 = {{3'd0}, MuxWrapper_15_Omuxes_0_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_15_i_mux_bus_0_0_rev_T_14 = {{1'd0}, _FDPE_15_i_mux_bus_0_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2692 = {{2'd0}, _FDPE_15_i_mux_bus_0_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_15_Omuxes_0_1 = MuxesWrapper_15_io_Omuxes_0_1; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_15_i_mux_bus_0_1_rev_T_2 = {MuxWrapper_15_Omuxes_0_1[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_15_i_mux_bus_0_1_rev_T_4 = {{1'd0}, MuxWrapper_15_Omuxes_0_1[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2694 = {_FDPE_15_i_mux_bus_0_1_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_15_i_mux_bus_0_1_rev_T_6 = {{1'd0}, _GEN_2694}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_15_i_mux_bus_0_1_rev_T_7 = _FDPE_15_i_mux_bus_0_1_rev_T_2 | _FDPE_15_i_mux_bus_0_1_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_15_i_mux_bus_0_1_rev_T_8 = {{2'd0}, MuxWrapper_15_Omuxes_0_1[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_15_i_mux_bus_0_1_rev_T_10 = {_FDPE_15_i_mux_bus_0_1_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2696 = {{2'd0}, _FDPE_15_i_mux_bus_0_1_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_15_i_mux_bus_0_1_rev_T_11 = _FDPE_15_i_mux_bus_0_1_rev_T_7 | _GEN_2696; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_15_i_mux_bus_0_1_rev_T_12 = {{3'd0}, MuxWrapper_15_Omuxes_0_1[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_15_i_mux_bus_0_1_rev_T_14 = {{1'd0}, _FDPE_15_i_mux_bus_0_1_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2698 = {{2'd0}, _FDPE_15_i_mux_bus_0_1_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_15_Omuxes_0_2 = MuxesWrapper_15_io_Omuxes_0_2; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_15_i_mux_bus_0_2_rev_T_2 = {MuxWrapper_15_Omuxes_0_2[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_15_i_mux_bus_0_2_rev_T_4 = {{1'd0}, MuxWrapper_15_Omuxes_0_2[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2700 = {_FDPE_15_i_mux_bus_0_2_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_15_i_mux_bus_0_2_rev_T_6 = {{1'd0}, _GEN_2700}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_15_i_mux_bus_0_2_rev_T_7 = _FDPE_15_i_mux_bus_0_2_rev_T_2 | _FDPE_15_i_mux_bus_0_2_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_15_i_mux_bus_0_2_rev_T_8 = {{2'd0}, MuxWrapper_15_Omuxes_0_2[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_15_i_mux_bus_0_2_rev_T_10 = {_FDPE_15_i_mux_bus_0_2_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2702 = {{2'd0}, _FDPE_15_i_mux_bus_0_2_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_15_i_mux_bus_0_2_rev_T_11 = _FDPE_15_i_mux_bus_0_2_rev_T_7 | _GEN_2702; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_15_i_mux_bus_0_2_rev_T_12 = {{3'd0}, MuxWrapper_15_Omuxes_0_2[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_15_i_mux_bus_0_2_rev_T_14 = {{1'd0}, _FDPE_15_i_mux_bus_0_2_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2704 = {{2'd0}, _FDPE_15_i_mux_bus_0_2_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_15_Omuxes_0_3 = MuxesWrapper_15_io_Omuxes_0_3; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_15_i_mux_bus_0_3_rev_T_2 = {MuxWrapper_15_Omuxes_0_3[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_15_i_mux_bus_0_3_rev_T_4 = {{1'd0}, MuxWrapper_15_Omuxes_0_3[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2706 = {_FDPE_15_i_mux_bus_0_3_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_15_i_mux_bus_0_3_rev_T_6 = {{1'd0}, _GEN_2706}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_15_i_mux_bus_0_3_rev_T_7 = _FDPE_15_i_mux_bus_0_3_rev_T_2 | _FDPE_15_i_mux_bus_0_3_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_15_i_mux_bus_0_3_rev_T_8 = {{2'd0}, MuxWrapper_15_Omuxes_0_3[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_15_i_mux_bus_0_3_rev_T_10 = {_FDPE_15_i_mux_bus_0_3_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2708 = {{2'd0}, _FDPE_15_i_mux_bus_0_3_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_15_i_mux_bus_0_3_rev_T_11 = _FDPE_15_i_mux_bus_0_3_rev_T_7 | _GEN_2708; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_15_i_mux_bus_0_3_rev_T_12 = {{3'd0}, MuxWrapper_15_Omuxes_0_3[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_15_i_mux_bus_0_3_rev_T_14 = {{1'd0}, _FDPE_15_i_mux_bus_0_3_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2710 = {{2'd0}, _FDPE_15_i_mux_bus_0_3_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_15_Omuxes_1_0 = MuxesWrapper_15_io_Omuxes_1_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_15_i_mux_bus_1_0_rev_T_2 = {MuxWrapper_15_Omuxes_1_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_15_i_mux_bus_1_0_rev_T_4 = {{1'd0}, MuxWrapper_15_Omuxes_1_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2712 = {_FDPE_15_i_mux_bus_1_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_15_i_mux_bus_1_0_rev_T_6 = {{1'd0}, _GEN_2712}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_15_i_mux_bus_1_0_rev_T_7 = _FDPE_15_i_mux_bus_1_0_rev_T_2 | _FDPE_15_i_mux_bus_1_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_15_i_mux_bus_1_0_rev_T_8 = {{2'd0}, MuxWrapper_15_Omuxes_1_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_15_i_mux_bus_1_0_rev_T_10 = {_FDPE_15_i_mux_bus_1_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2714 = {{2'd0}, _FDPE_15_i_mux_bus_1_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_15_i_mux_bus_1_0_rev_T_11 = _FDPE_15_i_mux_bus_1_0_rev_T_7 | _GEN_2714; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_15_i_mux_bus_1_0_rev_T_12 = {{3'd0}, MuxWrapper_15_Omuxes_1_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_15_i_mux_bus_1_0_rev_T_14 = {{1'd0}, _FDPE_15_i_mux_bus_1_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2716 = {{2'd0}, _FDPE_15_i_mux_bus_1_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_15_Omuxes_1_1 = MuxesWrapper_15_io_Omuxes_1_1; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_15_i_mux_bus_1_1_rev_T_2 = {MuxWrapper_15_Omuxes_1_1[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_15_i_mux_bus_1_1_rev_T_4 = {{1'd0}, MuxWrapper_15_Omuxes_1_1[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2718 = {_FDPE_15_i_mux_bus_1_1_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_15_i_mux_bus_1_1_rev_T_6 = {{1'd0}, _GEN_2718}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_15_i_mux_bus_1_1_rev_T_7 = _FDPE_15_i_mux_bus_1_1_rev_T_2 | _FDPE_15_i_mux_bus_1_1_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_15_i_mux_bus_1_1_rev_T_8 = {{2'd0}, MuxWrapper_15_Omuxes_1_1[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_15_i_mux_bus_1_1_rev_T_10 = {_FDPE_15_i_mux_bus_1_1_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2720 = {{2'd0}, _FDPE_15_i_mux_bus_1_1_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_15_i_mux_bus_1_1_rev_T_11 = _FDPE_15_i_mux_bus_1_1_rev_T_7 | _GEN_2720; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_15_i_mux_bus_1_1_rev_T_12 = {{3'd0}, MuxWrapper_15_Omuxes_1_1[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_15_i_mux_bus_1_1_rev_T_14 = {{1'd0}, _FDPE_15_i_mux_bus_1_1_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2722 = {{2'd0}, _FDPE_15_i_mux_bus_1_1_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_15_Omuxes_1_2 = MuxesWrapper_15_io_Omuxes_1_2; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_15_i_mux_bus_1_2_rev_T_2 = {MuxWrapper_15_Omuxes_1_2[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_15_i_mux_bus_1_2_rev_T_4 = {{1'd0}, MuxWrapper_15_Omuxes_1_2[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2724 = {_FDPE_15_i_mux_bus_1_2_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_15_i_mux_bus_1_2_rev_T_6 = {{1'd0}, _GEN_2724}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_15_i_mux_bus_1_2_rev_T_7 = _FDPE_15_i_mux_bus_1_2_rev_T_2 | _FDPE_15_i_mux_bus_1_2_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_15_i_mux_bus_1_2_rev_T_8 = {{2'd0}, MuxWrapper_15_Omuxes_1_2[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_15_i_mux_bus_1_2_rev_T_10 = {_FDPE_15_i_mux_bus_1_2_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2726 = {{2'd0}, _FDPE_15_i_mux_bus_1_2_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_15_i_mux_bus_1_2_rev_T_11 = _FDPE_15_i_mux_bus_1_2_rev_T_7 | _GEN_2726; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_15_i_mux_bus_1_2_rev_T_12 = {{3'd0}, MuxWrapper_15_Omuxes_1_2[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_15_i_mux_bus_1_2_rev_T_14 = {{1'd0}, _FDPE_15_i_mux_bus_1_2_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2728 = {{2'd0}, _FDPE_15_i_mux_bus_1_2_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_15_Omuxes_2_0 = MuxesWrapper_15_io_Omuxes_2_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_15_i_mux_bus_2_0_rev_T_2 = {MuxWrapper_15_Omuxes_2_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_15_i_mux_bus_2_0_rev_T_4 = {{1'd0}, MuxWrapper_15_Omuxes_2_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2730 = {_FDPE_15_i_mux_bus_2_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_15_i_mux_bus_2_0_rev_T_6 = {{1'd0}, _GEN_2730}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_15_i_mux_bus_2_0_rev_T_7 = _FDPE_15_i_mux_bus_2_0_rev_T_2 | _FDPE_15_i_mux_bus_2_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_15_i_mux_bus_2_0_rev_T_8 = {{2'd0}, MuxWrapper_15_Omuxes_2_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_15_i_mux_bus_2_0_rev_T_10 = {_FDPE_15_i_mux_bus_2_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2732 = {{2'd0}, _FDPE_15_i_mux_bus_2_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_15_i_mux_bus_2_0_rev_T_11 = _FDPE_15_i_mux_bus_2_0_rev_T_7 | _GEN_2732; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_15_i_mux_bus_2_0_rev_T_12 = {{3'd0}, MuxWrapper_15_Omuxes_2_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_15_i_mux_bus_2_0_rev_T_14 = {{1'd0}, _FDPE_15_i_mux_bus_2_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2734 = {{2'd0}, _FDPE_15_i_mux_bus_2_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_15_Omuxes_2_1 = MuxesWrapper_15_io_Omuxes_2_1; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_15_i_mux_bus_2_1_rev_T_2 = {MuxWrapper_15_Omuxes_2_1[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_15_i_mux_bus_2_1_rev_T_4 = {{1'd0}, MuxWrapper_15_Omuxes_2_1[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2736 = {_FDPE_15_i_mux_bus_2_1_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_15_i_mux_bus_2_1_rev_T_6 = {{1'd0}, _GEN_2736}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_15_i_mux_bus_2_1_rev_T_7 = _FDPE_15_i_mux_bus_2_1_rev_T_2 | _FDPE_15_i_mux_bus_2_1_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_15_i_mux_bus_2_1_rev_T_8 = {{2'd0}, MuxWrapper_15_Omuxes_2_1[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_15_i_mux_bus_2_1_rev_T_10 = {_FDPE_15_i_mux_bus_2_1_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2738 = {{2'd0}, _FDPE_15_i_mux_bus_2_1_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_15_i_mux_bus_2_1_rev_T_11 = _FDPE_15_i_mux_bus_2_1_rev_T_7 | _GEN_2738; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_15_i_mux_bus_2_1_rev_T_12 = {{3'd0}, MuxWrapper_15_Omuxes_2_1[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_15_i_mux_bus_2_1_rev_T_14 = {{1'd0}, _FDPE_15_i_mux_bus_2_1_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2740 = {{2'd0}, _FDPE_15_i_mux_bus_2_1_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] MuxWrapper_15_Omuxes_3_0 = MuxesWrapper_15_io_Omuxes_3_0; // @[FlexDPU.scala 124:{33,33}]
  wire [3:0] _FDPE_15_i_mux_bus_3_0_rev_T_2 = {MuxWrapper_15_Omuxes_3_0[0], 3'h0}; // @[FlexDPU.scala 68:35]
  wire [31:0] _FDPE_15_i_mux_bus_3_0_rev_T_4 = {{1'd0}, MuxWrapper_15_Omuxes_3_0[31:1]}; // @[FlexDPU.scala 68:24]
  wire [2:0] _GEN_2742 = {_FDPE_15_i_mux_bus_3_0_rev_T_4[0], 2'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_15_i_mux_bus_3_0_rev_T_6 = {{1'd0}, _GEN_2742}; // @[FlexDPU.scala 68:35]
  wire [3:0] _FDPE_15_i_mux_bus_3_0_rev_T_7 = _FDPE_15_i_mux_bus_3_0_rev_T_2 | _FDPE_15_i_mux_bus_3_0_rev_T_6; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_15_i_mux_bus_3_0_rev_T_8 = {{2'd0}, MuxWrapper_15_Omuxes_3_0[31:2]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_15_i_mux_bus_3_0_rev_T_10 = {_FDPE_15_i_mux_bus_3_0_rev_T_8[0], 1'h0}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2744 = {{2'd0}, _FDPE_15_i_mux_bus_3_0_rev_T_10}; // @[FlexDPU.scala 68:17]
  wire [3:0] _FDPE_15_i_mux_bus_3_0_rev_T_11 = _FDPE_15_i_mux_bus_3_0_rev_T_7 | _GEN_2744; // @[FlexDPU.scala 68:17]
  wire [31:0] _FDPE_15_i_mux_bus_3_0_rev_T_12 = {{3'd0}, MuxWrapper_15_Omuxes_3_0[31:3]}; // @[FlexDPU.scala 68:24]
  wire [1:0] _FDPE_15_i_mux_bus_3_0_rev_T_14 = {{1'd0}, _FDPE_15_i_mux_bus_3_0_rev_T_12[0]}; // @[FlexDPU.scala 68:35]
  wire [3:0] _GEN_2746 = {{2'd0}, _FDPE_15_i_mux_bus_3_0_rev_T_14}; // @[FlexDPU.scala 68:17]
  wire [31:0] _ModuleIndex_T_1 = ModuleIndex + 32'h1; // @[FlexDPU.scala 179:40]
  wire  PF_0_PF_Valid = PathFinder_io_PF_Valid; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] _GEN_268 = 3'h1 == ModuleIndex[2:0] ? io_Streaming_matrix_0_1 : io_Streaming_matrix_0_0; // @[FlexDPU.scala 189:{31,31}]
  wire [15:0] _GEN_269 = 3'h2 == ModuleIndex[2:0] ? io_Streaming_matrix_0_2 : _GEN_268; // @[FlexDPU.scala 189:{31,31}]
  wire [15:0] _GEN_270 = 3'h3 == ModuleIndex[2:0] ? io_Streaming_matrix_0_3 : _GEN_269; // @[FlexDPU.scala 189:{31,31}]
  wire [15:0] _GEN_271 = 3'h4 == ModuleIndex[2:0] ? io_Streaming_matrix_0_4 : _GEN_270; // @[FlexDPU.scala 189:{31,31}]
  wire [15:0] _GEN_272 = 3'h5 == ModuleIndex[2:0] ? io_Streaming_matrix_0_5 : _GEN_271; // @[FlexDPU.scala 189:{31,31}]
  wire [15:0] _GEN_273 = 3'h6 == ModuleIndex[2:0] ? io_Streaming_matrix_0_6 : _GEN_272; // @[FlexDPU.scala 189:{31,31}]
  wire [15:0] _GEN_274 = 3'h7 == ModuleIndex[2:0] ? io_Streaming_matrix_0_7 : _GEN_273; // @[FlexDPU.scala 189:{31,31}]
  wire [15:0] _GEN_276 = 3'h1 == ModuleIndex[2:0] ? io_Streaming_matrix_1_1 : io_Streaming_matrix_1_0; // @[FlexDPU.scala 189:{31,31}]
  wire [15:0] _GEN_277 = 3'h2 == ModuleIndex[2:0] ? io_Streaming_matrix_1_2 : _GEN_276; // @[FlexDPU.scala 189:{31,31}]
  wire [15:0] _GEN_278 = 3'h3 == ModuleIndex[2:0] ? io_Streaming_matrix_1_3 : _GEN_277; // @[FlexDPU.scala 189:{31,31}]
  wire [15:0] _GEN_279 = 3'h4 == ModuleIndex[2:0] ? io_Streaming_matrix_1_4 : _GEN_278; // @[FlexDPU.scala 189:{31,31}]
  wire [15:0] _GEN_280 = 3'h5 == ModuleIndex[2:0] ? io_Streaming_matrix_1_5 : _GEN_279; // @[FlexDPU.scala 189:{31,31}]
  wire [15:0] _GEN_281 = 3'h6 == ModuleIndex[2:0] ? io_Streaming_matrix_1_6 : _GEN_280; // @[FlexDPU.scala 189:{31,31}]
  wire [15:0] _GEN_282 = 3'h7 == ModuleIndex[2:0] ? io_Streaming_matrix_1_7 : _GEN_281; // @[FlexDPU.scala 189:{31,31}]
  wire [15:0] _GEN_284 = 3'h1 == ModuleIndex[2:0] ? io_Streaming_matrix_2_1 : io_Streaming_matrix_2_0; // @[FlexDPU.scala 189:{31,31}]
  wire [15:0] _GEN_285 = 3'h2 == ModuleIndex[2:0] ? io_Streaming_matrix_2_2 : _GEN_284; // @[FlexDPU.scala 189:{31,31}]
  wire [15:0] _GEN_286 = 3'h3 == ModuleIndex[2:0] ? io_Streaming_matrix_2_3 : _GEN_285; // @[FlexDPU.scala 189:{31,31}]
  wire [15:0] _GEN_287 = 3'h4 == ModuleIndex[2:0] ? io_Streaming_matrix_2_4 : _GEN_286; // @[FlexDPU.scala 189:{31,31}]
  wire [15:0] _GEN_288 = 3'h5 == ModuleIndex[2:0] ? io_Streaming_matrix_2_5 : _GEN_287; // @[FlexDPU.scala 189:{31,31}]
  wire [15:0] _GEN_289 = 3'h6 == ModuleIndex[2:0] ? io_Streaming_matrix_2_6 : _GEN_288; // @[FlexDPU.scala 189:{31,31}]
  wire [15:0] _GEN_290 = 3'h7 == ModuleIndex[2:0] ? io_Streaming_matrix_2_7 : _GEN_289; // @[FlexDPU.scala 189:{31,31}]
  wire [15:0] _GEN_292 = 3'h1 == ModuleIndex[2:0] ? io_Streaming_matrix_3_1 : io_Streaming_matrix_3_0; // @[FlexDPU.scala 189:{31,31}]
  wire [15:0] _GEN_293 = 3'h2 == ModuleIndex[2:0] ? io_Streaming_matrix_3_2 : _GEN_292; // @[FlexDPU.scala 189:{31,31}]
  wire [15:0] _GEN_294 = 3'h3 == ModuleIndex[2:0] ? io_Streaming_matrix_3_3 : _GEN_293; // @[FlexDPU.scala 189:{31,31}]
  wire [15:0] _GEN_295 = 3'h4 == ModuleIndex[2:0] ? io_Streaming_matrix_3_4 : _GEN_294; // @[FlexDPU.scala 189:{31,31}]
  wire [15:0] _GEN_296 = 3'h5 == ModuleIndex[2:0] ? io_Streaming_matrix_3_5 : _GEN_295; // @[FlexDPU.scala 189:{31,31}]
  wire [15:0] _GEN_297 = 3'h6 == ModuleIndex[2:0] ? io_Streaming_matrix_3_6 : _GEN_296; // @[FlexDPU.scala 189:{31,31}]
  wire [15:0] _GEN_298 = 3'h7 == ModuleIndex[2:0] ? io_Streaming_matrix_3_7 : _GEN_297; // @[FlexDPU.scala 189:{31,31}]
  wire [15:0] _GEN_300 = 3'h1 == ModuleIndex[2:0] ? io_Streaming_matrix_4_1 : io_Streaming_matrix_4_0; // @[FlexDPU.scala 189:{31,31}]
  wire [15:0] _GEN_301 = 3'h2 == ModuleIndex[2:0] ? io_Streaming_matrix_4_2 : _GEN_300; // @[FlexDPU.scala 189:{31,31}]
  wire [15:0] _GEN_302 = 3'h3 == ModuleIndex[2:0] ? io_Streaming_matrix_4_3 : _GEN_301; // @[FlexDPU.scala 189:{31,31}]
  wire [15:0] _GEN_303 = 3'h4 == ModuleIndex[2:0] ? io_Streaming_matrix_4_4 : _GEN_302; // @[FlexDPU.scala 189:{31,31}]
  wire [15:0] _GEN_304 = 3'h5 == ModuleIndex[2:0] ? io_Streaming_matrix_4_5 : _GEN_303; // @[FlexDPU.scala 189:{31,31}]
  wire [15:0] _GEN_305 = 3'h6 == ModuleIndex[2:0] ? io_Streaming_matrix_4_6 : _GEN_304; // @[FlexDPU.scala 189:{31,31}]
  wire [15:0] _GEN_306 = 3'h7 == ModuleIndex[2:0] ? io_Streaming_matrix_4_7 : _GEN_305; // @[FlexDPU.scala 189:{31,31}]
  wire [15:0] _GEN_308 = 3'h1 == ModuleIndex[2:0] ? io_Streaming_matrix_5_1 : io_Streaming_matrix_5_0; // @[FlexDPU.scala 189:{31,31}]
  wire [15:0] _GEN_309 = 3'h2 == ModuleIndex[2:0] ? io_Streaming_matrix_5_2 : _GEN_308; // @[FlexDPU.scala 189:{31,31}]
  wire [15:0] _GEN_310 = 3'h3 == ModuleIndex[2:0] ? io_Streaming_matrix_5_3 : _GEN_309; // @[FlexDPU.scala 189:{31,31}]
  wire [15:0] _GEN_311 = 3'h4 == ModuleIndex[2:0] ? io_Streaming_matrix_5_4 : _GEN_310; // @[FlexDPU.scala 189:{31,31}]
  wire [15:0] _GEN_312 = 3'h5 == ModuleIndex[2:0] ? io_Streaming_matrix_5_5 : _GEN_311; // @[FlexDPU.scala 189:{31,31}]
  wire [15:0] _GEN_313 = 3'h6 == ModuleIndex[2:0] ? io_Streaming_matrix_5_6 : _GEN_312; // @[FlexDPU.scala 189:{31,31}]
  wire [15:0] _GEN_314 = 3'h7 == ModuleIndex[2:0] ? io_Streaming_matrix_5_7 : _GEN_313; // @[FlexDPU.scala 189:{31,31}]
  wire [15:0] _GEN_316 = 3'h1 == ModuleIndex[2:0] ? io_Streaming_matrix_6_1 : io_Streaming_matrix_6_0; // @[FlexDPU.scala 189:{31,31}]
  wire [15:0] _GEN_317 = 3'h2 == ModuleIndex[2:0] ? io_Streaming_matrix_6_2 : _GEN_316; // @[FlexDPU.scala 189:{31,31}]
  wire [15:0] _GEN_318 = 3'h3 == ModuleIndex[2:0] ? io_Streaming_matrix_6_3 : _GEN_317; // @[FlexDPU.scala 189:{31,31}]
  wire [15:0] _GEN_319 = 3'h4 == ModuleIndex[2:0] ? io_Streaming_matrix_6_4 : _GEN_318; // @[FlexDPU.scala 189:{31,31}]
  wire [15:0] _GEN_320 = 3'h5 == ModuleIndex[2:0] ? io_Streaming_matrix_6_5 : _GEN_319; // @[FlexDPU.scala 189:{31,31}]
  wire [15:0] _GEN_321 = 3'h6 == ModuleIndex[2:0] ? io_Streaming_matrix_6_6 : _GEN_320; // @[FlexDPU.scala 189:{31,31}]
  wire [15:0] _GEN_322 = 3'h7 == ModuleIndex[2:0] ? io_Streaming_matrix_6_7 : _GEN_321; // @[FlexDPU.scala 189:{31,31}]
  wire [15:0] _GEN_324 = 3'h1 == ModuleIndex[2:0] ? io_Streaming_matrix_7_1 : io_Streaming_matrix_7_0; // @[FlexDPU.scala 189:{31,31}]
  wire [15:0] _GEN_325 = 3'h2 == ModuleIndex[2:0] ? io_Streaming_matrix_7_2 : _GEN_324; // @[FlexDPU.scala 189:{31,31}]
  wire [15:0] _GEN_326 = 3'h3 == ModuleIndex[2:0] ? io_Streaming_matrix_7_3 : _GEN_325; // @[FlexDPU.scala 189:{31,31}]
  wire [15:0] _GEN_327 = 3'h4 == ModuleIndex[2:0] ? io_Streaming_matrix_7_4 : _GEN_326; // @[FlexDPU.scala 189:{31,31}]
  wire [15:0] _GEN_328 = 3'h5 == ModuleIndex[2:0] ? io_Streaming_matrix_7_5 : _GEN_327; // @[FlexDPU.scala 189:{31,31}]
  wire [15:0] _GEN_329 = 3'h6 == ModuleIndex[2:0] ? io_Streaming_matrix_7_6 : _GEN_328; // @[FlexDPU.scala 189:{31,31}]
  wire [15:0] _GEN_330 = 3'h7 == ModuleIndex[2:0] ? io_Streaming_matrix_7_7 : _GEN_329; // @[FlexDPU.scala 189:{31,31}]
  wire [31:0] _GEN_397 = Statvalid & check ? PF1_Stream_Col_0 : 32'h0; // @[FlexDPU.scala 112:29 118:32 84:32]
  wire [31:0] _GEN_398 = Statvalid & check ? PF1_Stream_Col_1 : 32'h0; // @[FlexDPU.scala 112:29 118:32 84:32]
  wire [31:0] _GEN_399 = Statvalid & check ? PF1_Stream_Col_2 : 32'h0; // @[FlexDPU.scala 112:29 118:32 84:32]
  wire [31:0] _GEN_400 = Statvalid & check ? PF1_Stream_Col_3 : 32'h0; // @[FlexDPU.scala 112:29 118:32 84:32]
  wire [31:0] _GEN_401 = Statvalid & check ? PF1_Stream_Col_4 : 32'h0; // @[FlexDPU.scala 112:29 118:32 84:32]
  wire [31:0] _GEN_402 = Statvalid & check ? PF1_Stream_Col_5 : 32'h0; // @[FlexDPU.scala 112:29 118:32 84:32]
  wire [31:0] _GEN_403 = Statvalid & check ? PF1_Stream_Col_6 : 32'h0; // @[FlexDPU.scala 112:29 118:32 84:32]
  wire [31:0] _GEN_404 = Statvalid & check ? PF1_Stream_Col_7 : 32'h0; // @[FlexDPU.scala 112:29 118:32 84:32]
  wire [3:0] PF_15_i_mux_bus_0 = PathFinder_15_io_i_mux_bus_0; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_15_i_mux_bus_1 = PathFinder_15_io_i_mux_bus_1; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_15_i_mux_bus_2 = PathFinder_15_io_i_mux_bus_2; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_15_i_mux_bus_3 = PathFinder_15_io_i_mux_bus_3; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_15_Source_0 = PathFinder_15_io_Source_0; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_15_Source_1 = PathFinder_15_io_Source_1; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_15_Source_2 = PathFinder_15_io_Source_2; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_15_Source_3 = PathFinder_15_io_Source_3; // @[FlexDPU.scala 77:{21,21}]
  wire [1:0] _GEN_554 = Statvalid & check ? 2'h2 : 2'h0; // @[FlexDPU.scala 112:29 117:21 83:21]
  wire [1:0] _GEN_627 = Statvalid & check ? 2'h3 : 2'h0; // @[FlexDPU.scala 112:29 117:21 83:21]
  wire [2:0] _GEN_700 = Statvalid & check ? 3'h4 : 3'h0; // @[FlexDPU.scala 112:29 117:21 83:21]
  wire [2:0] _GEN_773 = Statvalid & check ? 3'h5 : 3'h0; // @[FlexDPU.scala 112:29 117:21 83:21]
  wire [2:0] _GEN_846 = Statvalid & check ? 3'h6 : 3'h0; // @[FlexDPU.scala 112:29 117:21 83:21]
  wire [2:0] _GEN_919 = Statvalid & check ? 3'h7 : 3'h0; // @[FlexDPU.scala 112:29 117:21 83:21]
  wire [3:0] _GEN_992 = Statvalid & check ? 4'h8 : 4'h0; // @[FlexDPU.scala 112:29 117:21 83:21]
  wire [3:0] _GEN_1065 = Statvalid & check ? 4'h9 : 4'h0; // @[FlexDPU.scala 112:29 117:21 83:21]
  wire [3:0] _GEN_1138 = Statvalid & check ? 4'ha : 4'h0; // @[FlexDPU.scala 112:29 117:21 83:21]
  wire [3:0] _GEN_1211 = Statvalid & check ? 4'hb : 4'h0; // @[FlexDPU.scala 112:29 117:21 83:21]
  wire [3:0] _GEN_1284 = Statvalid & check ? 4'hc : 4'h0; // @[FlexDPU.scala 112:29 117:21 83:21]
  wire [3:0] _GEN_1357 = Statvalid & check ? 4'hd : 4'h0; // @[FlexDPU.scala 112:29 117:21 83:21]
  wire [3:0] _GEN_1430 = Statvalid & check ? 4'he : 4'h0; // @[FlexDPU.scala 112:29 117:21 83:21]
  wire [3:0] _GEN_1503 = Statvalid & check ? 4'hf : 4'h0; // @[FlexDPU.scala 112:29 117:21 83:21]
  wire [3:0] PF_0_i_mux_bus_0 = PathFinder_io_i_mux_bus_0; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_0_i_mux_bus_1 = PathFinder_io_i_mux_bus_1; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_0_i_mux_bus_2 = PathFinder_io_i_mux_bus_2; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_0_i_mux_bus_3 = PathFinder_io_i_mux_bus_3; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_0_Source_0 = PathFinder_io_Source_0; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_0_Source_1 = PathFinder_io_Source_1; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_0_Source_2 = PathFinder_io_Source_2; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_0_Source_3 = PathFinder_io_Source_3; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_1_i_mux_bus_0 = PathFinder_1_io_i_mux_bus_0; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_1_i_mux_bus_1 = PathFinder_1_io_i_mux_bus_1; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_1_i_mux_bus_2 = PathFinder_1_io_i_mux_bus_2; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_1_i_mux_bus_3 = PathFinder_1_io_i_mux_bus_3; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_1_Source_0 = PathFinder_1_io_Source_0; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_1_Source_1 = PathFinder_1_io_Source_1; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_1_Source_2 = PathFinder_1_io_Source_2; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_1_Source_3 = PathFinder_1_io_Source_3; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_2_i_mux_bus_0 = PathFinder_2_io_i_mux_bus_0; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_2_i_mux_bus_1 = PathFinder_2_io_i_mux_bus_1; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_2_i_mux_bus_2 = PathFinder_2_io_i_mux_bus_2; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_2_i_mux_bus_3 = PathFinder_2_io_i_mux_bus_3; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_2_Source_0 = PathFinder_2_io_Source_0; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_2_Source_1 = PathFinder_2_io_Source_1; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_2_Source_2 = PathFinder_2_io_Source_2; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_2_Source_3 = PathFinder_2_io_Source_3; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_3_i_mux_bus_0 = PathFinder_3_io_i_mux_bus_0; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_3_i_mux_bus_1 = PathFinder_3_io_i_mux_bus_1; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_3_i_mux_bus_2 = PathFinder_3_io_i_mux_bus_2; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_3_i_mux_bus_3 = PathFinder_3_io_i_mux_bus_3; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_3_Source_0 = PathFinder_3_io_Source_0; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_3_Source_1 = PathFinder_3_io_Source_1; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_3_Source_2 = PathFinder_3_io_Source_2; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_3_Source_3 = PathFinder_3_io_Source_3; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_4_i_mux_bus_0 = PathFinder_4_io_i_mux_bus_0; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_4_i_mux_bus_1 = PathFinder_4_io_i_mux_bus_1; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_4_i_mux_bus_2 = PathFinder_4_io_i_mux_bus_2; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_4_i_mux_bus_3 = PathFinder_4_io_i_mux_bus_3; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_4_Source_0 = PathFinder_4_io_Source_0; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_4_Source_1 = PathFinder_4_io_Source_1; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_4_Source_2 = PathFinder_4_io_Source_2; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_4_Source_3 = PathFinder_4_io_Source_3; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_5_i_mux_bus_0 = PathFinder_5_io_i_mux_bus_0; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_5_i_mux_bus_1 = PathFinder_5_io_i_mux_bus_1; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_5_i_mux_bus_2 = PathFinder_5_io_i_mux_bus_2; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_5_i_mux_bus_3 = PathFinder_5_io_i_mux_bus_3; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_5_Source_0 = PathFinder_5_io_Source_0; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_5_Source_1 = PathFinder_5_io_Source_1; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_5_Source_2 = PathFinder_5_io_Source_2; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_5_Source_3 = PathFinder_5_io_Source_3; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_6_i_mux_bus_0 = PathFinder_6_io_i_mux_bus_0; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_6_i_mux_bus_1 = PathFinder_6_io_i_mux_bus_1; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_6_i_mux_bus_2 = PathFinder_6_io_i_mux_bus_2; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_6_i_mux_bus_3 = PathFinder_6_io_i_mux_bus_3; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_6_Source_0 = PathFinder_6_io_Source_0; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_6_Source_1 = PathFinder_6_io_Source_1; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_6_Source_2 = PathFinder_6_io_Source_2; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_6_Source_3 = PathFinder_6_io_Source_3; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_7_i_mux_bus_0 = PathFinder_7_io_i_mux_bus_0; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_7_i_mux_bus_1 = PathFinder_7_io_i_mux_bus_1; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_7_i_mux_bus_2 = PathFinder_7_io_i_mux_bus_2; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_7_i_mux_bus_3 = PathFinder_7_io_i_mux_bus_3; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_7_Source_0 = PathFinder_7_io_Source_0; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_7_Source_1 = PathFinder_7_io_Source_1; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_7_Source_2 = PathFinder_7_io_Source_2; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_7_Source_3 = PathFinder_7_io_Source_3; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_8_i_mux_bus_0 = PathFinder_8_io_i_mux_bus_0; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_8_i_mux_bus_1 = PathFinder_8_io_i_mux_bus_1; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_8_i_mux_bus_2 = PathFinder_8_io_i_mux_bus_2; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_8_i_mux_bus_3 = PathFinder_8_io_i_mux_bus_3; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_8_Source_0 = PathFinder_8_io_Source_0; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_8_Source_1 = PathFinder_8_io_Source_1; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_8_Source_2 = PathFinder_8_io_Source_2; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_8_Source_3 = PathFinder_8_io_Source_3; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_9_i_mux_bus_0 = PathFinder_9_io_i_mux_bus_0; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_9_i_mux_bus_1 = PathFinder_9_io_i_mux_bus_1; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_9_i_mux_bus_2 = PathFinder_9_io_i_mux_bus_2; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_9_i_mux_bus_3 = PathFinder_9_io_i_mux_bus_3; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_9_Source_0 = PathFinder_9_io_Source_0; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_9_Source_1 = PathFinder_9_io_Source_1; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_9_Source_2 = PathFinder_9_io_Source_2; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_9_Source_3 = PathFinder_9_io_Source_3; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_10_i_mux_bus_0 = PathFinder_10_io_i_mux_bus_0; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_10_i_mux_bus_1 = PathFinder_10_io_i_mux_bus_1; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_10_i_mux_bus_2 = PathFinder_10_io_i_mux_bus_2; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_10_i_mux_bus_3 = PathFinder_10_io_i_mux_bus_3; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_10_Source_0 = PathFinder_10_io_Source_0; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_10_Source_1 = PathFinder_10_io_Source_1; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_10_Source_2 = PathFinder_10_io_Source_2; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_10_Source_3 = PathFinder_10_io_Source_3; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_11_i_mux_bus_0 = PathFinder_11_io_i_mux_bus_0; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_11_i_mux_bus_1 = PathFinder_11_io_i_mux_bus_1; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_11_i_mux_bus_2 = PathFinder_11_io_i_mux_bus_2; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_11_i_mux_bus_3 = PathFinder_11_io_i_mux_bus_3; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_11_Source_0 = PathFinder_11_io_Source_0; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_11_Source_1 = PathFinder_11_io_Source_1; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_11_Source_2 = PathFinder_11_io_Source_2; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_11_Source_3 = PathFinder_11_io_Source_3; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_12_i_mux_bus_0 = PathFinder_12_io_i_mux_bus_0; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_12_i_mux_bus_1 = PathFinder_12_io_i_mux_bus_1; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_12_i_mux_bus_2 = PathFinder_12_io_i_mux_bus_2; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_12_i_mux_bus_3 = PathFinder_12_io_i_mux_bus_3; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_12_Source_0 = PathFinder_12_io_Source_0; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_12_Source_1 = PathFinder_12_io_Source_1; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_12_Source_2 = PathFinder_12_io_Source_2; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_12_Source_3 = PathFinder_12_io_Source_3; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_13_i_mux_bus_0 = PathFinder_13_io_i_mux_bus_0; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_13_i_mux_bus_1 = PathFinder_13_io_i_mux_bus_1; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_13_i_mux_bus_2 = PathFinder_13_io_i_mux_bus_2; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_13_i_mux_bus_3 = PathFinder_13_io_i_mux_bus_3; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_13_Source_0 = PathFinder_13_io_Source_0; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_13_Source_1 = PathFinder_13_io_Source_1; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_13_Source_2 = PathFinder_13_io_Source_2; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_13_Source_3 = PathFinder_13_io_Source_3; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_14_i_mux_bus_0 = PathFinder_14_io_i_mux_bus_0; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_14_i_mux_bus_1 = PathFinder_14_io_i_mux_bus_1; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_14_i_mux_bus_2 = PathFinder_14_io_i_mux_bus_2; // @[FlexDPU.scala 77:{21,21}]
  wire [3:0] PF_14_i_mux_bus_3 = PathFinder_14_io_i_mux_bus_3; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_14_Source_0 = PathFinder_14_io_Source_0; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_14_Source_1 = PathFinder_14_io_Source_1; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_14_Source_2 = PathFinder_14_io_Source_2; // @[FlexDPU.scala 77:{21,21}]
  wire [15:0] PF_14_Source_3 = PathFinder_14_io_Source_3; // @[FlexDPU.scala 77:{21,21}]
  wire [31:0] MuxWrapper_0_Osrc_0 = MuxesWrapper_io_Osrc_0; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_0_Osrc_1 = MuxesWrapper_io_Osrc_1; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_0_Osrc_2 = MuxesWrapper_io_Osrc_2; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_0_Osrc_3 = MuxesWrapper_io_Osrc_3; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_1_Osrc_0 = MuxesWrapper_1_io_Osrc_0; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_1_Osrc_1 = MuxesWrapper_1_io_Osrc_1; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_1_Osrc_2 = MuxesWrapper_1_io_Osrc_2; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_1_Osrc_3 = MuxesWrapper_1_io_Osrc_3; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_2_Osrc_0 = MuxesWrapper_2_io_Osrc_0; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_2_Osrc_1 = MuxesWrapper_2_io_Osrc_1; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_2_Osrc_2 = MuxesWrapper_2_io_Osrc_2; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_2_Osrc_3 = MuxesWrapper_2_io_Osrc_3; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_3_Osrc_0 = MuxesWrapper_3_io_Osrc_0; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_3_Osrc_1 = MuxesWrapper_3_io_Osrc_1; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_3_Osrc_2 = MuxesWrapper_3_io_Osrc_2; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_3_Osrc_3 = MuxesWrapper_3_io_Osrc_3; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_4_Osrc_0 = MuxesWrapper_4_io_Osrc_0; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_4_Osrc_1 = MuxesWrapper_4_io_Osrc_1; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_4_Osrc_2 = MuxesWrapper_4_io_Osrc_2; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_4_Osrc_3 = MuxesWrapper_4_io_Osrc_3; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_5_Osrc_0 = MuxesWrapper_5_io_Osrc_0; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_5_Osrc_1 = MuxesWrapper_5_io_Osrc_1; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_5_Osrc_2 = MuxesWrapper_5_io_Osrc_2; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_5_Osrc_3 = MuxesWrapper_5_io_Osrc_3; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_6_Osrc_0 = MuxesWrapper_6_io_Osrc_0; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_6_Osrc_1 = MuxesWrapper_6_io_Osrc_1; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_6_Osrc_2 = MuxesWrapper_6_io_Osrc_2; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_6_Osrc_3 = MuxesWrapper_6_io_Osrc_3; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_7_Osrc_0 = MuxesWrapper_7_io_Osrc_0; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_7_Osrc_1 = MuxesWrapper_7_io_Osrc_1; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_7_Osrc_2 = MuxesWrapper_7_io_Osrc_2; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_7_Osrc_3 = MuxesWrapper_7_io_Osrc_3; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_8_Osrc_0 = MuxesWrapper_8_io_Osrc_0; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_8_Osrc_1 = MuxesWrapper_8_io_Osrc_1; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_8_Osrc_2 = MuxesWrapper_8_io_Osrc_2; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_8_Osrc_3 = MuxesWrapper_8_io_Osrc_3; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_9_Osrc_0 = MuxesWrapper_9_io_Osrc_0; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_9_Osrc_1 = MuxesWrapper_9_io_Osrc_1; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_9_Osrc_2 = MuxesWrapper_9_io_Osrc_2; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_9_Osrc_3 = MuxesWrapper_9_io_Osrc_3; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_10_Osrc_0 = MuxesWrapper_10_io_Osrc_0; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_10_Osrc_1 = MuxesWrapper_10_io_Osrc_1; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_10_Osrc_2 = MuxesWrapper_10_io_Osrc_2; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_10_Osrc_3 = MuxesWrapper_10_io_Osrc_3; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_11_Osrc_0 = MuxesWrapper_11_io_Osrc_0; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_11_Osrc_1 = MuxesWrapper_11_io_Osrc_1; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_11_Osrc_2 = MuxesWrapper_11_io_Osrc_2; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_11_Osrc_3 = MuxesWrapper_11_io_Osrc_3; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_12_Osrc_0 = MuxesWrapper_12_io_Osrc_0; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_12_Osrc_1 = MuxesWrapper_12_io_Osrc_1; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_12_Osrc_2 = MuxesWrapper_12_io_Osrc_2; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_12_Osrc_3 = MuxesWrapper_12_io_Osrc_3; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_13_Osrc_0 = MuxesWrapper_13_io_Osrc_0; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_13_Osrc_1 = MuxesWrapper_13_io_Osrc_1; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_13_Osrc_2 = MuxesWrapper_13_io_Osrc_2; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_13_Osrc_3 = MuxesWrapper_13_io_Osrc_3; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_14_Osrc_0 = MuxesWrapper_14_io_Osrc_0; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_14_Osrc_1 = MuxesWrapper_14_io_Osrc_1; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_14_Osrc_2 = MuxesWrapper_14_io_Osrc_2; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_14_Osrc_3 = MuxesWrapper_14_io_Osrc_3; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_15_Osrc_0 = MuxesWrapper_15_io_Osrc_0; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_15_Osrc_1 = MuxesWrapper_15_io_Osrc_1; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_15_Osrc_2 = MuxesWrapper_15_io_Osrc_2; // @[FlexDPU.scala 124:{33,33}]
  wire [31:0] MuxWrapper_15_Osrc_3 = MuxesWrapper_15_io_Osrc_3; // @[FlexDPU.scala 124:{33,33}]
  wire [15:0] FDPE_0_o_adder_0 = flexdpecom4_io_o_adder_0; // @[FlexDPU.scala 132:{27,27}]
  wire [15:0] FDPE_0_o_adder_1 = flexdpecom4_io_o_adder_1; // @[FlexDPU.scala 132:{27,27}]
  wire [15:0] FDPE_0_o_adder_2 = flexdpecom4_io_o_adder_2; // @[FlexDPU.scala 132:{27,27}]
  wire [15:0] FDPE_1_o_adder_0 = flexdpecom4_1_io_o_adder_0; // @[FlexDPU.scala 132:{27,27}]
  wire [15:0] FDPE_1_o_adder_1 = flexdpecom4_1_io_o_adder_1; // @[FlexDPU.scala 132:{27,27}]
  wire [15:0] FDPE_1_o_adder_2 = flexdpecom4_1_io_o_adder_2; // @[FlexDPU.scala 132:{27,27}]
  wire [15:0] FDPE_2_o_adder_0 = flexdpecom4_2_io_o_adder_0; // @[FlexDPU.scala 132:{27,27}]
  wire [15:0] FDPE_2_o_adder_1 = flexdpecom4_2_io_o_adder_1; // @[FlexDPU.scala 132:{27,27}]
  wire [15:0] FDPE_2_o_adder_2 = flexdpecom4_2_io_o_adder_2; // @[FlexDPU.scala 132:{27,27}]
  wire [15:0] FDPE_3_o_adder_0 = flexdpecom4_3_io_o_adder_0; // @[FlexDPU.scala 132:{27,27}]
  wire [15:0] FDPE_3_o_adder_1 = flexdpecom4_3_io_o_adder_1; // @[FlexDPU.scala 132:{27,27}]
  wire [15:0] FDPE_3_o_adder_2 = flexdpecom4_3_io_o_adder_2; // @[FlexDPU.scala 132:{27,27}]
  wire [15:0] FDPE_4_o_adder_0 = flexdpecom4_4_io_o_adder_0; // @[FlexDPU.scala 132:{27,27}]
  wire [15:0] FDPE_4_o_adder_1 = flexdpecom4_4_io_o_adder_1; // @[FlexDPU.scala 132:{27,27}]
  wire [15:0] FDPE_4_o_adder_2 = flexdpecom4_4_io_o_adder_2; // @[FlexDPU.scala 132:{27,27}]
  wire [15:0] FDPE_5_o_adder_0 = flexdpecom4_5_io_o_adder_0; // @[FlexDPU.scala 132:{27,27}]
  wire [15:0] FDPE_5_o_adder_1 = flexdpecom4_5_io_o_adder_1; // @[FlexDPU.scala 132:{27,27}]
  wire [15:0] FDPE_5_o_adder_2 = flexdpecom4_5_io_o_adder_2; // @[FlexDPU.scala 132:{27,27}]
  wire [15:0] FDPE_6_o_adder_0 = flexdpecom4_6_io_o_adder_0; // @[FlexDPU.scala 132:{27,27}]
  wire [15:0] FDPE_6_o_adder_1 = flexdpecom4_6_io_o_adder_1; // @[FlexDPU.scala 132:{27,27}]
  wire [15:0] FDPE_6_o_adder_2 = flexdpecom4_6_io_o_adder_2; // @[FlexDPU.scala 132:{27,27}]
  wire [15:0] FDPE_7_o_adder_0 = flexdpecom4_7_io_o_adder_0; // @[FlexDPU.scala 132:{27,27}]
  wire [15:0] FDPE_7_o_adder_1 = flexdpecom4_7_io_o_adder_1; // @[FlexDPU.scala 132:{27,27}]
  wire [15:0] FDPE_7_o_adder_2 = flexdpecom4_7_io_o_adder_2; // @[FlexDPU.scala 132:{27,27}]
  wire [15:0] FDPE_8_o_adder_0 = flexdpecom4_8_io_o_adder_0; // @[FlexDPU.scala 132:{27,27}]
  wire [15:0] FDPE_8_o_adder_1 = flexdpecom4_8_io_o_adder_1; // @[FlexDPU.scala 132:{27,27}]
  wire [15:0] FDPE_8_o_adder_2 = flexdpecom4_8_io_o_adder_2; // @[FlexDPU.scala 132:{27,27}]
  wire [15:0] FDPE_9_o_adder_0 = flexdpecom4_9_io_o_adder_0; // @[FlexDPU.scala 132:{27,27}]
  wire [15:0] FDPE_9_o_adder_1 = flexdpecom4_9_io_o_adder_1; // @[FlexDPU.scala 132:{27,27}]
  wire [15:0] FDPE_9_o_adder_2 = flexdpecom4_9_io_o_adder_2; // @[FlexDPU.scala 132:{27,27}]
  wire [15:0] FDPE_10_o_adder_0 = flexdpecom4_10_io_o_adder_0; // @[FlexDPU.scala 132:{27,27}]
  wire [15:0] FDPE_10_o_adder_1 = flexdpecom4_10_io_o_adder_1; // @[FlexDPU.scala 132:{27,27}]
  wire [15:0] FDPE_10_o_adder_2 = flexdpecom4_10_io_o_adder_2; // @[FlexDPU.scala 132:{27,27}]
  wire [15:0] FDPE_11_o_adder_0 = flexdpecom4_11_io_o_adder_0; // @[FlexDPU.scala 132:{27,27}]
  wire [15:0] FDPE_11_o_adder_1 = flexdpecom4_11_io_o_adder_1; // @[FlexDPU.scala 132:{27,27}]
  wire [15:0] FDPE_11_o_adder_2 = flexdpecom4_11_io_o_adder_2; // @[FlexDPU.scala 132:{27,27}]
  wire [15:0] FDPE_12_o_adder_0 = flexdpecom4_12_io_o_adder_0; // @[FlexDPU.scala 132:{27,27}]
  wire [15:0] FDPE_12_o_adder_1 = flexdpecom4_12_io_o_adder_1; // @[FlexDPU.scala 132:{27,27}]
  wire [15:0] FDPE_12_o_adder_2 = flexdpecom4_12_io_o_adder_2; // @[FlexDPU.scala 132:{27,27}]
  wire [15:0] FDPE_13_o_adder_0 = flexdpecom4_13_io_o_adder_0; // @[FlexDPU.scala 132:{27,27}]
  wire [15:0] FDPE_13_o_adder_1 = flexdpecom4_13_io_o_adder_1; // @[FlexDPU.scala 132:{27,27}]
  wire [15:0] FDPE_13_o_adder_2 = flexdpecom4_13_io_o_adder_2; // @[FlexDPU.scala 132:{27,27}]
  wire [15:0] FDPE_14_o_adder_0 = flexdpecom4_14_io_o_adder_0; // @[FlexDPU.scala 132:{27,27}]
  wire [15:0] FDPE_14_o_adder_1 = flexdpecom4_14_io_o_adder_1; // @[FlexDPU.scala 132:{27,27}]
  wire [15:0] FDPE_14_o_adder_2 = flexdpecom4_14_io_o_adder_2; // @[FlexDPU.scala 132:{27,27}]
  wire [15:0] FDPE_15_o_adder_0 = flexdpecom4_15_io_o_adder_0; // @[FlexDPU.scala 132:{27,27}]
  wire [15:0] FDPE_15_o_adder_1 = flexdpecom4_15_io_o_adder_1; // @[FlexDPU.scala 132:{27,27}]
  wire [15:0] FDPE_15_o_adder_2 = flexdpecom4_15_io_o_adder_2; // @[FlexDPU.scala 132:{27,27}]
  PathFinder PathFinder ( // @[FlexDPU.scala 77:41]
    .clock(PathFinder_clock),
    .reset(PathFinder_reset),
    .io_Stationary_matrix_0_0(PathFinder_io_Stationary_matrix_0_0),
    .io_Stationary_matrix_0_1(PathFinder_io_Stationary_matrix_0_1),
    .io_Stationary_matrix_0_2(PathFinder_io_Stationary_matrix_0_2),
    .io_Stationary_matrix_0_3(PathFinder_io_Stationary_matrix_0_3),
    .io_Stationary_matrix_0_4(PathFinder_io_Stationary_matrix_0_4),
    .io_Stationary_matrix_0_5(PathFinder_io_Stationary_matrix_0_5),
    .io_Stationary_matrix_0_6(PathFinder_io_Stationary_matrix_0_6),
    .io_Stationary_matrix_0_7(PathFinder_io_Stationary_matrix_0_7),
    .io_Stationary_matrix_1_0(PathFinder_io_Stationary_matrix_1_0),
    .io_Stationary_matrix_1_1(PathFinder_io_Stationary_matrix_1_1),
    .io_Stationary_matrix_1_2(PathFinder_io_Stationary_matrix_1_2),
    .io_Stationary_matrix_1_3(PathFinder_io_Stationary_matrix_1_3),
    .io_Stationary_matrix_1_4(PathFinder_io_Stationary_matrix_1_4),
    .io_Stationary_matrix_1_5(PathFinder_io_Stationary_matrix_1_5),
    .io_Stationary_matrix_1_6(PathFinder_io_Stationary_matrix_1_6),
    .io_Stationary_matrix_1_7(PathFinder_io_Stationary_matrix_1_7),
    .io_Stationary_matrix_2_0(PathFinder_io_Stationary_matrix_2_0),
    .io_Stationary_matrix_2_1(PathFinder_io_Stationary_matrix_2_1),
    .io_Stationary_matrix_2_2(PathFinder_io_Stationary_matrix_2_2),
    .io_Stationary_matrix_2_3(PathFinder_io_Stationary_matrix_2_3),
    .io_Stationary_matrix_2_4(PathFinder_io_Stationary_matrix_2_4),
    .io_Stationary_matrix_2_5(PathFinder_io_Stationary_matrix_2_5),
    .io_Stationary_matrix_2_6(PathFinder_io_Stationary_matrix_2_6),
    .io_Stationary_matrix_2_7(PathFinder_io_Stationary_matrix_2_7),
    .io_Stationary_matrix_3_0(PathFinder_io_Stationary_matrix_3_0),
    .io_Stationary_matrix_3_1(PathFinder_io_Stationary_matrix_3_1),
    .io_Stationary_matrix_3_2(PathFinder_io_Stationary_matrix_3_2),
    .io_Stationary_matrix_3_3(PathFinder_io_Stationary_matrix_3_3),
    .io_Stationary_matrix_3_4(PathFinder_io_Stationary_matrix_3_4),
    .io_Stationary_matrix_3_5(PathFinder_io_Stationary_matrix_3_5),
    .io_Stationary_matrix_3_6(PathFinder_io_Stationary_matrix_3_6),
    .io_Stationary_matrix_3_7(PathFinder_io_Stationary_matrix_3_7),
    .io_Stationary_matrix_4_0(PathFinder_io_Stationary_matrix_4_0),
    .io_Stationary_matrix_4_1(PathFinder_io_Stationary_matrix_4_1),
    .io_Stationary_matrix_4_2(PathFinder_io_Stationary_matrix_4_2),
    .io_Stationary_matrix_4_3(PathFinder_io_Stationary_matrix_4_3),
    .io_Stationary_matrix_4_4(PathFinder_io_Stationary_matrix_4_4),
    .io_Stationary_matrix_4_5(PathFinder_io_Stationary_matrix_4_5),
    .io_Stationary_matrix_4_6(PathFinder_io_Stationary_matrix_4_6),
    .io_Stationary_matrix_4_7(PathFinder_io_Stationary_matrix_4_7),
    .io_Stationary_matrix_5_0(PathFinder_io_Stationary_matrix_5_0),
    .io_Stationary_matrix_5_1(PathFinder_io_Stationary_matrix_5_1),
    .io_Stationary_matrix_5_2(PathFinder_io_Stationary_matrix_5_2),
    .io_Stationary_matrix_5_3(PathFinder_io_Stationary_matrix_5_3),
    .io_Stationary_matrix_5_4(PathFinder_io_Stationary_matrix_5_4),
    .io_Stationary_matrix_5_5(PathFinder_io_Stationary_matrix_5_5),
    .io_Stationary_matrix_5_6(PathFinder_io_Stationary_matrix_5_6),
    .io_Stationary_matrix_5_7(PathFinder_io_Stationary_matrix_5_7),
    .io_Stationary_matrix_6_0(PathFinder_io_Stationary_matrix_6_0),
    .io_Stationary_matrix_6_1(PathFinder_io_Stationary_matrix_6_1),
    .io_Stationary_matrix_6_2(PathFinder_io_Stationary_matrix_6_2),
    .io_Stationary_matrix_6_3(PathFinder_io_Stationary_matrix_6_3),
    .io_Stationary_matrix_6_4(PathFinder_io_Stationary_matrix_6_4),
    .io_Stationary_matrix_6_5(PathFinder_io_Stationary_matrix_6_5),
    .io_Stationary_matrix_6_6(PathFinder_io_Stationary_matrix_6_6),
    .io_Stationary_matrix_6_7(PathFinder_io_Stationary_matrix_6_7),
    .io_Stationary_matrix_7_0(PathFinder_io_Stationary_matrix_7_0),
    .io_Stationary_matrix_7_1(PathFinder_io_Stationary_matrix_7_1),
    .io_Stationary_matrix_7_2(PathFinder_io_Stationary_matrix_7_2),
    .io_Stationary_matrix_7_3(PathFinder_io_Stationary_matrix_7_3),
    .io_Stationary_matrix_7_4(PathFinder_io_Stationary_matrix_7_4),
    .io_Stationary_matrix_7_5(PathFinder_io_Stationary_matrix_7_5),
    .io_Stationary_matrix_7_6(PathFinder_io_Stationary_matrix_7_6),
    .io_Stationary_matrix_7_7(PathFinder_io_Stationary_matrix_7_7),
    .io_Streaming_matrix_0(PathFinder_io_Streaming_matrix_0),
    .io_Streaming_matrix_1(PathFinder_io_Streaming_matrix_1),
    .io_Streaming_matrix_2(PathFinder_io_Streaming_matrix_2),
    .io_Streaming_matrix_3(PathFinder_io_Streaming_matrix_3),
    .io_Streaming_matrix_4(PathFinder_io_Streaming_matrix_4),
    .io_Streaming_matrix_5(PathFinder_io_Streaming_matrix_5),
    .io_Streaming_matrix_6(PathFinder_io_Streaming_matrix_6),
    .io_Streaming_matrix_7(PathFinder_io_Streaming_matrix_7),
    .io_i_mux_bus_0(PathFinder_io_i_mux_bus_0),
    .io_i_mux_bus_1(PathFinder_io_i_mux_bus_1),
    .io_i_mux_bus_2(PathFinder_io_i_mux_bus_2),
    .io_i_mux_bus_3(PathFinder_io_i_mux_bus_3),
    .io_Source_0(PathFinder_io_Source_0),
    .io_Source_1(PathFinder_io_Source_1),
    .io_Source_2(PathFinder_io_Source_2),
    .io_Source_3(PathFinder_io_Source_3),
    .io_PF_Valid(PathFinder_io_PF_Valid),
    .io_NoDPE(PathFinder_io_NoDPE),
    .io_DataValid(PathFinder_io_DataValid)
  );
  PathFinder PathFinder_1 ( // @[FlexDPU.scala 77:41]
    .clock(PathFinder_1_clock),
    .reset(PathFinder_1_reset),
    .io_Stationary_matrix_0_0(PathFinder_1_io_Stationary_matrix_0_0),
    .io_Stationary_matrix_0_1(PathFinder_1_io_Stationary_matrix_0_1),
    .io_Stationary_matrix_0_2(PathFinder_1_io_Stationary_matrix_0_2),
    .io_Stationary_matrix_0_3(PathFinder_1_io_Stationary_matrix_0_3),
    .io_Stationary_matrix_0_4(PathFinder_1_io_Stationary_matrix_0_4),
    .io_Stationary_matrix_0_5(PathFinder_1_io_Stationary_matrix_0_5),
    .io_Stationary_matrix_0_6(PathFinder_1_io_Stationary_matrix_0_6),
    .io_Stationary_matrix_0_7(PathFinder_1_io_Stationary_matrix_0_7),
    .io_Stationary_matrix_1_0(PathFinder_1_io_Stationary_matrix_1_0),
    .io_Stationary_matrix_1_1(PathFinder_1_io_Stationary_matrix_1_1),
    .io_Stationary_matrix_1_2(PathFinder_1_io_Stationary_matrix_1_2),
    .io_Stationary_matrix_1_3(PathFinder_1_io_Stationary_matrix_1_3),
    .io_Stationary_matrix_1_4(PathFinder_1_io_Stationary_matrix_1_4),
    .io_Stationary_matrix_1_5(PathFinder_1_io_Stationary_matrix_1_5),
    .io_Stationary_matrix_1_6(PathFinder_1_io_Stationary_matrix_1_6),
    .io_Stationary_matrix_1_7(PathFinder_1_io_Stationary_matrix_1_7),
    .io_Stationary_matrix_2_0(PathFinder_1_io_Stationary_matrix_2_0),
    .io_Stationary_matrix_2_1(PathFinder_1_io_Stationary_matrix_2_1),
    .io_Stationary_matrix_2_2(PathFinder_1_io_Stationary_matrix_2_2),
    .io_Stationary_matrix_2_3(PathFinder_1_io_Stationary_matrix_2_3),
    .io_Stationary_matrix_2_4(PathFinder_1_io_Stationary_matrix_2_4),
    .io_Stationary_matrix_2_5(PathFinder_1_io_Stationary_matrix_2_5),
    .io_Stationary_matrix_2_6(PathFinder_1_io_Stationary_matrix_2_6),
    .io_Stationary_matrix_2_7(PathFinder_1_io_Stationary_matrix_2_7),
    .io_Stationary_matrix_3_0(PathFinder_1_io_Stationary_matrix_3_0),
    .io_Stationary_matrix_3_1(PathFinder_1_io_Stationary_matrix_3_1),
    .io_Stationary_matrix_3_2(PathFinder_1_io_Stationary_matrix_3_2),
    .io_Stationary_matrix_3_3(PathFinder_1_io_Stationary_matrix_3_3),
    .io_Stationary_matrix_3_4(PathFinder_1_io_Stationary_matrix_3_4),
    .io_Stationary_matrix_3_5(PathFinder_1_io_Stationary_matrix_3_5),
    .io_Stationary_matrix_3_6(PathFinder_1_io_Stationary_matrix_3_6),
    .io_Stationary_matrix_3_7(PathFinder_1_io_Stationary_matrix_3_7),
    .io_Stationary_matrix_4_0(PathFinder_1_io_Stationary_matrix_4_0),
    .io_Stationary_matrix_4_1(PathFinder_1_io_Stationary_matrix_4_1),
    .io_Stationary_matrix_4_2(PathFinder_1_io_Stationary_matrix_4_2),
    .io_Stationary_matrix_4_3(PathFinder_1_io_Stationary_matrix_4_3),
    .io_Stationary_matrix_4_4(PathFinder_1_io_Stationary_matrix_4_4),
    .io_Stationary_matrix_4_5(PathFinder_1_io_Stationary_matrix_4_5),
    .io_Stationary_matrix_4_6(PathFinder_1_io_Stationary_matrix_4_6),
    .io_Stationary_matrix_4_7(PathFinder_1_io_Stationary_matrix_4_7),
    .io_Stationary_matrix_5_0(PathFinder_1_io_Stationary_matrix_5_0),
    .io_Stationary_matrix_5_1(PathFinder_1_io_Stationary_matrix_5_1),
    .io_Stationary_matrix_5_2(PathFinder_1_io_Stationary_matrix_5_2),
    .io_Stationary_matrix_5_3(PathFinder_1_io_Stationary_matrix_5_3),
    .io_Stationary_matrix_5_4(PathFinder_1_io_Stationary_matrix_5_4),
    .io_Stationary_matrix_5_5(PathFinder_1_io_Stationary_matrix_5_5),
    .io_Stationary_matrix_5_6(PathFinder_1_io_Stationary_matrix_5_6),
    .io_Stationary_matrix_5_7(PathFinder_1_io_Stationary_matrix_5_7),
    .io_Stationary_matrix_6_0(PathFinder_1_io_Stationary_matrix_6_0),
    .io_Stationary_matrix_6_1(PathFinder_1_io_Stationary_matrix_6_1),
    .io_Stationary_matrix_6_2(PathFinder_1_io_Stationary_matrix_6_2),
    .io_Stationary_matrix_6_3(PathFinder_1_io_Stationary_matrix_6_3),
    .io_Stationary_matrix_6_4(PathFinder_1_io_Stationary_matrix_6_4),
    .io_Stationary_matrix_6_5(PathFinder_1_io_Stationary_matrix_6_5),
    .io_Stationary_matrix_6_6(PathFinder_1_io_Stationary_matrix_6_6),
    .io_Stationary_matrix_6_7(PathFinder_1_io_Stationary_matrix_6_7),
    .io_Stationary_matrix_7_0(PathFinder_1_io_Stationary_matrix_7_0),
    .io_Stationary_matrix_7_1(PathFinder_1_io_Stationary_matrix_7_1),
    .io_Stationary_matrix_7_2(PathFinder_1_io_Stationary_matrix_7_2),
    .io_Stationary_matrix_7_3(PathFinder_1_io_Stationary_matrix_7_3),
    .io_Stationary_matrix_7_4(PathFinder_1_io_Stationary_matrix_7_4),
    .io_Stationary_matrix_7_5(PathFinder_1_io_Stationary_matrix_7_5),
    .io_Stationary_matrix_7_6(PathFinder_1_io_Stationary_matrix_7_6),
    .io_Stationary_matrix_7_7(PathFinder_1_io_Stationary_matrix_7_7),
    .io_Streaming_matrix_0(PathFinder_1_io_Streaming_matrix_0),
    .io_Streaming_matrix_1(PathFinder_1_io_Streaming_matrix_1),
    .io_Streaming_matrix_2(PathFinder_1_io_Streaming_matrix_2),
    .io_Streaming_matrix_3(PathFinder_1_io_Streaming_matrix_3),
    .io_Streaming_matrix_4(PathFinder_1_io_Streaming_matrix_4),
    .io_Streaming_matrix_5(PathFinder_1_io_Streaming_matrix_5),
    .io_Streaming_matrix_6(PathFinder_1_io_Streaming_matrix_6),
    .io_Streaming_matrix_7(PathFinder_1_io_Streaming_matrix_7),
    .io_i_mux_bus_0(PathFinder_1_io_i_mux_bus_0),
    .io_i_mux_bus_1(PathFinder_1_io_i_mux_bus_1),
    .io_i_mux_bus_2(PathFinder_1_io_i_mux_bus_2),
    .io_i_mux_bus_3(PathFinder_1_io_i_mux_bus_3),
    .io_Source_0(PathFinder_1_io_Source_0),
    .io_Source_1(PathFinder_1_io_Source_1),
    .io_Source_2(PathFinder_1_io_Source_2),
    .io_Source_3(PathFinder_1_io_Source_3),
    .io_PF_Valid(PathFinder_1_io_PF_Valid),
    .io_NoDPE(PathFinder_1_io_NoDPE),
    .io_DataValid(PathFinder_1_io_DataValid)
  );
  PathFinder PathFinder_2 ( // @[FlexDPU.scala 77:41]
    .clock(PathFinder_2_clock),
    .reset(PathFinder_2_reset),
    .io_Stationary_matrix_0_0(PathFinder_2_io_Stationary_matrix_0_0),
    .io_Stationary_matrix_0_1(PathFinder_2_io_Stationary_matrix_0_1),
    .io_Stationary_matrix_0_2(PathFinder_2_io_Stationary_matrix_0_2),
    .io_Stationary_matrix_0_3(PathFinder_2_io_Stationary_matrix_0_3),
    .io_Stationary_matrix_0_4(PathFinder_2_io_Stationary_matrix_0_4),
    .io_Stationary_matrix_0_5(PathFinder_2_io_Stationary_matrix_0_5),
    .io_Stationary_matrix_0_6(PathFinder_2_io_Stationary_matrix_0_6),
    .io_Stationary_matrix_0_7(PathFinder_2_io_Stationary_matrix_0_7),
    .io_Stationary_matrix_1_0(PathFinder_2_io_Stationary_matrix_1_0),
    .io_Stationary_matrix_1_1(PathFinder_2_io_Stationary_matrix_1_1),
    .io_Stationary_matrix_1_2(PathFinder_2_io_Stationary_matrix_1_2),
    .io_Stationary_matrix_1_3(PathFinder_2_io_Stationary_matrix_1_3),
    .io_Stationary_matrix_1_4(PathFinder_2_io_Stationary_matrix_1_4),
    .io_Stationary_matrix_1_5(PathFinder_2_io_Stationary_matrix_1_5),
    .io_Stationary_matrix_1_6(PathFinder_2_io_Stationary_matrix_1_6),
    .io_Stationary_matrix_1_7(PathFinder_2_io_Stationary_matrix_1_7),
    .io_Stationary_matrix_2_0(PathFinder_2_io_Stationary_matrix_2_0),
    .io_Stationary_matrix_2_1(PathFinder_2_io_Stationary_matrix_2_1),
    .io_Stationary_matrix_2_2(PathFinder_2_io_Stationary_matrix_2_2),
    .io_Stationary_matrix_2_3(PathFinder_2_io_Stationary_matrix_2_3),
    .io_Stationary_matrix_2_4(PathFinder_2_io_Stationary_matrix_2_4),
    .io_Stationary_matrix_2_5(PathFinder_2_io_Stationary_matrix_2_5),
    .io_Stationary_matrix_2_6(PathFinder_2_io_Stationary_matrix_2_6),
    .io_Stationary_matrix_2_7(PathFinder_2_io_Stationary_matrix_2_7),
    .io_Stationary_matrix_3_0(PathFinder_2_io_Stationary_matrix_3_0),
    .io_Stationary_matrix_3_1(PathFinder_2_io_Stationary_matrix_3_1),
    .io_Stationary_matrix_3_2(PathFinder_2_io_Stationary_matrix_3_2),
    .io_Stationary_matrix_3_3(PathFinder_2_io_Stationary_matrix_3_3),
    .io_Stationary_matrix_3_4(PathFinder_2_io_Stationary_matrix_3_4),
    .io_Stationary_matrix_3_5(PathFinder_2_io_Stationary_matrix_3_5),
    .io_Stationary_matrix_3_6(PathFinder_2_io_Stationary_matrix_3_6),
    .io_Stationary_matrix_3_7(PathFinder_2_io_Stationary_matrix_3_7),
    .io_Stationary_matrix_4_0(PathFinder_2_io_Stationary_matrix_4_0),
    .io_Stationary_matrix_4_1(PathFinder_2_io_Stationary_matrix_4_1),
    .io_Stationary_matrix_4_2(PathFinder_2_io_Stationary_matrix_4_2),
    .io_Stationary_matrix_4_3(PathFinder_2_io_Stationary_matrix_4_3),
    .io_Stationary_matrix_4_4(PathFinder_2_io_Stationary_matrix_4_4),
    .io_Stationary_matrix_4_5(PathFinder_2_io_Stationary_matrix_4_5),
    .io_Stationary_matrix_4_6(PathFinder_2_io_Stationary_matrix_4_6),
    .io_Stationary_matrix_4_7(PathFinder_2_io_Stationary_matrix_4_7),
    .io_Stationary_matrix_5_0(PathFinder_2_io_Stationary_matrix_5_0),
    .io_Stationary_matrix_5_1(PathFinder_2_io_Stationary_matrix_5_1),
    .io_Stationary_matrix_5_2(PathFinder_2_io_Stationary_matrix_5_2),
    .io_Stationary_matrix_5_3(PathFinder_2_io_Stationary_matrix_5_3),
    .io_Stationary_matrix_5_4(PathFinder_2_io_Stationary_matrix_5_4),
    .io_Stationary_matrix_5_5(PathFinder_2_io_Stationary_matrix_5_5),
    .io_Stationary_matrix_5_6(PathFinder_2_io_Stationary_matrix_5_6),
    .io_Stationary_matrix_5_7(PathFinder_2_io_Stationary_matrix_5_7),
    .io_Stationary_matrix_6_0(PathFinder_2_io_Stationary_matrix_6_0),
    .io_Stationary_matrix_6_1(PathFinder_2_io_Stationary_matrix_6_1),
    .io_Stationary_matrix_6_2(PathFinder_2_io_Stationary_matrix_6_2),
    .io_Stationary_matrix_6_3(PathFinder_2_io_Stationary_matrix_6_3),
    .io_Stationary_matrix_6_4(PathFinder_2_io_Stationary_matrix_6_4),
    .io_Stationary_matrix_6_5(PathFinder_2_io_Stationary_matrix_6_5),
    .io_Stationary_matrix_6_6(PathFinder_2_io_Stationary_matrix_6_6),
    .io_Stationary_matrix_6_7(PathFinder_2_io_Stationary_matrix_6_7),
    .io_Stationary_matrix_7_0(PathFinder_2_io_Stationary_matrix_7_0),
    .io_Stationary_matrix_7_1(PathFinder_2_io_Stationary_matrix_7_1),
    .io_Stationary_matrix_7_2(PathFinder_2_io_Stationary_matrix_7_2),
    .io_Stationary_matrix_7_3(PathFinder_2_io_Stationary_matrix_7_3),
    .io_Stationary_matrix_7_4(PathFinder_2_io_Stationary_matrix_7_4),
    .io_Stationary_matrix_7_5(PathFinder_2_io_Stationary_matrix_7_5),
    .io_Stationary_matrix_7_6(PathFinder_2_io_Stationary_matrix_7_6),
    .io_Stationary_matrix_7_7(PathFinder_2_io_Stationary_matrix_7_7),
    .io_Streaming_matrix_0(PathFinder_2_io_Streaming_matrix_0),
    .io_Streaming_matrix_1(PathFinder_2_io_Streaming_matrix_1),
    .io_Streaming_matrix_2(PathFinder_2_io_Streaming_matrix_2),
    .io_Streaming_matrix_3(PathFinder_2_io_Streaming_matrix_3),
    .io_Streaming_matrix_4(PathFinder_2_io_Streaming_matrix_4),
    .io_Streaming_matrix_5(PathFinder_2_io_Streaming_matrix_5),
    .io_Streaming_matrix_6(PathFinder_2_io_Streaming_matrix_6),
    .io_Streaming_matrix_7(PathFinder_2_io_Streaming_matrix_7),
    .io_i_mux_bus_0(PathFinder_2_io_i_mux_bus_0),
    .io_i_mux_bus_1(PathFinder_2_io_i_mux_bus_1),
    .io_i_mux_bus_2(PathFinder_2_io_i_mux_bus_2),
    .io_i_mux_bus_3(PathFinder_2_io_i_mux_bus_3),
    .io_Source_0(PathFinder_2_io_Source_0),
    .io_Source_1(PathFinder_2_io_Source_1),
    .io_Source_2(PathFinder_2_io_Source_2),
    .io_Source_3(PathFinder_2_io_Source_3),
    .io_PF_Valid(PathFinder_2_io_PF_Valid),
    .io_NoDPE(PathFinder_2_io_NoDPE),
    .io_DataValid(PathFinder_2_io_DataValid)
  );
  PathFinder PathFinder_3 ( // @[FlexDPU.scala 77:41]
    .clock(PathFinder_3_clock),
    .reset(PathFinder_3_reset),
    .io_Stationary_matrix_0_0(PathFinder_3_io_Stationary_matrix_0_0),
    .io_Stationary_matrix_0_1(PathFinder_3_io_Stationary_matrix_0_1),
    .io_Stationary_matrix_0_2(PathFinder_3_io_Stationary_matrix_0_2),
    .io_Stationary_matrix_0_3(PathFinder_3_io_Stationary_matrix_0_3),
    .io_Stationary_matrix_0_4(PathFinder_3_io_Stationary_matrix_0_4),
    .io_Stationary_matrix_0_5(PathFinder_3_io_Stationary_matrix_0_5),
    .io_Stationary_matrix_0_6(PathFinder_3_io_Stationary_matrix_0_6),
    .io_Stationary_matrix_0_7(PathFinder_3_io_Stationary_matrix_0_7),
    .io_Stationary_matrix_1_0(PathFinder_3_io_Stationary_matrix_1_0),
    .io_Stationary_matrix_1_1(PathFinder_3_io_Stationary_matrix_1_1),
    .io_Stationary_matrix_1_2(PathFinder_3_io_Stationary_matrix_1_2),
    .io_Stationary_matrix_1_3(PathFinder_3_io_Stationary_matrix_1_3),
    .io_Stationary_matrix_1_4(PathFinder_3_io_Stationary_matrix_1_4),
    .io_Stationary_matrix_1_5(PathFinder_3_io_Stationary_matrix_1_5),
    .io_Stationary_matrix_1_6(PathFinder_3_io_Stationary_matrix_1_6),
    .io_Stationary_matrix_1_7(PathFinder_3_io_Stationary_matrix_1_7),
    .io_Stationary_matrix_2_0(PathFinder_3_io_Stationary_matrix_2_0),
    .io_Stationary_matrix_2_1(PathFinder_3_io_Stationary_matrix_2_1),
    .io_Stationary_matrix_2_2(PathFinder_3_io_Stationary_matrix_2_2),
    .io_Stationary_matrix_2_3(PathFinder_3_io_Stationary_matrix_2_3),
    .io_Stationary_matrix_2_4(PathFinder_3_io_Stationary_matrix_2_4),
    .io_Stationary_matrix_2_5(PathFinder_3_io_Stationary_matrix_2_5),
    .io_Stationary_matrix_2_6(PathFinder_3_io_Stationary_matrix_2_6),
    .io_Stationary_matrix_2_7(PathFinder_3_io_Stationary_matrix_2_7),
    .io_Stationary_matrix_3_0(PathFinder_3_io_Stationary_matrix_3_0),
    .io_Stationary_matrix_3_1(PathFinder_3_io_Stationary_matrix_3_1),
    .io_Stationary_matrix_3_2(PathFinder_3_io_Stationary_matrix_3_2),
    .io_Stationary_matrix_3_3(PathFinder_3_io_Stationary_matrix_3_3),
    .io_Stationary_matrix_3_4(PathFinder_3_io_Stationary_matrix_3_4),
    .io_Stationary_matrix_3_5(PathFinder_3_io_Stationary_matrix_3_5),
    .io_Stationary_matrix_3_6(PathFinder_3_io_Stationary_matrix_3_6),
    .io_Stationary_matrix_3_7(PathFinder_3_io_Stationary_matrix_3_7),
    .io_Stationary_matrix_4_0(PathFinder_3_io_Stationary_matrix_4_0),
    .io_Stationary_matrix_4_1(PathFinder_3_io_Stationary_matrix_4_1),
    .io_Stationary_matrix_4_2(PathFinder_3_io_Stationary_matrix_4_2),
    .io_Stationary_matrix_4_3(PathFinder_3_io_Stationary_matrix_4_3),
    .io_Stationary_matrix_4_4(PathFinder_3_io_Stationary_matrix_4_4),
    .io_Stationary_matrix_4_5(PathFinder_3_io_Stationary_matrix_4_5),
    .io_Stationary_matrix_4_6(PathFinder_3_io_Stationary_matrix_4_6),
    .io_Stationary_matrix_4_7(PathFinder_3_io_Stationary_matrix_4_7),
    .io_Stationary_matrix_5_0(PathFinder_3_io_Stationary_matrix_5_0),
    .io_Stationary_matrix_5_1(PathFinder_3_io_Stationary_matrix_5_1),
    .io_Stationary_matrix_5_2(PathFinder_3_io_Stationary_matrix_5_2),
    .io_Stationary_matrix_5_3(PathFinder_3_io_Stationary_matrix_5_3),
    .io_Stationary_matrix_5_4(PathFinder_3_io_Stationary_matrix_5_4),
    .io_Stationary_matrix_5_5(PathFinder_3_io_Stationary_matrix_5_5),
    .io_Stationary_matrix_5_6(PathFinder_3_io_Stationary_matrix_5_6),
    .io_Stationary_matrix_5_7(PathFinder_3_io_Stationary_matrix_5_7),
    .io_Stationary_matrix_6_0(PathFinder_3_io_Stationary_matrix_6_0),
    .io_Stationary_matrix_6_1(PathFinder_3_io_Stationary_matrix_6_1),
    .io_Stationary_matrix_6_2(PathFinder_3_io_Stationary_matrix_6_2),
    .io_Stationary_matrix_6_3(PathFinder_3_io_Stationary_matrix_6_3),
    .io_Stationary_matrix_6_4(PathFinder_3_io_Stationary_matrix_6_4),
    .io_Stationary_matrix_6_5(PathFinder_3_io_Stationary_matrix_6_5),
    .io_Stationary_matrix_6_6(PathFinder_3_io_Stationary_matrix_6_6),
    .io_Stationary_matrix_6_7(PathFinder_3_io_Stationary_matrix_6_7),
    .io_Stationary_matrix_7_0(PathFinder_3_io_Stationary_matrix_7_0),
    .io_Stationary_matrix_7_1(PathFinder_3_io_Stationary_matrix_7_1),
    .io_Stationary_matrix_7_2(PathFinder_3_io_Stationary_matrix_7_2),
    .io_Stationary_matrix_7_3(PathFinder_3_io_Stationary_matrix_7_3),
    .io_Stationary_matrix_7_4(PathFinder_3_io_Stationary_matrix_7_4),
    .io_Stationary_matrix_7_5(PathFinder_3_io_Stationary_matrix_7_5),
    .io_Stationary_matrix_7_6(PathFinder_3_io_Stationary_matrix_7_6),
    .io_Stationary_matrix_7_7(PathFinder_3_io_Stationary_matrix_7_7),
    .io_Streaming_matrix_0(PathFinder_3_io_Streaming_matrix_0),
    .io_Streaming_matrix_1(PathFinder_3_io_Streaming_matrix_1),
    .io_Streaming_matrix_2(PathFinder_3_io_Streaming_matrix_2),
    .io_Streaming_matrix_3(PathFinder_3_io_Streaming_matrix_3),
    .io_Streaming_matrix_4(PathFinder_3_io_Streaming_matrix_4),
    .io_Streaming_matrix_5(PathFinder_3_io_Streaming_matrix_5),
    .io_Streaming_matrix_6(PathFinder_3_io_Streaming_matrix_6),
    .io_Streaming_matrix_7(PathFinder_3_io_Streaming_matrix_7),
    .io_i_mux_bus_0(PathFinder_3_io_i_mux_bus_0),
    .io_i_mux_bus_1(PathFinder_3_io_i_mux_bus_1),
    .io_i_mux_bus_2(PathFinder_3_io_i_mux_bus_2),
    .io_i_mux_bus_3(PathFinder_3_io_i_mux_bus_3),
    .io_Source_0(PathFinder_3_io_Source_0),
    .io_Source_1(PathFinder_3_io_Source_1),
    .io_Source_2(PathFinder_3_io_Source_2),
    .io_Source_3(PathFinder_3_io_Source_3),
    .io_PF_Valid(PathFinder_3_io_PF_Valid),
    .io_NoDPE(PathFinder_3_io_NoDPE),
    .io_DataValid(PathFinder_3_io_DataValid)
  );
  PathFinder PathFinder_4 ( // @[FlexDPU.scala 77:41]
    .clock(PathFinder_4_clock),
    .reset(PathFinder_4_reset),
    .io_Stationary_matrix_0_0(PathFinder_4_io_Stationary_matrix_0_0),
    .io_Stationary_matrix_0_1(PathFinder_4_io_Stationary_matrix_0_1),
    .io_Stationary_matrix_0_2(PathFinder_4_io_Stationary_matrix_0_2),
    .io_Stationary_matrix_0_3(PathFinder_4_io_Stationary_matrix_0_3),
    .io_Stationary_matrix_0_4(PathFinder_4_io_Stationary_matrix_0_4),
    .io_Stationary_matrix_0_5(PathFinder_4_io_Stationary_matrix_0_5),
    .io_Stationary_matrix_0_6(PathFinder_4_io_Stationary_matrix_0_6),
    .io_Stationary_matrix_0_7(PathFinder_4_io_Stationary_matrix_0_7),
    .io_Stationary_matrix_1_0(PathFinder_4_io_Stationary_matrix_1_0),
    .io_Stationary_matrix_1_1(PathFinder_4_io_Stationary_matrix_1_1),
    .io_Stationary_matrix_1_2(PathFinder_4_io_Stationary_matrix_1_2),
    .io_Stationary_matrix_1_3(PathFinder_4_io_Stationary_matrix_1_3),
    .io_Stationary_matrix_1_4(PathFinder_4_io_Stationary_matrix_1_4),
    .io_Stationary_matrix_1_5(PathFinder_4_io_Stationary_matrix_1_5),
    .io_Stationary_matrix_1_6(PathFinder_4_io_Stationary_matrix_1_6),
    .io_Stationary_matrix_1_7(PathFinder_4_io_Stationary_matrix_1_7),
    .io_Stationary_matrix_2_0(PathFinder_4_io_Stationary_matrix_2_0),
    .io_Stationary_matrix_2_1(PathFinder_4_io_Stationary_matrix_2_1),
    .io_Stationary_matrix_2_2(PathFinder_4_io_Stationary_matrix_2_2),
    .io_Stationary_matrix_2_3(PathFinder_4_io_Stationary_matrix_2_3),
    .io_Stationary_matrix_2_4(PathFinder_4_io_Stationary_matrix_2_4),
    .io_Stationary_matrix_2_5(PathFinder_4_io_Stationary_matrix_2_5),
    .io_Stationary_matrix_2_6(PathFinder_4_io_Stationary_matrix_2_6),
    .io_Stationary_matrix_2_7(PathFinder_4_io_Stationary_matrix_2_7),
    .io_Stationary_matrix_3_0(PathFinder_4_io_Stationary_matrix_3_0),
    .io_Stationary_matrix_3_1(PathFinder_4_io_Stationary_matrix_3_1),
    .io_Stationary_matrix_3_2(PathFinder_4_io_Stationary_matrix_3_2),
    .io_Stationary_matrix_3_3(PathFinder_4_io_Stationary_matrix_3_3),
    .io_Stationary_matrix_3_4(PathFinder_4_io_Stationary_matrix_3_4),
    .io_Stationary_matrix_3_5(PathFinder_4_io_Stationary_matrix_3_5),
    .io_Stationary_matrix_3_6(PathFinder_4_io_Stationary_matrix_3_6),
    .io_Stationary_matrix_3_7(PathFinder_4_io_Stationary_matrix_3_7),
    .io_Stationary_matrix_4_0(PathFinder_4_io_Stationary_matrix_4_0),
    .io_Stationary_matrix_4_1(PathFinder_4_io_Stationary_matrix_4_1),
    .io_Stationary_matrix_4_2(PathFinder_4_io_Stationary_matrix_4_2),
    .io_Stationary_matrix_4_3(PathFinder_4_io_Stationary_matrix_4_3),
    .io_Stationary_matrix_4_4(PathFinder_4_io_Stationary_matrix_4_4),
    .io_Stationary_matrix_4_5(PathFinder_4_io_Stationary_matrix_4_5),
    .io_Stationary_matrix_4_6(PathFinder_4_io_Stationary_matrix_4_6),
    .io_Stationary_matrix_4_7(PathFinder_4_io_Stationary_matrix_4_7),
    .io_Stationary_matrix_5_0(PathFinder_4_io_Stationary_matrix_5_0),
    .io_Stationary_matrix_5_1(PathFinder_4_io_Stationary_matrix_5_1),
    .io_Stationary_matrix_5_2(PathFinder_4_io_Stationary_matrix_5_2),
    .io_Stationary_matrix_5_3(PathFinder_4_io_Stationary_matrix_5_3),
    .io_Stationary_matrix_5_4(PathFinder_4_io_Stationary_matrix_5_4),
    .io_Stationary_matrix_5_5(PathFinder_4_io_Stationary_matrix_5_5),
    .io_Stationary_matrix_5_6(PathFinder_4_io_Stationary_matrix_5_6),
    .io_Stationary_matrix_5_7(PathFinder_4_io_Stationary_matrix_5_7),
    .io_Stationary_matrix_6_0(PathFinder_4_io_Stationary_matrix_6_0),
    .io_Stationary_matrix_6_1(PathFinder_4_io_Stationary_matrix_6_1),
    .io_Stationary_matrix_6_2(PathFinder_4_io_Stationary_matrix_6_2),
    .io_Stationary_matrix_6_3(PathFinder_4_io_Stationary_matrix_6_3),
    .io_Stationary_matrix_6_4(PathFinder_4_io_Stationary_matrix_6_4),
    .io_Stationary_matrix_6_5(PathFinder_4_io_Stationary_matrix_6_5),
    .io_Stationary_matrix_6_6(PathFinder_4_io_Stationary_matrix_6_6),
    .io_Stationary_matrix_6_7(PathFinder_4_io_Stationary_matrix_6_7),
    .io_Stationary_matrix_7_0(PathFinder_4_io_Stationary_matrix_7_0),
    .io_Stationary_matrix_7_1(PathFinder_4_io_Stationary_matrix_7_1),
    .io_Stationary_matrix_7_2(PathFinder_4_io_Stationary_matrix_7_2),
    .io_Stationary_matrix_7_3(PathFinder_4_io_Stationary_matrix_7_3),
    .io_Stationary_matrix_7_4(PathFinder_4_io_Stationary_matrix_7_4),
    .io_Stationary_matrix_7_5(PathFinder_4_io_Stationary_matrix_7_5),
    .io_Stationary_matrix_7_6(PathFinder_4_io_Stationary_matrix_7_6),
    .io_Stationary_matrix_7_7(PathFinder_4_io_Stationary_matrix_7_7),
    .io_Streaming_matrix_0(PathFinder_4_io_Streaming_matrix_0),
    .io_Streaming_matrix_1(PathFinder_4_io_Streaming_matrix_1),
    .io_Streaming_matrix_2(PathFinder_4_io_Streaming_matrix_2),
    .io_Streaming_matrix_3(PathFinder_4_io_Streaming_matrix_3),
    .io_Streaming_matrix_4(PathFinder_4_io_Streaming_matrix_4),
    .io_Streaming_matrix_5(PathFinder_4_io_Streaming_matrix_5),
    .io_Streaming_matrix_6(PathFinder_4_io_Streaming_matrix_6),
    .io_Streaming_matrix_7(PathFinder_4_io_Streaming_matrix_7),
    .io_i_mux_bus_0(PathFinder_4_io_i_mux_bus_0),
    .io_i_mux_bus_1(PathFinder_4_io_i_mux_bus_1),
    .io_i_mux_bus_2(PathFinder_4_io_i_mux_bus_2),
    .io_i_mux_bus_3(PathFinder_4_io_i_mux_bus_3),
    .io_Source_0(PathFinder_4_io_Source_0),
    .io_Source_1(PathFinder_4_io_Source_1),
    .io_Source_2(PathFinder_4_io_Source_2),
    .io_Source_3(PathFinder_4_io_Source_3),
    .io_PF_Valid(PathFinder_4_io_PF_Valid),
    .io_NoDPE(PathFinder_4_io_NoDPE),
    .io_DataValid(PathFinder_4_io_DataValid)
  );
  PathFinder PathFinder_5 ( // @[FlexDPU.scala 77:41]
    .clock(PathFinder_5_clock),
    .reset(PathFinder_5_reset),
    .io_Stationary_matrix_0_0(PathFinder_5_io_Stationary_matrix_0_0),
    .io_Stationary_matrix_0_1(PathFinder_5_io_Stationary_matrix_0_1),
    .io_Stationary_matrix_0_2(PathFinder_5_io_Stationary_matrix_0_2),
    .io_Stationary_matrix_0_3(PathFinder_5_io_Stationary_matrix_0_3),
    .io_Stationary_matrix_0_4(PathFinder_5_io_Stationary_matrix_0_4),
    .io_Stationary_matrix_0_5(PathFinder_5_io_Stationary_matrix_0_5),
    .io_Stationary_matrix_0_6(PathFinder_5_io_Stationary_matrix_0_6),
    .io_Stationary_matrix_0_7(PathFinder_5_io_Stationary_matrix_0_7),
    .io_Stationary_matrix_1_0(PathFinder_5_io_Stationary_matrix_1_0),
    .io_Stationary_matrix_1_1(PathFinder_5_io_Stationary_matrix_1_1),
    .io_Stationary_matrix_1_2(PathFinder_5_io_Stationary_matrix_1_2),
    .io_Stationary_matrix_1_3(PathFinder_5_io_Stationary_matrix_1_3),
    .io_Stationary_matrix_1_4(PathFinder_5_io_Stationary_matrix_1_4),
    .io_Stationary_matrix_1_5(PathFinder_5_io_Stationary_matrix_1_5),
    .io_Stationary_matrix_1_6(PathFinder_5_io_Stationary_matrix_1_6),
    .io_Stationary_matrix_1_7(PathFinder_5_io_Stationary_matrix_1_7),
    .io_Stationary_matrix_2_0(PathFinder_5_io_Stationary_matrix_2_0),
    .io_Stationary_matrix_2_1(PathFinder_5_io_Stationary_matrix_2_1),
    .io_Stationary_matrix_2_2(PathFinder_5_io_Stationary_matrix_2_2),
    .io_Stationary_matrix_2_3(PathFinder_5_io_Stationary_matrix_2_3),
    .io_Stationary_matrix_2_4(PathFinder_5_io_Stationary_matrix_2_4),
    .io_Stationary_matrix_2_5(PathFinder_5_io_Stationary_matrix_2_5),
    .io_Stationary_matrix_2_6(PathFinder_5_io_Stationary_matrix_2_6),
    .io_Stationary_matrix_2_7(PathFinder_5_io_Stationary_matrix_2_7),
    .io_Stationary_matrix_3_0(PathFinder_5_io_Stationary_matrix_3_0),
    .io_Stationary_matrix_3_1(PathFinder_5_io_Stationary_matrix_3_1),
    .io_Stationary_matrix_3_2(PathFinder_5_io_Stationary_matrix_3_2),
    .io_Stationary_matrix_3_3(PathFinder_5_io_Stationary_matrix_3_3),
    .io_Stationary_matrix_3_4(PathFinder_5_io_Stationary_matrix_3_4),
    .io_Stationary_matrix_3_5(PathFinder_5_io_Stationary_matrix_3_5),
    .io_Stationary_matrix_3_6(PathFinder_5_io_Stationary_matrix_3_6),
    .io_Stationary_matrix_3_7(PathFinder_5_io_Stationary_matrix_3_7),
    .io_Stationary_matrix_4_0(PathFinder_5_io_Stationary_matrix_4_0),
    .io_Stationary_matrix_4_1(PathFinder_5_io_Stationary_matrix_4_1),
    .io_Stationary_matrix_4_2(PathFinder_5_io_Stationary_matrix_4_2),
    .io_Stationary_matrix_4_3(PathFinder_5_io_Stationary_matrix_4_3),
    .io_Stationary_matrix_4_4(PathFinder_5_io_Stationary_matrix_4_4),
    .io_Stationary_matrix_4_5(PathFinder_5_io_Stationary_matrix_4_5),
    .io_Stationary_matrix_4_6(PathFinder_5_io_Stationary_matrix_4_6),
    .io_Stationary_matrix_4_7(PathFinder_5_io_Stationary_matrix_4_7),
    .io_Stationary_matrix_5_0(PathFinder_5_io_Stationary_matrix_5_0),
    .io_Stationary_matrix_5_1(PathFinder_5_io_Stationary_matrix_5_1),
    .io_Stationary_matrix_5_2(PathFinder_5_io_Stationary_matrix_5_2),
    .io_Stationary_matrix_5_3(PathFinder_5_io_Stationary_matrix_5_3),
    .io_Stationary_matrix_5_4(PathFinder_5_io_Stationary_matrix_5_4),
    .io_Stationary_matrix_5_5(PathFinder_5_io_Stationary_matrix_5_5),
    .io_Stationary_matrix_5_6(PathFinder_5_io_Stationary_matrix_5_6),
    .io_Stationary_matrix_5_7(PathFinder_5_io_Stationary_matrix_5_7),
    .io_Stationary_matrix_6_0(PathFinder_5_io_Stationary_matrix_6_0),
    .io_Stationary_matrix_6_1(PathFinder_5_io_Stationary_matrix_6_1),
    .io_Stationary_matrix_6_2(PathFinder_5_io_Stationary_matrix_6_2),
    .io_Stationary_matrix_6_3(PathFinder_5_io_Stationary_matrix_6_3),
    .io_Stationary_matrix_6_4(PathFinder_5_io_Stationary_matrix_6_4),
    .io_Stationary_matrix_6_5(PathFinder_5_io_Stationary_matrix_6_5),
    .io_Stationary_matrix_6_6(PathFinder_5_io_Stationary_matrix_6_6),
    .io_Stationary_matrix_6_7(PathFinder_5_io_Stationary_matrix_6_7),
    .io_Stationary_matrix_7_0(PathFinder_5_io_Stationary_matrix_7_0),
    .io_Stationary_matrix_7_1(PathFinder_5_io_Stationary_matrix_7_1),
    .io_Stationary_matrix_7_2(PathFinder_5_io_Stationary_matrix_7_2),
    .io_Stationary_matrix_7_3(PathFinder_5_io_Stationary_matrix_7_3),
    .io_Stationary_matrix_7_4(PathFinder_5_io_Stationary_matrix_7_4),
    .io_Stationary_matrix_7_5(PathFinder_5_io_Stationary_matrix_7_5),
    .io_Stationary_matrix_7_6(PathFinder_5_io_Stationary_matrix_7_6),
    .io_Stationary_matrix_7_7(PathFinder_5_io_Stationary_matrix_7_7),
    .io_Streaming_matrix_0(PathFinder_5_io_Streaming_matrix_0),
    .io_Streaming_matrix_1(PathFinder_5_io_Streaming_matrix_1),
    .io_Streaming_matrix_2(PathFinder_5_io_Streaming_matrix_2),
    .io_Streaming_matrix_3(PathFinder_5_io_Streaming_matrix_3),
    .io_Streaming_matrix_4(PathFinder_5_io_Streaming_matrix_4),
    .io_Streaming_matrix_5(PathFinder_5_io_Streaming_matrix_5),
    .io_Streaming_matrix_6(PathFinder_5_io_Streaming_matrix_6),
    .io_Streaming_matrix_7(PathFinder_5_io_Streaming_matrix_7),
    .io_i_mux_bus_0(PathFinder_5_io_i_mux_bus_0),
    .io_i_mux_bus_1(PathFinder_5_io_i_mux_bus_1),
    .io_i_mux_bus_2(PathFinder_5_io_i_mux_bus_2),
    .io_i_mux_bus_3(PathFinder_5_io_i_mux_bus_3),
    .io_Source_0(PathFinder_5_io_Source_0),
    .io_Source_1(PathFinder_5_io_Source_1),
    .io_Source_2(PathFinder_5_io_Source_2),
    .io_Source_3(PathFinder_5_io_Source_3),
    .io_PF_Valid(PathFinder_5_io_PF_Valid),
    .io_NoDPE(PathFinder_5_io_NoDPE),
    .io_DataValid(PathFinder_5_io_DataValid)
  );
  PathFinder PathFinder_6 ( // @[FlexDPU.scala 77:41]
    .clock(PathFinder_6_clock),
    .reset(PathFinder_6_reset),
    .io_Stationary_matrix_0_0(PathFinder_6_io_Stationary_matrix_0_0),
    .io_Stationary_matrix_0_1(PathFinder_6_io_Stationary_matrix_0_1),
    .io_Stationary_matrix_0_2(PathFinder_6_io_Stationary_matrix_0_2),
    .io_Stationary_matrix_0_3(PathFinder_6_io_Stationary_matrix_0_3),
    .io_Stationary_matrix_0_4(PathFinder_6_io_Stationary_matrix_0_4),
    .io_Stationary_matrix_0_5(PathFinder_6_io_Stationary_matrix_0_5),
    .io_Stationary_matrix_0_6(PathFinder_6_io_Stationary_matrix_0_6),
    .io_Stationary_matrix_0_7(PathFinder_6_io_Stationary_matrix_0_7),
    .io_Stationary_matrix_1_0(PathFinder_6_io_Stationary_matrix_1_0),
    .io_Stationary_matrix_1_1(PathFinder_6_io_Stationary_matrix_1_1),
    .io_Stationary_matrix_1_2(PathFinder_6_io_Stationary_matrix_1_2),
    .io_Stationary_matrix_1_3(PathFinder_6_io_Stationary_matrix_1_3),
    .io_Stationary_matrix_1_4(PathFinder_6_io_Stationary_matrix_1_4),
    .io_Stationary_matrix_1_5(PathFinder_6_io_Stationary_matrix_1_5),
    .io_Stationary_matrix_1_6(PathFinder_6_io_Stationary_matrix_1_6),
    .io_Stationary_matrix_1_7(PathFinder_6_io_Stationary_matrix_1_7),
    .io_Stationary_matrix_2_0(PathFinder_6_io_Stationary_matrix_2_0),
    .io_Stationary_matrix_2_1(PathFinder_6_io_Stationary_matrix_2_1),
    .io_Stationary_matrix_2_2(PathFinder_6_io_Stationary_matrix_2_2),
    .io_Stationary_matrix_2_3(PathFinder_6_io_Stationary_matrix_2_3),
    .io_Stationary_matrix_2_4(PathFinder_6_io_Stationary_matrix_2_4),
    .io_Stationary_matrix_2_5(PathFinder_6_io_Stationary_matrix_2_5),
    .io_Stationary_matrix_2_6(PathFinder_6_io_Stationary_matrix_2_6),
    .io_Stationary_matrix_2_7(PathFinder_6_io_Stationary_matrix_2_7),
    .io_Stationary_matrix_3_0(PathFinder_6_io_Stationary_matrix_3_0),
    .io_Stationary_matrix_3_1(PathFinder_6_io_Stationary_matrix_3_1),
    .io_Stationary_matrix_3_2(PathFinder_6_io_Stationary_matrix_3_2),
    .io_Stationary_matrix_3_3(PathFinder_6_io_Stationary_matrix_3_3),
    .io_Stationary_matrix_3_4(PathFinder_6_io_Stationary_matrix_3_4),
    .io_Stationary_matrix_3_5(PathFinder_6_io_Stationary_matrix_3_5),
    .io_Stationary_matrix_3_6(PathFinder_6_io_Stationary_matrix_3_6),
    .io_Stationary_matrix_3_7(PathFinder_6_io_Stationary_matrix_3_7),
    .io_Stationary_matrix_4_0(PathFinder_6_io_Stationary_matrix_4_0),
    .io_Stationary_matrix_4_1(PathFinder_6_io_Stationary_matrix_4_1),
    .io_Stationary_matrix_4_2(PathFinder_6_io_Stationary_matrix_4_2),
    .io_Stationary_matrix_4_3(PathFinder_6_io_Stationary_matrix_4_3),
    .io_Stationary_matrix_4_4(PathFinder_6_io_Stationary_matrix_4_4),
    .io_Stationary_matrix_4_5(PathFinder_6_io_Stationary_matrix_4_5),
    .io_Stationary_matrix_4_6(PathFinder_6_io_Stationary_matrix_4_6),
    .io_Stationary_matrix_4_7(PathFinder_6_io_Stationary_matrix_4_7),
    .io_Stationary_matrix_5_0(PathFinder_6_io_Stationary_matrix_5_0),
    .io_Stationary_matrix_5_1(PathFinder_6_io_Stationary_matrix_5_1),
    .io_Stationary_matrix_5_2(PathFinder_6_io_Stationary_matrix_5_2),
    .io_Stationary_matrix_5_3(PathFinder_6_io_Stationary_matrix_5_3),
    .io_Stationary_matrix_5_4(PathFinder_6_io_Stationary_matrix_5_4),
    .io_Stationary_matrix_5_5(PathFinder_6_io_Stationary_matrix_5_5),
    .io_Stationary_matrix_5_6(PathFinder_6_io_Stationary_matrix_5_6),
    .io_Stationary_matrix_5_7(PathFinder_6_io_Stationary_matrix_5_7),
    .io_Stationary_matrix_6_0(PathFinder_6_io_Stationary_matrix_6_0),
    .io_Stationary_matrix_6_1(PathFinder_6_io_Stationary_matrix_6_1),
    .io_Stationary_matrix_6_2(PathFinder_6_io_Stationary_matrix_6_2),
    .io_Stationary_matrix_6_3(PathFinder_6_io_Stationary_matrix_6_3),
    .io_Stationary_matrix_6_4(PathFinder_6_io_Stationary_matrix_6_4),
    .io_Stationary_matrix_6_5(PathFinder_6_io_Stationary_matrix_6_5),
    .io_Stationary_matrix_6_6(PathFinder_6_io_Stationary_matrix_6_6),
    .io_Stationary_matrix_6_7(PathFinder_6_io_Stationary_matrix_6_7),
    .io_Stationary_matrix_7_0(PathFinder_6_io_Stationary_matrix_7_0),
    .io_Stationary_matrix_7_1(PathFinder_6_io_Stationary_matrix_7_1),
    .io_Stationary_matrix_7_2(PathFinder_6_io_Stationary_matrix_7_2),
    .io_Stationary_matrix_7_3(PathFinder_6_io_Stationary_matrix_7_3),
    .io_Stationary_matrix_7_4(PathFinder_6_io_Stationary_matrix_7_4),
    .io_Stationary_matrix_7_5(PathFinder_6_io_Stationary_matrix_7_5),
    .io_Stationary_matrix_7_6(PathFinder_6_io_Stationary_matrix_7_6),
    .io_Stationary_matrix_7_7(PathFinder_6_io_Stationary_matrix_7_7),
    .io_Streaming_matrix_0(PathFinder_6_io_Streaming_matrix_0),
    .io_Streaming_matrix_1(PathFinder_6_io_Streaming_matrix_1),
    .io_Streaming_matrix_2(PathFinder_6_io_Streaming_matrix_2),
    .io_Streaming_matrix_3(PathFinder_6_io_Streaming_matrix_3),
    .io_Streaming_matrix_4(PathFinder_6_io_Streaming_matrix_4),
    .io_Streaming_matrix_5(PathFinder_6_io_Streaming_matrix_5),
    .io_Streaming_matrix_6(PathFinder_6_io_Streaming_matrix_6),
    .io_Streaming_matrix_7(PathFinder_6_io_Streaming_matrix_7),
    .io_i_mux_bus_0(PathFinder_6_io_i_mux_bus_0),
    .io_i_mux_bus_1(PathFinder_6_io_i_mux_bus_1),
    .io_i_mux_bus_2(PathFinder_6_io_i_mux_bus_2),
    .io_i_mux_bus_3(PathFinder_6_io_i_mux_bus_3),
    .io_Source_0(PathFinder_6_io_Source_0),
    .io_Source_1(PathFinder_6_io_Source_1),
    .io_Source_2(PathFinder_6_io_Source_2),
    .io_Source_3(PathFinder_6_io_Source_3),
    .io_PF_Valid(PathFinder_6_io_PF_Valid),
    .io_NoDPE(PathFinder_6_io_NoDPE),
    .io_DataValid(PathFinder_6_io_DataValid)
  );
  PathFinder PathFinder_7 ( // @[FlexDPU.scala 77:41]
    .clock(PathFinder_7_clock),
    .reset(PathFinder_7_reset),
    .io_Stationary_matrix_0_0(PathFinder_7_io_Stationary_matrix_0_0),
    .io_Stationary_matrix_0_1(PathFinder_7_io_Stationary_matrix_0_1),
    .io_Stationary_matrix_0_2(PathFinder_7_io_Stationary_matrix_0_2),
    .io_Stationary_matrix_0_3(PathFinder_7_io_Stationary_matrix_0_3),
    .io_Stationary_matrix_0_4(PathFinder_7_io_Stationary_matrix_0_4),
    .io_Stationary_matrix_0_5(PathFinder_7_io_Stationary_matrix_0_5),
    .io_Stationary_matrix_0_6(PathFinder_7_io_Stationary_matrix_0_6),
    .io_Stationary_matrix_0_7(PathFinder_7_io_Stationary_matrix_0_7),
    .io_Stationary_matrix_1_0(PathFinder_7_io_Stationary_matrix_1_0),
    .io_Stationary_matrix_1_1(PathFinder_7_io_Stationary_matrix_1_1),
    .io_Stationary_matrix_1_2(PathFinder_7_io_Stationary_matrix_1_2),
    .io_Stationary_matrix_1_3(PathFinder_7_io_Stationary_matrix_1_3),
    .io_Stationary_matrix_1_4(PathFinder_7_io_Stationary_matrix_1_4),
    .io_Stationary_matrix_1_5(PathFinder_7_io_Stationary_matrix_1_5),
    .io_Stationary_matrix_1_6(PathFinder_7_io_Stationary_matrix_1_6),
    .io_Stationary_matrix_1_7(PathFinder_7_io_Stationary_matrix_1_7),
    .io_Stationary_matrix_2_0(PathFinder_7_io_Stationary_matrix_2_0),
    .io_Stationary_matrix_2_1(PathFinder_7_io_Stationary_matrix_2_1),
    .io_Stationary_matrix_2_2(PathFinder_7_io_Stationary_matrix_2_2),
    .io_Stationary_matrix_2_3(PathFinder_7_io_Stationary_matrix_2_3),
    .io_Stationary_matrix_2_4(PathFinder_7_io_Stationary_matrix_2_4),
    .io_Stationary_matrix_2_5(PathFinder_7_io_Stationary_matrix_2_5),
    .io_Stationary_matrix_2_6(PathFinder_7_io_Stationary_matrix_2_6),
    .io_Stationary_matrix_2_7(PathFinder_7_io_Stationary_matrix_2_7),
    .io_Stationary_matrix_3_0(PathFinder_7_io_Stationary_matrix_3_0),
    .io_Stationary_matrix_3_1(PathFinder_7_io_Stationary_matrix_3_1),
    .io_Stationary_matrix_3_2(PathFinder_7_io_Stationary_matrix_3_2),
    .io_Stationary_matrix_3_3(PathFinder_7_io_Stationary_matrix_3_3),
    .io_Stationary_matrix_3_4(PathFinder_7_io_Stationary_matrix_3_4),
    .io_Stationary_matrix_3_5(PathFinder_7_io_Stationary_matrix_3_5),
    .io_Stationary_matrix_3_6(PathFinder_7_io_Stationary_matrix_3_6),
    .io_Stationary_matrix_3_7(PathFinder_7_io_Stationary_matrix_3_7),
    .io_Stationary_matrix_4_0(PathFinder_7_io_Stationary_matrix_4_0),
    .io_Stationary_matrix_4_1(PathFinder_7_io_Stationary_matrix_4_1),
    .io_Stationary_matrix_4_2(PathFinder_7_io_Stationary_matrix_4_2),
    .io_Stationary_matrix_4_3(PathFinder_7_io_Stationary_matrix_4_3),
    .io_Stationary_matrix_4_4(PathFinder_7_io_Stationary_matrix_4_4),
    .io_Stationary_matrix_4_5(PathFinder_7_io_Stationary_matrix_4_5),
    .io_Stationary_matrix_4_6(PathFinder_7_io_Stationary_matrix_4_6),
    .io_Stationary_matrix_4_7(PathFinder_7_io_Stationary_matrix_4_7),
    .io_Stationary_matrix_5_0(PathFinder_7_io_Stationary_matrix_5_0),
    .io_Stationary_matrix_5_1(PathFinder_7_io_Stationary_matrix_5_1),
    .io_Stationary_matrix_5_2(PathFinder_7_io_Stationary_matrix_5_2),
    .io_Stationary_matrix_5_3(PathFinder_7_io_Stationary_matrix_5_3),
    .io_Stationary_matrix_5_4(PathFinder_7_io_Stationary_matrix_5_4),
    .io_Stationary_matrix_5_5(PathFinder_7_io_Stationary_matrix_5_5),
    .io_Stationary_matrix_5_6(PathFinder_7_io_Stationary_matrix_5_6),
    .io_Stationary_matrix_5_7(PathFinder_7_io_Stationary_matrix_5_7),
    .io_Stationary_matrix_6_0(PathFinder_7_io_Stationary_matrix_6_0),
    .io_Stationary_matrix_6_1(PathFinder_7_io_Stationary_matrix_6_1),
    .io_Stationary_matrix_6_2(PathFinder_7_io_Stationary_matrix_6_2),
    .io_Stationary_matrix_6_3(PathFinder_7_io_Stationary_matrix_6_3),
    .io_Stationary_matrix_6_4(PathFinder_7_io_Stationary_matrix_6_4),
    .io_Stationary_matrix_6_5(PathFinder_7_io_Stationary_matrix_6_5),
    .io_Stationary_matrix_6_6(PathFinder_7_io_Stationary_matrix_6_6),
    .io_Stationary_matrix_6_7(PathFinder_7_io_Stationary_matrix_6_7),
    .io_Stationary_matrix_7_0(PathFinder_7_io_Stationary_matrix_7_0),
    .io_Stationary_matrix_7_1(PathFinder_7_io_Stationary_matrix_7_1),
    .io_Stationary_matrix_7_2(PathFinder_7_io_Stationary_matrix_7_2),
    .io_Stationary_matrix_7_3(PathFinder_7_io_Stationary_matrix_7_3),
    .io_Stationary_matrix_7_4(PathFinder_7_io_Stationary_matrix_7_4),
    .io_Stationary_matrix_7_5(PathFinder_7_io_Stationary_matrix_7_5),
    .io_Stationary_matrix_7_6(PathFinder_7_io_Stationary_matrix_7_6),
    .io_Stationary_matrix_7_7(PathFinder_7_io_Stationary_matrix_7_7),
    .io_Streaming_matrix_0(PathFinder_7_io_Streaming_matrix_0),
    .io_Streaming_matrix_1(PathFinder_7_io_Streaming_matrix_1),
    .io_Streaming_matrix_2(PathFinder_7_io_Streaming_matrix_2),
    .io_Streaming_matrix_3(PathFinder_7_io_Streaming_matrix_3),
    .io_Streaming_matrix_4(PathFinder_7_io_Streaming_matrix_4),
    .io_Streaming_matrix_5(PathFinder_7_io_Streaming_matrix_5),
    .io_Streaming_matrix_6(PathFinder_7_io_Streaming_matrix_6),
    .io_Streaming_matrix_7(PathFinder_7_io_Streaming_matrix_7),
    .io_i_mux_bus_0(PathFinder_7_io_i_mux_bus_0),
    .io_i_mux_bus_1(PathFinder_7_io_i_mux_bus_1),
    .io_i_mux_bus_2(PathFinder_7_io_i_mux_bus_2),
    .io_i_mux_bus_3(PathFinder_7_io_i_mux_bus_3),
    .io_Source_0(PathFinder_7_io_Source_0),
    .io_Source_1(PathFinder_7_io_Source_1),
    .io_Source_2(PathFinder_7_io_Source_2),
    .io_Source_3(PathFinder_7_io_Source_3),
    .io_PF_Valid(PathFinder_7_io_PF_Valid),
    .io_NoDPE(PathFinder_7_io_NoDPE),
    .io_DataValid(PathFinder_7_io_DataValid)
  );
  PathFinder PathFinder_8 ( // @[FlexDPU.scala 77:41]
    .clock(PathFinder_8_clock),
    .reset(PathFinder_8_reset),
    .io_Stationary_matrix_0_0(PathFinder_8_io_Stationary_matrix_0_0),
    .io_Stationary_matrix_0_1(PathFinder_8_io_Stationary_matrix_0_1),
    .io_Stationary_matrix_0_2(PathFinder_8_io_Stationary_matrix_0_2),
    .io_Stationary_matrix_0_3(PathFinder_8_io_Stationary_matrix_0_3),
    .io_Stationary_matrix_0_4(PathFinder_8_io_Stationary_matrix_0_4),
    .io_Stationary_matrix_0_5(PathFinder_8_io_Stationary_matrix_0_5),
    .io_Stationary_matrix_0_6(PathFinder_8_io_Stationary_matrix_0_6),
    .io_Stationary_matrix_0_7(PathFinder_8_io_Stationary_matrix_0_7),
    .io_Stationary_matrix_1_0(PathFinder_8_io_Stationary_matrix_1_0),
    .io_Stationary_matrix_1_1(PathFinder_8_io_Stationary_matrix_1_1),
    .io_Stationary_matrix_1_2(PathFinder_8_io_Stationary_matrix_1_2),
    .io_Stationary_matrix_1_3(PathFinder_8_io_Stationary_matrix_1_3),
    .io_Stationary_matrix_1_4(PathFinder_8_io_Stationary_matrix_1_4),
    .io_Stationary_matrix_1_5(PathFinder_8_io_Stationary_matrix_1_5),
    .io_Stationary_matrix_1_6(PathFinder_8_io_Stationary_matrix_1_6),
    .io_Stationary_matrix_1_7(PathFinder_8_io_Stationary_matrix_1_7),
    .io_Stationary_matrix_2_0(PathFinder_8_io_Stationary_matrix_2_0),
    .io_Stationary_matrix_2_1(PathFinder_8_io_Stationary_matrix_2_1),
    .io_Stationary_matrix_2_2(PathFinder_8_io_Stationary_matrix_2_2),
    .io_Stationary_matrix_2_3(PathFinder_8_io_Stationary_matrix_2_3),
    .io_Stationary_matrix_2_4(PathFinder_8_io_Stationary_matrix_2_4),
    .io_Stationary_matrix_2_5(PathFinder_8_io_Stationary_matrix_2_5),
    .io_Stationary_matrix_2_6(PathFinder_8_io_Stationary_matrix_2_6),
    .io_Stationary_matrix_2_7(PathFinder_8_io_Stationary_matrix_2_7),
    .io_Stationary_matrix_3_0(PathFinder_8_io_Stationary_matrix_3_0),
    .io_Stationary_matrix_3_1(PathFinder_8_io_Stationary_matrix_3_1),
    .io_Stationary_matrix_3_2(PathFinder_8_io_Stationary_matrix_3_2),
    .io_Stationary_matrix_3_3(PathFinder_8_io_Stationary_matrix_3_3),
    .io_Stationary_matrix_3_4(PathFinder_8_io_Stationary_matrix_3_4),
    .io_Stationary_matrix_3_5(PathFinder_8_io_Stationary_matrix_3_5),
    .io_Stationary_matrix_3_6(PathFinder_8_io_Stationary_matrix_3_6),
    .io_Stationary_matrix_3_7(PathFinder_8_io_Stationary_matrix_3_7),
    .io_Stationary_matrix_4_0(PathFinder_8_io_Stationary_matrix_4_0),
    .io_Stationary_matrix_4_1(PathFinder_8_io_Stationary_matrix_4_1),
    .io_Stationary_matrix_4_2(PathFinder_8_io_Stationary_matrix_4_2),
    .io_Stationary_matrix_4_3(PathFinder_8_io_Stationary_matrix_4_3),
    .io_Stationary_matrix_4_4(PathFinder_8_io_Stationary_matrix_4_4),
    .io_Stationary_matrix_4_5(PathFinder_8_io_Stationary_matrix_4_5),
    .io_Stationary_matrix_4_6(PathFinder_8_io_Stationary_matrix_4_6),
    .io_Stationary_matrix_4_7(PathFinder_8_io_Stationary_matrix_4_7),
    .io_Stationary_matrix_5_0(PathFinder_8_io_Stationary_matrix_5_0),
    .io_Stationary_matrix_5_1(PathFinder_8_io_Stationary_matrix_5_1),
    .io_Stationary_matrix_5_2(PathFinder_8_io_Stationary_matrix_5_2),
    .io_Stationary_matrix_5_3(PathFinder_8_io_Stationary_matrix_5_3),
    .io_Stationary_matrix_5_4(PathFinder_8_io_Stationary_matrix_5_4),
    .io_Stationary_matrix_5_5(PathFinder_8_io_Stationary_matrix_5_5),
    .io_Stationary_matrix_5_6(PathFinder_8_io_Stationary_matrix_5_6),
    .io_Stationary_matrix_5_7(PathFinder_8_io_Stationary_matrix_5_7),
    .io_Stationary_matrix_6_0(PathFinder_8_io_Stationary_matrix_6_0),
    .io_Stationary_matrix_6_1(PathFinder_8_io_Stationary_matrix_6_1),
    .io_Stationary_matrix_6_2(PathFinder_8_io_Stationary_matrix_6_2),
    .io_Stationary_matrix_6_3(PathFinder_8_io_Stationary_matrix_6_3),
    .io_Stationary_matrix_6_4(PathFinder_8_io_Stationary_matrix_6_4),
    .io_Stationary_matrix_6_5(PathFinder_8_io_Stationary_matrix_6_5),
    .io_Stationary_matrix_6_6(PathFinder_8_io_Stationary_matrix_6_6),
    .io_Stationary_matrix_6_7(PathFinder_8_io_Stationary_matrix_6_7),
    .io_Stationary_matrix_7_0(PathFinder_8_io_Stationary_matrix_7_0),
    .io_Stationary_matrix_7_1(PathFinder_8_io_Stationary_matrix_7_1),
    .io_Stationary_matrix_7_2(PathFinder_8_io_Stationary_matrix_7_2),
    .io_Stationary_matrix_7_3(PathFinder_8_io_Stationary_matrix_7_3),
    .io_Stationary_matrix_7_4(PathFinder_8_io_Stationary_matrix_7_4),
    .io_Stationary_matrix_7_5(PathFinder_8_io_Stationary_matrix_7_5),
    .io_Stationary_matrix_7_6(PathFinder_8_io_Stationary_matrix_7_6),
    .io_Stationary_matrix_7_7(PathFinder_8_io_Stationary_matrix_7_7),
    .io_Streaming_matrix_0(PathFinder_8_io_Streaming_matrix_0),
    .io_Streaming_matrix_1(PathFinder_8_io_Streaming_matrix_1),
    .io_Streaming_matrix_2(PathFinder_8_io_Streaming_matrix_2),
    .io_Streaming_matrix_3(PathFinder_8_io_Streaming_matrix_3),
    .io_Streaming_matrix_4(PathFinder_8_io_Streaming_matrix_4),
    .io_Streaming_matrix_5(PathFinder_8_io_Streaming_matrix_5),
    .io_Streaming_matrix_6(PathFinder_8_io_Streaming_matrix_6),
    .io_Streaming_matrix_7(PathFinder_8_io_Streaming_matrix_7),
    .io_i_mux_bus_0(PathFinder_8_io_i_mux_bus_0),
    .io_i_mux_bus_1(PathFinder_8_io_i_mux_bus_1),
    .io_i_mux_bus_2(PathFinder_8_io_i_mux_bus_2),
    .io_i_mux_bus_3(PathFinder_8_io_i_mux_bus_3),
    .io_Source_0(PathFinder_8_io_Source_0),
    .io_Source_1(PathFinder_8_io_Source_1),
    .io_Source_2(PathFinder_8_io_Source_2),
    .io_Source_3(PathFinder_8_io_Source_3),
    .io_PF_Valid(PathFinder_8_io_PF_Valid),
    .io_NoDPE(PathFinder_8_io_NoDPE),
    .io_DataValid(PathFinder_8_io_DataValid)
  );
  PathFinder PathFinder_9 ( // @[FlexDPU.scala 77:41]
    .clock(PathFinder_9_clock),
    .reset(PathFinder_9_reset),
    .io_Stationary_matrix_0_0(PathFinder_9_io_Stationary_matrix_0_0),
    .io_Stationary_matrix_0_1(PathFinder_9_io_Stationary_matrix_0_1),
    .io_Stationary_matrix_0_2(PathFinder_9_io_Stationary_matrix_0_2),
    .io_Stationary_matrix_0_3(PathFinder_9_io_Stationary_matrix_0_3),
    .io_Stationary_matrix_0_4(PathFinder_9_io_Stationary_matrix_0_4),
    .io_Stationary_matrix_0_5(PathFinder_9_io_Stationary_matrix_0_5),
    .io_Stationary_matrix_0_6(PathFinder_9_io_Stationary_matrix_0_6),
    .io_Stationary_matrix_0_7(PathFinder_9_io_Stationary_matrix_0_7),
    .io_Stationary_matrix_1_0(PathFinder_9_io_Stationary_matrix_1_0),
    .io_Stationary_matrix_1_1(PathFinder_9_io_Stationary_matrix_1_1),
    .io_Stationary_matrix_1_2(PathFinder_9_io_Stationary_matrix_1_2),
    .io_Stationary_matrix_1_3(PathFinder_9_io_Stationary_matrix_1_3),
    .io_Stationary_matrix_1_4(PathFinder_9_io_Stationary_matrix_1_4),
    .io_Stationary_matrix_1_5(PathFinder_9_io_Stationary_matrix_1_5),
    .io_Stationary_matrix_1_6(PathFinder_9_io_Stationary_matrix_1_6),
    .io_Stationary_matrix_1_7(PathFinder_9_io_Stationary_matrix_1_7),
    .io_Stationary_matrix_2_0(PathFinder_9_io_Stationary_matrix_2_0),
    .io_Stationary_matrix_2_1(PathFinder_9_io_Stationary_matrix_2_1),
    .io_Stationary_matrix_2_2(PathFinder_9_io_Stationary_matrix_2_2),
    .io_Stationary_matrix_2_3(PathFinder_9_io_Stationary_matrix_2_3),
    .io_Stationary_matrix_2_4(PathFinder_9_io_Stationary_matrix_2_4),
    .io_Stationary_matrix_2_5(PathFinder_9_io_Stationary_matrix_2_5),
    .io_Stationary_matrix_2_6(PathFinder_9_io_Stationary_matrix_2_6),
    .io_Stationary_matrix_2_7(PathFinder_9_io_Stationary_matrix_2_7),
    .io_Stationary_matrix_3_0(PathFinder_9_io_Stationary_matrix_3_0),
    .io_Stationary_matrix_3_1(PathFinder_9_io_Stationary_matrix_3_1),
    .io_Stationary_matrix_3_2(PathFinder_9_io_Stationary_matrix_3_2),
    .io_Stationary_matrix_3_3(PathFinder_9_io_Stationary_matrix_3_3),
    .io_Stationary_matrix_3_4(PathFinder_9_io_Stationary_matrix_3_4),
    .io_Stationary_matrix_3_5(PathFinder_9_io_Stationary_matrix_3_5),
    .io_Stationary_matrix_3_6(PathFinder_9_io_Stationary_matrix_3_6),
    .io_Stationary_matrix_3_7(PathFinder_9_io_Stationary_matrix_3_7),
    .io_Stationary_matrix_4_0(PathFinder_9_io_Stationary_matrix_4_0),
    .io_Stationary_matrix_4_1(PathFinder_9_io_Stationary_matrix_4_1),
    .io_Stationary_matrix_4_2(PathFinder_9_io_Stationary_matrix_4_2),
    .io_Stationary_matrix_4_3(PathFinder_9_io_Stationary_matrix_4_3),
    .io_Stationary_matrix_4_4(PathFinder_9_io_Stationary_matrix_4_4),
    .io_Stationary_matrix_4_5(PathFinder_9_io_Stationary_matrix_4_5),
    .io_Stationary_matrix_4_6(PathFinder_9_io_Stationary_matrix_4_6),
    .io_Stationary_matrix_4_7(PathFinder_9_io_Stationary_matrix_4_7),
    .io_Stationary_matrix_5_0(PathFinder_9_io_Stationary_matrix_5_0),
    .io_Stationary_matrix_5_1(PathFinder_9_io_Stationary_matrix_5_1),
    .io_Stationary_matrix_5_2(PathFinder_9_io_Stationary_matrix_5_2),
    .io_Stationary_matrix_5_3(PathFinder_9_io_Stationary_matrix_5_3),
    .io_Stationary_matrix_5_4(PathFinder_9_io_Stationary_matrix_5_4),
    .io_Stationary_matrix_5_5(PathFinder_9_io_Stationary_matrix_5_5),
    .io_Stationary_matrix_5_6(PathFinder_9_io_Stationary_matrix_5_6),
    .io_Stationary_matrix_5_7(PathFinder_9_io_Stationary_matrix_5_7),
    .io_Stationary_matrix_6_0(PathFinder_9_io_Stationary_matrix_6_0),
    .io_Stationary_matrix_6_1(PathFinder_9_io_Stationary_matrix_6_1),
    .io_Stationary_matrix_6_2(PathFinder_9_io_Stationary_matrix_6_2),
    .io_Stationary_matrix_6_3(PathFinder_9_io_Stationary_matrix_6_3),
    .io_Stationary_matrix_6_4(PathFinder_9_io_Stationary_matrix_6_4),
    .io_Stationary_matrix_6_5(PathFinder_9_io_Stationary_matrix_6_5),
    .io_Stationary_matrix_6_6(PathFinder_9_io_Stationary_matrix_6_6),
    .io_Stationary_matrix_6_7(PathFinder_9_io_Stationary_matrix_6_7),
    .io_Stationary_matrix_7_0(PathFinder_9_io_Stationary_matrix_7_0),
    .io_Stationary_matrix_7_1(PathFinder_9_io_Stationary_matrix_7_1),
    .io_Stationary_matrix_7_2(PathFinder_9_io_Stationary_matrix_7_2),
    .io_Stationary_matrix_7_3(PathFinder_9_io_Stationary_matrix_7_3),
    .io_Stationary_matrix_7_4(PathFinder_9_io_Stationary_matrix_7_4),
    .io_Stationary_matrix_7_5(PathFinder_9_io_Stationary_matrix_7_5),
    .io_Stationary_matrix_7_6(PathFinder_9_io_Stationary_matrix_7_6),
    .io_Stationary_matrix_7_7(PathFinder_9_io_Stationary_matrix_7_7),
    .io_Streaming_matrix_0(PathFinder_9_io_Streaming_matrix_0),
    .io_Streaming_matrix_1(PathFinder_9_io_Streaming_matrix_1),
    .io_Streaming_matrix_2(PathFinder_9_io_Streaming_matrix_2),
    .io_Streaming_matrix_3(PathFinder_9_io_Streaming_matrix_3),
    .io_Streaming_matrix_4(PathFinder_9_io_Streaming_matrix_4),
    .io_Streaming_matrix_5(PathFinder_9_io_Streaming_matrix_5),
    .io_Streaming_matrix_6(PathFinder_9_io_Streaming_matrix_6),
    .io_Streaming_matrix_7(PathFinder_9_io_Streaming_matrix_7),
    .io_i_mux_bus_0(PathFinder_9_io_i_mux_bus_0),
    .io_i_mux_bus_1(PathFinder_9_io_i_mux_bus_1),
    .io_i_mux_bus_2(PathFinder_9_io_i_mux_bus_2),
    .io_i_mux_bus_3(PathFinder_9_io_i_mux_bus_3),
    .io_Source_0(PathFinder_9_io_Source_0),
    .io_Source_1(PathFinder_9_io_Source_1),
    .io_Source_2(PathFinder_9_io_Source_2),
    .io_Source_3(PathFinder_9_io_Source_3),
    .io_PF_Valid(PathFinder_9_io_PF_Valid),
    .io_NoDPE(PathFinder_9_io_NoDPE),
    .io_DataValid(PathFinder_9_io_DataValid)
  );
  PathFinder PathFinder_10 ( // @[FlexDPU.scala 77:41]
    .clock(PathFinder_10_clock),
    .reset(PathFinder_10_reset),
    .io_Stationary_matrix_0_0(PathFinder_10_io_Stationary_matrix_0_0),
    .io_Stationary_matrix_0_1(PathFinder_10_io_Stationary_matrix_0_1),
    .io_Stationary_matrix_0_2(PathFinder_10_io_Stationary_matrix_0_2),
    .io_Stationary_matrix_0_3(PathFinder_10_io_Stationary_matrix_0_3),
    .io_Stationary_matrix_0_4(PathFinder_10_io_Stationary_matrix_0_4),
    .io_Stationary_matrix_0_5(PathFinder_10_io_Stationary_matrix_0_5),
    .io_Stationary_matrix_0_6(PathFinder_10_io_Stationary_matrix_0_6),
    .io_Stationary_matrix_0_7(PathFinder_10_io_Stationary_matrix_0_7),
    .io_Stationary_matrix_1_0(PathFinder_10_io_Stationary_matrix_1_0),
    .io_Stationary_matrix_1_1(PathFinder_10_io_Stationary_matrix_1_1),
    .io_Stationary_matrix_1_2(PathFinder_10_io_Stationary_matrix_1_2),
    .io_Stationary_matrix_1_3(PathFinder_10_io_Stationary_matrix_1_3),
    .io_Stationary_matrix_1_4(PathFinder_10_io_Stationary_matrix_1_4),
    .io_Stationary_matrix_1_5(PathFinder_10_io_Stationary_matrix_1_5),
    .io_Stationary_matrix_1_6(PathFinder_10_io_Stationary_matrix_1_6),
    .io_Stationary_matrix_1_7(PathFinder_10_io_Stationary_matrix_1_7),
    .io_Stationary_matrix_2_0(PathFinder_10_io_Stationary_matrix_2_0),
    .io_Stationary_matrix_2_1(PathFinder_10_io_Stationary_matrix_2_1),
    .io_Stationary_matrix_2_2(PathFinder_10_io_Stationary_matrix_2_2),
    .io_Stationary_matrix_2_3(PathFinder_10_io_Stationary_matrix_2_3),
    .io_Stationary_matrix_2_4(PathFinder_10_io_Stationary_matrix_2_4),
    .io_Stationary_matrix_2_5(PathFinder_10_io_Stationary_matrix_2_5),
    .io_Stationary_matrix_2_6(PathFinder_10_io_Stationary_matrix_2_6),
    .io_Stationary_matrix_2_7(PathFinder_10_io_Stationary_matrix_2_7),
    .io_Stationary_matrix_3_0(PathFinder_10_io_Stationary_matrix_3_0),
    .io_Stationary_matrix_3_1(PathFinder_10_io_Stationary_matrix_3_1),
    .io_Stationary_matrix_3_2(PathFinder_10_io_Stationary_matrix_3_2),
    .io_Stationary_matrix_3_3(PathFinder_10_io_Stationary_matrix_3_3),
    .io_Stationary_matrix_3_4(PathFinder_10_io_Stationary_matrix_3_4),
    .io_Stationary_matrix_3_5(PathFinder_10_io_Stationary_matrix_3_5),
    .io_Stationary_matrix_3_6(PathFinder_10_io_Stationary_matrix_3_6),
    .io_Stationary_matrix_3_7(PathFinder_10_io_Stationary_matrix_3_7),
    .io_Stationary_matrix_4_0(PathFinder_10_io_Stationary_matrix_4_0),
    .io_Stationary_matrix_4_1(PathFinder_10_io_Stationary_matrix_4_1),
    .io_Stationary_matrix_4_2(PathFinder_10_io_Stationary_matrix_4_2),
    .io_Stationary_matrix_4_3(PathFinder_10_io_Stationary_matrix_4_3),
    .io_Stationary_matrix_4_4(PathFinder_10_io_Stationary_matrix_4_4),
    .io_Stationary_matrix_4_5(PathFinder_10_io_Stationary_matrix_4_5),
    .io_Stationary_matrix_4_6(PathFinder_10_io_Stationary_matrix_4_6),
    .io_Stationary_matrix_4_7(PathFinder_10_io_Stationary_matrix_4_7),
    .io_Stationary_matrix_5_0(PathFinder_10_io_Stationary_matrix_5_0),
    .io_Stationary_matrix_5_1(PathFinder_10_io_Stationary_matrix_5_1),
    .io_Stationary_matrix_5_2(PathFinder_10_io_Stationary_matrix_5_2),
    .io_Stationary_matrix_5_3(PathFinder_10_io_Stationary_matrix_5_3),
    .io_Stationary_matrix_5_4(PathFinder_10_io_Stationary_matrix_5_4),
    .io_Stationary_matrix_5_5(PathFinder_10_io_Stationary_matrix_5_5),
    .io_Stationary_matrix_5_6(PathFinder_10_io_Stationary_matrix_5_6),
    .io_Stationary_matrix_5_7(PathFinder_10_io_Stationary_matrix_5_7),
    .io_Stationary_matrix_6_0(PathFinder_10_io_Stationary_matrix_6_0),
    .io_Stationary_matrix_6_1(PathFinder_10_io_Stationary_matrix_6_1),
    .io_Stationary_matrix_6_2(PathFinder_10_io_Stationary_matrix_6_2),
    .io_Stationary_matrix_6_3(PathFinder_10_io_Stationary_matrix_6_3),
    .io_Stationary_matrix_6_4(PathFinder_10_io_Stationary_matrix_6_4),
    .io_Stationary_matrix_6_5(PathFinder_10_io_Stationary_matrix_6_5),
    .io_Stationary_matrix_6_6(PathFinder_10_io_Stationary_matrix_6_6),
    .io_Stationary_matrix_6_7(PathFinder_10_io_Stationary_matrix_6_7),
    .io_Stationary_matrix_7_0(PathFinder_10_io_Stationary_matrix_7_0),
    .io_Stationary_matrix_7_1(PathFinder_10_io_Stationary_matrix_7_1),
    .io_Stationary_matrix_7_2(PathFinder_10_io_Stationary_matrix_7_2),
    .io_Stationary_matrix_7_3(PathFinder_10_io_Stationary_matrix_7_3),
    .io_Stationary_matrix_7_4(PathFinder_10_io_Stationary_matrix_7_4),
    .io_Stationary_matrix_7_5(PathFinder_10_io_Stationary_matrix_7_5),
    .io_Stationary_matrix_7_6(PathFinder_10_io_Stationary_matrix_7_6),
    .io_Stationary_matrix_7_7(PathFinder_10_io_Stationary_matrix_7_7),
    .io_Streaming_matrix_0(PathFinder_10_io_Streaming_matrix_0),
    .io_Streaming_matrix_1(PathFinder_10_io_Streaming_matrix_1),
    .io_Streaming_matrix_2(PathFinder_10_io_Streaming_matrix_2),
    .io_Streaming_matrix_3(PathFinder_10_io_Streaming_matrix_3),
    .io_Streaming_matrix_4(PathFinder_10_io_Streaming_matrix_4),
    .io_Streaming_matrix_5(PathFinder_10_io_Streaming_matrix_5),
    .io_Streaming_matrix_6(PathFinder_10_io_Streaming_matrix_6),
    .io_Streaming_matrix_7(PathFinder_10_io_Streaming_matrix_7),
    .io_i_mux_bus_0(PathFinder_10_io_i_mux_bus_0),
    .io_i_mux_bus_1(PathFinder_10_io_i_mux_bus_1),
    .io_i_mux_bus_2(PathFinder_10_io_i_mux_bus_2),
    .io_i_mux_bus_3(PathFinder_10_io_i_mux_bus_3),
    .io_Source_0(PathFinder_10_io_Source_0),
    .io_Source_1(PathFinder_10_io_Source_1),
    .io_Source_2(PathFinder_10_io_Source_2),
    .io_Source_3(PathFinder_10_io_Source_3),
    .io_PF_Valid(PathFinder_10_io_PF_Valid),
    .io_NoDPE(PathFinder_10_io_NoDPE),
    .io_DataValid(PathFinder_10_io_DataValid)
  );
  PathFinder PathFinder_11 ( // @[FlexDPU.scala 77:41]
    .clock(PathFinder_11_clock),
    .reset(PathFinder_11_reset),
    .io_Stationary_matrix_0_0(PathFinder_11_io_Stationary_matrix_0_0),
    .io_Stationary_matrix_0_1(PathFinder_11_io_Stationary_matrix_0_1),
    .io_Stationary_matrix_0_2(PathFinder_11_io_Stationary_matrix_0_2),
    .io_Stationary_matrix_0_3(PathFinder_11_io_Stationary_matrix_0_3),
    .io_Stationary_matrix_0_4(PathFinder_11_io_Stationary_matrix_0_4),
    .io_Stationary_matrix_0_5(PathFinder_11_io_Stationary_matrix_0_5),
    .io_Stationary_matrix_0_6(PathFinder_11_io_Stationary_matrix_0_6),
    .io_Stationary_matrix_0_7(PathFinder_11_io_Stationary_matrix_0_7),
    .io_Stationary_matrix_1_0(PathFinder_11_io_Stationary_matrix_1_0),
    .io_Stationary_matrix_1_1(PathFinder_11_io_Stationary_matrix_1_1),
    .io_Stationary_matrix_1_2(PathFinder_11_io_Stationary_matrix_1_2),
    .io_Stationary_matrix_1_3(PathFinder_11_io_Stationary_matrix_1_3),
    .io_Stationary_matrix_1_4(PathFinder_11_io_Stationary_matrix_1_4),
    .io_Stationary_matrix_1_5(PathFinder_11_io_Stationary_matrix_1_5),
    .io_Stationary_matrix_1_6(PathFinder_11_io_Stationary_matrix_1_6),
    .io_Stationary_matrix_1_7(PathFinder_11_io_Stationary_matrix_1_7),
    .io_Stationary_matrix_2_0(PathFinder_11_io_Stationary_matrix_2_0),
    .io_Stationary_matrix_2_1(PathFinder_11_io_Stationary_matrix_2_1),
    .io_Stationary_matrix_2_2(PathFinder_11_io_Stationary_matrix_2_2),
    .io_Stationary_matrix_2_3(PathFinder_11_io_Stationary_matrix_2_3),
    .io_Stationary_matrix_2_4(PathFinder_11_io_Stationary_matrix_2_4),
    .io_Stationary_matrix_2_5(PathFinder_11_io_Stationary_matrix_2_5),
    .io_Stationary_matrix_2_6(PathFinder_11_io_Stationary_matrix_2_6),
    .io_Stationary_matrix_2_7(PathFinder_11_io_Stationary_matrix_2_7),
    .io_Stationary_matrix_3_0(PathFinder_11_io_Stationary_matrix_3_0),
    .io_Stationary_matrix_3_1(PathFinder_11_io_Stationary_matrix_3_1),
    .io_Stationary_matrix_3_2(PathFinder_11_io_Stationary_matrix_3_2),
    .io_Stationary_matrix_3_3(PathFinder_11_io_Stationary_matrix_3_3),
    .io_Stationary_matrix_3_4(PathFinder_11_io_Stationary_matrix_3_4),
    .io_Stationary_matrix_3_5(PathFinder_11_io_Stationary_matrix_3_5),
    .io_Stationary_matrix_3_6(PathFinder_11_io_Stationary_matrix_3_6),
    .io_Stationary_matrix_3_7(PathFinder_11_io_Stationary_matrix_3_7),
    .io_Stationary_matrix_4_0(PathFinder_11_io_Stationary_matrix_4_0),
    .io_Stationary_matrix_4_1(PathFinder_11_io_Stationary_matrix_4_1),
    .io_Stationary_matrix_4_2(PathFinder_11_io_Stationary_matrix_4_2),
    .io_Stationary_matrix_4_3(PathFinder_11_io_Stationary_matrix_4_3),
    .io_Stationary_matrix_4_4(PathFinder_11_io_Stationary_matrix_4_4),
    .io_Stationary_matrix_4_5(PathFinder_11_io_Stationary_matrix_4_5),
    .io_Stationary_matrix_4_6(PathFinder_11_io_Stationary_matrix_4_6),
    .io_Stationary_matrix_4_7(PathFinder_11_io_Stationary_matrix_4_7),
    .io_Stationary_matrix_5_0(PathFinder_11_io_Stationary_matrix_5_0),
    .io_Stationary_matrix_5_1(PathFinder_11_io_Stationary_matrix_5_1),
    .io_Stationary_matrix_5_2(PathFinder_11_io_Stationary_matrix_5_2),
    .io_Stationary_matrix_5_3(PathFinder_11_io_Stationary_matrix_5_3),
    .io_Stationary_matrix_5_4(PathFinder_11_io_Stationary_matrix_5_4),
    .io_Stationary_matrix_5_5(PathFinder_11_io_Stationary_matrix_5_5),
    .io_Stationary_matrix_5_6(PathFinder_11_io_Stationary_matrix_5_6),
    .io_Stationary_matrix_5_7(PathFinder_11_io_Stationary_matrix_5_7),
    .io_Stationary_matrix_6_0(PathFinder_11_io_Stationary_matrix_6_0),
    .io_Stationary_matrix_6_1(PathFinder_11_io_Stationary_matrix_6_1),
    .io_Stationary_matrix_6_2(PathFinder_11_io_Stationary_matrix_6_2),
    .io_Stationary_matrix_6_3(PathFinder_11_io_Stationary_matrix_6_3),
    .io_Stationary_matrix_6_4(PathFinder_11_io_Stationary_matrix_6_4),
    .io_Stationary_matrix_6_5(PathFinder_11_io_Stationary_matrix_6_5),
    .io_Stationary_matrix_6_6(PathFinder_11_io_Stationary_matrix_6_6),
    .io_Stationary_matrix_6_7(PathFinder_11_io_Stationary_matrix_6_7),
    .io_Stationary_matrix_7_0(PathFinder_11_io_Stationary_matrix_7_0),
    .io_Stationary_matrix_7_1(PathFinder_11_io_Stationary_matrix_7_1),
    .io_Stationary_matrix_7_2(PathFinder_11_io_Stationary_matrix_7_2),
    .io_Stationary_matrix_7_3(PathFinder_11_io_Stationary_matrix_7_3),
    .io_Stationary_matrix_7_4(PathFinder_11_io_Stationary_matrix_7_4),
    .io_Stationary_matrix_7_5(PathFinder_11_io_Stationary_matrix_7_5),
    .io_Stationary_matrix_7_6(PathFinder_11_io_Stationary_matrix_7_6),
    .io_Stationary_matrix_7_7(PathFinder_11_io_Stationary_matrix_7_7),
    .io_Streaming_matrix_0(PathFinder_11_io_Streaming_matrix_0),
    .io_Streaming_matrix_1(PathFinder_11_io_Streaming_matrix_1),
    .io_Streaming_matrix_2(PathFinder_11_io_Streaming_matrix_2),
    .io_Streaming_matrix_3(PathFinder_11_io_Streaming_matrix_3),
    .io_Streaming_matrix_4(PathFinder_11_io_Streaming_matrix_4),
    .io_Streaming_matrix_5(PathFinder_11_io_Streaming_matrix_5),
    .io_Streaming_matrix_6(PathFinder_11_io_Streaming_matrix_6),
    .io_Streaming_matrix_7(PathFinder_11_io_Streaming_matrix_7),
    .io_i_mux_bus_0(PathFinder_11_io_i_mux_bus_0),
    .io_i_mux_bus_1(PathFinder_11_io_i_mux_bus_1),
    .io_i_mux_bus_2(PathFinder_11_io_i_mux_bus_2),
    .io_i_mux_bus_3(PathFinder_11_io_i_mux_bus_3),
    .io_Source_0(PathFinder_11_io_Source_0),
    .io_Source_1(PathFinder_11_io_Source_1),
    .io_Source_2(PathFinder_11_io_Source_2),
    .io_Source_3(PathFinder_11_io_Source_3),
    .io_PF_Valid(PathFinder_11_io_PF_Valid),
    .io_NoDPE(PathFinder_11_io_NoDPE),
    .io_DataValid(PathFinder_11_io_DataValid)
  );
  PathFinder PathFinder_12 ( // @[FlexDPU.scala 77:41]
    .clock(PathFinder_12_clock),
    .reset(PathFinder_12_reset),
    .io_Stationary_matrix_0_0(PathFinder_12_io_Stationary_matrix_0_0),
    .io_Stationary_matrix_0_1(PathFinder_12_io_Stationary_matrix_0_1),
    .io_Stationary_matrix_0_2(PathFinder_12_io_Stationary_matrix_0_2),
    .io_Stationary_matrix_0_3(PathFinder_12_io_Stationary_matrix_0_3),
    .io_Stationary_matrix_0_4(PathFinder_12_io_Stationary_matrix_0_4),
    .io_Stationary_matrix_0_5(PathFinder_12_io_Stationary_matrix_0_5),
    .io_Stationary_matrix_0_6(PathFinder_12_io_Stationary_matrix_0_6),
    .io_Stationary_matrix_0_7(PathFinder_12_io_Stationary_matrix_0_7),
    .io_Stationary_matrix_1_0(PathFinder_12_io_Stationary_matrix_1_0),
    .io_Stationary_matrix_1_1(PathFinder_12_io_Stationary_matrix_1_1),
    .io_Stationary_matrix_1_2(PathFinder_12_io_Stationary_matrix_1_2),
    .io_Stationary_matrix_1_3(PathFinder_12_io_Stationary_matrix_1_3),
    .io_Stationary_matrix_1_4(PathFinder_12_io_Stationary_matrix_1_4),
    .io_Stationary_matrix_1_5(PathFinder_12_io_Stationary_matrix_1_5),
    .io_Stationary_matrix_1_6(PathFinder_12_io_Stationary_matrix_1_6),
    .io_Stationary_matrix_1_7(PathFinder_12_io_Stationary_matrix_1_7),
    .io_Stationary_matrix_2_0(PathFinder_12_io_Stationary_matrix_2_0),
    .io_Stationary_matrix_2_1(PathFinder_12_io_Stationary_matrix_2_1),
    .io_Stationary_matrix_2_2(PathFinder_12_io_Stationary_matrix_2_2),
    .io_Stationary_matrix_2_3(PathFinder_12_io_Stationary_matrix_2_3),
    .io_Stationary_matrix_2_4(PathFinder_12_io_Stationary_matrix_2_4),
    .io_Stationary_matrix_2_5(PathFinder_12_io_Stationary_matrix_2_5),
    .io_Stationary_matrix_2_6(PathFinder_12_io_Stationary_matrix_2_6),
    .io_Stationary_matrix_2_7(PathFinder_12_io_Stationary_matrix_2_7),
    .io_Stationary_matrix_3_0(PathFinder_12_io_Stationary_matrix_3_0),
    .io_Stationary_matrix_3_1(PathFinder_12_io_Stationary_matrix_3_1),
    .io_Stationary_matrix_3_2(PathFinder_12_io_Stationary_matrix_3_2),
    .io_Stationary_matrix_3_3(PathFinder_12_io_Stationary_matrix_3_3),
    .io_Stationary_matrix_3_4(PathFinder_12_io_Stationary_matrix_3_4),
    .io_Stationary_matrix_3_5(PathFinder_12_io_Stationary_matrix_3_5),
    .io_Stationary_matrix_3_6(PathFinder_12_io_Stationary_matrix_3_6),
    .io_Stationary_matrix_3_7(PathFinder_12_io_Stationary_matrix_3_7),
    .io_Stationary_matrix_4_0(PathFinder_12_io_Stationary_matrix_4_0),
    .io_Stationary_matrix_4_1(PathFinder_12_io_Stationary_matrix_4_1),
    .io_Stationary_matrix_4_2(PathFinder_12_io_Stationary_matrix_4_2),
    .io_Stationary_matrix_4_3(PathFinder_12_io_Stationary_matrix_4_3),
    .io_Stationary_matrix_4_4(PathFinder_12_io_Stationary_matrix_4_4),
    .io_Stationary_matrix_4_5(PathFinder_12_io_Stationary_matrix_4_5),
    .io_Stationary_matrix_4_6(PathFinder_12_io_Stationary_matrix_4_6),
    .io_Stationary_matrix_4_7(PathFinder_12_io_Stationary_matrix_4_7),
    .io_Stationary_matrix_5_0(PathFinder_12_io_Stationary_matrix_5_0),
    .io_Stationary_matrix_5_1(PathFinder_12_io_Stationary_matrix_5_1),
    .io_Stationary_matrix_5_2(PathFinder_12_io_Stationary_matrix_5_2),
    .io_Stationary_matrix_5_3(PathFinder_12_io_Stationary_matrix_5_3),
    .io_Stationary_matrix_5_4(PathFinder_12_io_Stationary_matrix_5_4),
    .io_Stationary_matrix_5_5(PathFinder_12_io_Stationary_matrix_5_5),
    .io_Stationary_matrix_5_6(PathFinder_12_io_Stationary_matrix_5_6),
    .io_Stationary_matrix_5_7(PathFinder_12_io_Stationary_matrix_5_7),
    .io_Stationary_matrix_6_0(PathFinder_12_io_Stationary_matrix_6_0),
    .io_Stationary_matrix_6_1(PathFinder_12_io_Stationary_matrix_6_1),
    .io_Stationary_matrix_6_2(PathFinder_12_io_Stationary_matrix_6_2),
    .io_Stationary_matrix_6_3(PathFinder_12_io_Stationary_matrix_6_3),
    .io_Stationary_matrix_6_4(PathFinder_12_io_Stationary_matrix_6_4),
    .io_Stationary_matrix_6_5(PathFinder_12_io_Stationary_matrix_6_5),
    .io_Stationary_matrix_6_6(PathFinder_12_io_Stationary_matrix_6_6),
    .io_Stationary_matrix_6_7(PathFinder_12_io_Stationary_matrix_6_7),
    .io_Stationary_matrix_7_0(PathFinder_12_io_Stationary_matrix_7_0),
    .io_Stationary_matrix_7_1(PathFinder_12_io_Stationary_matrix_7_1),
    .io_Stationary_matrix_7_2(PathFinder_12_io_Stationary_matrix_7_2),
    .io_Stationary_matrix_7_3(PathFinder_12_io_Stationary_matrix_7_3),
    .io_Stationary_matrix_7_4(PathFinder_12_io_Stationary_matrix_7_4),
    .io_Stationary_matrix_7_5(PathFinder_12_io_Stationary_matrix_7_5),
    .io_Stationary_matrix_7_6(PathFinder_12_io_Stationary_matrix_7_6),
    .io_Stationary_matrix_7_7(PathFinder_12_io_Stationary_matrix_7_7),
    .io_Streaming_matrix_0(PathFinder_12_io_Streaming_matrix_0),
    .io_Streaming_matrix_1(PathFinder_12_io_Streaming_matrix_1),
    .io_Streaming_matrix_2(PathFinder_12_io_Streaming_matrix_2),
    .io_Streaming_matrix_3(PathFinder_12_io_Streaming_matrix_3),
    .io_Streaming_matrix_4(PathFinder_12_io_Streaming_matrix_4),
    .io_Streaming_matrix_5(PathFinder_12_io_Streaming_matrix_5),
    .io_Streaming_matrix_6(PathFinder_12_io_Streaming_matrix_6),
    .io_Streaming_matrix_7(PathFinder_12_io_Streaming_matrix_7),
    .io_i_mux_bus_0(PathFinder_12_io_i_mux_bus_0),
    .io_i_mux_bus_1(PathFinder_12_io_i_mux_bus_1),
    .io_i_mux_bus_2(PathFinder_12_io_i_mux_bus_2),
    .io_i_mux_bus_3(PathFinder_12_io_i_mux_bus_3),
    .io_Source_0(PathFinder_12_io_Source_0),
    .io_Source_1(PathFinder_12_io_Source_1),
    .io_Source_2(PathFinder_12_io_Source_2),
    .io_Source_3(PathFinder_12_io_Source_3),
    .io_PF_Valid(PathFinder_12_io_PF_Valid),
    .io_NoDPE(PathFinder_12_io_NoDPE),
    .io_DataValid(PathFinder_12_io_DataValid)
  );
  PathFinder PathFinder_13 ( // @[FlexDPU.scala 77:41]
    .clock(PathFinder_13_clock),
    .reset(PathFinder_13_reset),
    .io_Stationary_matrix_0_0(PathFinder_13_io_Stationary_matrix_0_0),
    .io_Stationary_matrix_0_1(PathFinder_13_io_Stationary_matrix_0_1),
    .io_Stationary_matrix_0_2(PathFinder_13_io_Stationary_matrix_0_2),
    .io_Stationary_matrix_0_3(PathFinder_13_io_Stationary_matrix_0_3),
    .io_Stationary_matrix_0_4(PathFinder_13_io_Stationary_matrix_0_4),
    .io_Stationary_matrix_0_5(PathFinder_13_io_Stationary_matrix_0_5),
    .io_Stationary_matrix_0_6(PathFinder_13_io_Stationary_matrix_0_6),
    .io_Stationary_matrix_0_7(PathFinder_13_io_Stationary_matrix_0_7),
    .io_Stationary_matrix_1_0(PathFinder_13_io_Stationary_matrix_1_0),
    .io_Stationary_matrix_1_1(PathFinder_13_io_Stationary_matrix_1_1),
    .io_Stationary_matrix_1_2(PathFinder_13_io_Stationary_matrix_1_2),
    .io_Stationary_matrix_1_3(PathFinder_13_io_Stationary_matrix_1_3),
    .io_Stationary_matrix_1_4(PathFinder_13_io_Stationary_matrix_1_4),
    .io_Stationary_matrix_1_5(PathFinder_13_io_Stationary_matrix_1_5),
    .io_Stationary_matrix_1_6(PathFinder_13_io_Stationary_matrix_1_6),
    .io_Stationary_matrix_1_7(PathFinder_13_io_Stationary_matrix_1_7),
    .io_Stationary_matrix_2_0(PathFinder_13_io_Stationary_matrix_2_0),
    .io_Stationary_matrix_2_1(PathFinder_13_io_Stationary_matrix_2_1),
    .io_Stationary_matrix_2_2(PathFinder_13_io_Stationary_matrix_2_2),
    .io_Stationary_matrix_2_3(PathFinder_13_io_Stationary_matrix_2_3),
    .io_Stationary_matrix_2_4(PathFinder_13_io_Stationary_matrix_2_4),
    .io_Stationary_matrix_2_5(PathFinder_13_io_Stationary_matrix_2_5),
    .io_Stationary_matrix_2_6(PathFinder_13_io_Stationary_matrix_2_6),
    .io_Stationary_matrix_2_7(PathFinder_13_io_Stationary_matrix_2_7),
    .io_Stationary_matrix_3_0(PathFinder_13_io_Stationary_matrix_3_0),
    .io_Stationary_matrix_3_1(PathFinder_13_io_Stationary_matrix_3_1),
    .io_Stationary_matrix_3_2(PathFinder_13_io_Stationary_matrix_3_2),
    .io_Stationary_matrix_3_3(PathFinder_13_io_Stationary_matrix_3_3),
    .io_Stationary_matrix_3_4(PathFinder_13_io_Stationary_matrix_3_4),
    .io_Stationary_matrix_3_5(PathFinder_13_io_Stationary_matrix_3_5),
    .io_Stationary_matrix_3_6(PathFinder_13_io_Stationary_matrix_3_6),
    .io_Stationary_matrix_3_7(PathFinder_13_io_Stationary_matrix_3_7),
    .io_Stationary_matrix_4_0(PathFinder_13_io_Stationary_matrix_4_0),
    .io_Stationary_matrix_4_1(PathFinder_13_io_Stationary_matrix_4_1),
    .io_Stationary_matrix_4_2(PathFinder_13_io_Stationary_matrix_4_2),
    .io_Stationary_matrix_4_3(PathFinder_13_io_Stationary_matrix_4_3),
    .io_Stationary_matrix_4_4(PathFinder_13_io_Stationary_matrix_4_4),
    .io_Stationary_matrix_4_5(PathFinder_13_io_Stationary_matrix_4_5),
    .io_Stationary_matrix_4_6(PathFinder_13_io_Stationary_matrix_4_6),
    .io_Stationary_matrix_4_7(PathFinder_13_io_Stationary_matrix_4_7),
    .io_Stationary_matrix_5_0(PathFinder_13_io_Stationary_matrix_5_0),
    .io_Stationary_matrix_5_1(PathFinder_13_io_Stationary_matrix_5_1),
    .io_Stationary_matrix_5_2(PathFinder_13_io_Stationary_matrix_5_2),
    .io_Stationary_matrix_5_3(PathFinder_13_io_Stationary_matrix_5_3),
    .io_Stationary_matrix_5_4(PathFinder_13_io_Stationary_matrix_5_4),
    .io_Stationary_matrix_5_5(PathFinder_13_io_Stationary_matrix_5_5),
    .io_Stationary_matrix_5_6(PathFinder_13_io_Stationary_matrix_5_6),
    .io_Stationary_matrix_5_7(PathFinder_13_io_Stationary_matrix_5_7),
    .io_Stationary_matrix_6_0(PathFinder_13_io_Stationary_matrix_6_0),
    .io_Stationary_matrix_6_1(PathFinder_13_io_Stationary_matrix_6_1),
    .io_Stationary_matrix_6_2(PathFinder_13_io_Stationary_matrix_6_2),
    .io_Stationary_matrix_6_3(PathFinder_13_io_Stationary_matrix_6_3),
    .io_Stationary_matrix_6_4(PathFinder_13_io_Stationary_matrix_6_4),
    .io_Stationary_matrix_6_5(PathFinder_13_io_Stationary_matrix_6_5),
    .io_Stationary_matrix_6_6(PathFinder_13_io_Stationary_matrix_6_6),
    .io_Stationary_matrix_6_7(PathFinder_13_io_Stationary_matrix_6_7),
    .io_Stationary_matrix_7_0(PathFinder_13_io_Stationary_matrix_7_0),
    .io_Stationary_matrix_7_1(PathFinder_13_io_Stationary_matrix_7_1),
    .io_Stationary_matrix_7_2(PathFinder_13_io_Stationary_matrix_7_2),
    .io_Stationary_matrix_7_3(PathFinder_13_io_Stationary_matrix_7_3),
    .io_Stationary_matrix_7_4(PathFinder_13_io_Stationary_matrix_7_4),
    .io_Stationary_matrix_7_5(PathFinder_13_io_Stationary_matrix_7_5),
    .io_Stationary_matrix_7_6(PathFinder_13_io_Stationary_matrix_7_6),
    .io_Stationary_matrix_7_7(PathFinder_13_io_Stationary_matrix_7_7),
    .io_Streaming_matrix_0(PathFinder_13_io_Streaming_matrix_0),
    .io_Streaming_matrix_1(PathFinder_13_io_Streaming_matrix_1),
    .io_Streaming_matrix_2(PathFinder_13_io_Streaming_matrix_2),
    .io_Streaming_matrix_3(PathFinder_13_io_Streaming_matrix_3),
    .io_Streaming_matrix_4(PathFinder_13_io_Streaming_matrix_4),
    .io_Streaming_matrix_5(PathFinder_13_io_Streaming_matrix_5),
    .io_Streaming_matrix_6(PathFinder_13_io_Streaming_matrix_6),
    .io_Streaming_matrix_7(PathFinder_13_io_Streaming_matrix_7),
    .io_i_mux_bus_0(PathFinder_13_io_i_mux_bus_0),
    .io_i_mux_bus_1(PathFinder_13_io_i_mux_bus_1),
    .io_i_mux_bus_2(PathFinder_13_io_i_mux_bus_2),
    .io_i_mux_bus_3(PathFinder_13_io_i_mux_bus_3),
    .io_Source_0(PathFinder_13_io_Source_0),
    .io_Source_1(PathFinder_13_io_Source_1),
    .io_Source_2(PathFinder_13_io_Source_2),
    .io_Source_3(PathFinder_13_io_Source_3),
    .io_PF_Valid(PathFinder_13_io_PF_Valid),
    .io_NoDPE(PathFinder_13_io_NoDPE),
    .io_DataValid(PathFinder_13_io_DataValid)
  );
  PathFinder PathFinder_14 ( // @[FlexDPU.scala 77:41]
    .clock(PathFinder_14_clock),
    .reset(PathFinder_14_reset),
    .io_Stationary_matrix_0_0(PathFinder_14_io_Stationary_matrix_0_0),
    .io_Stationary_matrix_0_1(PathFinder_14_io_Stationary_matrix_0_1),
    .io_Stationary_matrix_0_2(PathFinder_14_io_Stationary_matrix_0_2),
    .io_Stationary_matrix_0_3(PathFinder_14_io_Stationary_matrix_0_3),
    .io_Stationary_matrix_0_4(PathFinder_14_io_Stationary_matrix_0_4),
    .io_Stationary_matrix_0_5(PathFinder_14_io_Stationary_matrix_0_5),
    .io_Stationary_matrix_0_6(PathFinder_14_io_Stationary_matrix_0_6),
    .io_Stationary_matrix_0_7(PathFinder_14_io_Stationary_matrix_0_7),
    .io_Stationary_matrix_1_0(PathFinder_14_io_Stationary_matrix_1_0),
    .io_Stationary_matrix_1_1(PathFinder_14_io_Stationary_matrix_1_1),
    .io_Stationary_matrix_1_2(PathFinder_14_io_Stationary_matrix_1_2),
    .io_Stationary_matrix_1_3(PathFinder_14_io_Stationary_matrix_1_3),
    .io_Stationary_matrix_1_4(PathFinder_14_io_Stationary_matrix_1_4),
    .io_Stationary_matrix_1_5(PathFinder_14_io_Stationary_matrix_1_5),
    .io_Stationary_matrix_1_6(PathFinder_14_io_Stationary_matrix_1_6),
    .io_Stationary_matrix_1_7(PathFinder_14_io_Stationary_matrix_1_7),
    .io_Stationary_matrix_2_0(PathFinder_14_io_Stationary_matrix_2_0),
    .io_Stationary_matrix_2_1(PathFinder_14_io_Stationary_matrix_2_1),
    .io_Stationary_matrix_2_2(PathFinder_14_io_Stationary_matrix_2_2),
    .io_Stationary_matrix_2_3(PathFinder_14_io_Stationary_matrix_2_3),
    .io_Stationary_matrix_2_4(PathFinder_14_io_Stationary_matrix_2_4),
    .io_Stationary_matrix_2_5(PathFinder_14_io_Stationary_matrix_2_5),
    .io_Stationary_matrix_2_6(PathFinder_14_io_Stationary_matrix_2_6),
    .io_Stationary_matrix_2_7(PathFinder_14_io_Stationary_matrix_2_7),
    .io_Stationary_matrix_3_0(PathFinder_14_io_Stationary_matrix_3_0),
    .io_Stationary_matrix_3_1(PathFinder_14_io_Stationary_matrix_3_1),
    .io_Stationary_matrix_3_2(PathFinder_14_io_Stationary_matrix_3_2),
    .io_Stationary_matrix_3_3(PathFinder_14_io_Stationary_matrix_3_3),
    .io_Stationary_matrix_3_4(PathFinder_14_io_Stationary_matrix_3_4),
    .io_Stationary_matrix_3_5(PathFinder_14_io_Stationary_matrix_3_5),
    .io_Stationary_matrix_3_6(PathFinder_14_io_Stationary_matrix_3_6),
    .io_Stationary_matrix_3_7(PathFinder_14_io_Stationary_matrix_3_7),
    .io_Stationary_matrix_4_0(PathFinder_14_io_Stationary_matrix_4_0),
    .io_Stationary_matrix_4_1(PathFinder_14_io_Stationary_matrix_4_1),
    .io_Stationary_matrix_4_2(PathFinder_14_io_Stationary_matrix_4_2),
    .io_Stationary_matrix_4_3(PathFinder_14_io_Stationary_matrix_4_3),
    .io_Stationary_matrix_4_4(PathFinder_14_io_Stationary_matrix_4_4),
    .io_Stationary_matrix_4_5(PathFinder_14_io_Stationary_matrix_4_5),
    .io_Stationary_matrix_4_6(PathFinder_14_io_Stationary_matrix_4_6),
    .io_Stationary_matrix_4_7(PathFinder_14_io_Stationary_matrix_4_7),
    .io_Stationary_matrix_5_0(PathFinder_14_io_Stationary_matrix_5_0),
    .io_Stationary_matrix_5_1(PathFinder_14_io_Stationary_matrix_5_1),
    .io_Stationary_matrix_5_2(PathFinder_14_io_Stationary_matrix_5_2),
    .io_Stationary_matrix_5_3(PathFinder_14_io_Stationary_matrix_5_3),
    .io_Stationary_matrix_5_4(PathFinder_14_io_Stationary_matrix_5_4),
    .io_Stationary_matrix_5_5(PathFinder_14_io_Stationary_matrix_5_5),
    .io_Stationary_matrix_5_6(PathFinder_14_io_Stationary_matrix_5_6),
    .io_Stationary_matrix_5_7(PathFinder_14_io_Stationary_matrix_5_7),
    .io_Stationary_matrix_6_0(PathFinder_14_io_Stationary_matrix_6_0),
    .io_Stationary_matrix_6_1(PathFinder_14_io_Stationary_matrix_6_1),
    .io_Stationary_matrix_6_2(PathFinder_14_io_Stationary_matrix_6_2),
    .io_Stationary_matrix_6_3(PathFinder_14_io_Stationary_matrix_6_3),
    .io_Stationary_matrix_6_4(PathFinder_14_io_Stationary_matrix_6_4),
    .io_Stationary_matrix_6_5(PathFinder_14_io_Stationary_matrix_6_5),
    .io_Stationary_matrix_6_6(PathFinder_14_io_Stationary_matrix_6_6),
    .io_Stationary_matrix_6_7(PathFinder_14_io_Stationary_matrix_6_7),
    .io_Stationary_matrix_7_0(PathFinder_14_io_Stationary_matrix_7_0),
    .io_Stationary_matrix_7_1(PathFinder_14_io_Stationary_matrix_7_1),
    .io_Stationary_matrix_7_2(PathFinder_14_io_Stationary_matrix_7_2),
    .io_Stationary_matrix_7_3(PathFinder_14_io_Stationary_matrix_7_3),
    .io_Stationary_matrix_7_4(PathFinder_14_io_Stationary_matrix_7_4),
    .io_Stationary_matrix_7_5(PathFinder_14_io_Stationary_matrix_7_5),
    .io_Stationary_matrix_7_6(PathFinder_14_io_Stationary_matrix_7_6),
    .io_Stationary_matrix_7_7(PathFinder_14_io_Stationary_matrix_7_7),
    .io_Streaming_matrix_0(PathFinder_14_io_Streaming_matrix_0),
    .io_Streaming_matrix_1(PathFinder_14_io_Streaming_matrix_1),
    .io_Streaming_matrix_2(PathFinder_14_io_Streaming_matrix_2),
    .io_Streaming_matrix_3(PathFinder_14_io_Streaming_matrix_3),
    .io_Streaming_matrix_4(PathFinder_14_io_Streaming_matrix_4),
    .io_Streaming_matrix_5(PathFinder_14_io_Streaming_matrix_5),
    .io_Streaming_matrix_6(PathFinder_14_io_Streaming_matrix_6),
    .io_Streaming_matrix_7(PathFinder_14_io_Streaming_matrix_7),
    .io_i_mux_bus_0(PathFinder_14_io_i_mux_bus_0),
    .io_i_mux_bus_1(PathFinder_14_io_i_mux_bus_1),
    .io_i_mux_bus_2(PathFinder_14_io_i_mux_bus_2),
    .io_i_mux_bus_3(PathFinder_14_io_i_mux_bus_3),
    .io_Source_0(PathFinder_14_io_Source_0),
    .io_Source_1(PathFinder_14_io_Source_1),
    .io_Source_2(PathFinder_14_io_Source_2),
    .io_Source_3(PathFinder_14_io_Source_3),
    .io_PF_Valid(PathFinder_14_io_PF_Valid),
    .io_NoDPE(PathFinder_14_io_NoDPE),
    .io_DataValid(PathFinder_14_io_DataValid)
  );
  PathFinder PathFinder_15 ( // @[FlexDPU.scala 77:41]
    .clock(PathFinder_15_clock),
    .reset(PathFinder_15_reset),
    .io_Stationary_matrix_0_0(PathFinder_15_io_Stationary_matrix_0_0),
    .io_Stationary_matrix_0_1(PathFinder_15_io_Stationary_matrix_0_1),
    .io_Stationary_matrix_0_2(PathFinder_15_io_Stationary_matrix_0_2),
    .io_Stationary_matrix_0_3(PathFinder_15_io_Stationary_matrix_0_3),
    .io_Stationary_matrix_0_4(PathFinder_15_io_Stationary_matrix_0_4),
    .io_Stationary_matrix_0_5(PathFinder_15_io_Stationary_matrix_0_5),
    .io_Stationary_matrix_0_6(PathFinder_15_io_Stationary_matrix_0_6),
    .io_Stationary_matrix_0_7(PathFinder_15_io_Stationary_matrix_0_7),
    .io_Stationary_matrix_1_0(PathFinder_15_io_Stationary_matrix_1_0),
    .io_Stationary_matrix_1_1(PathFinder_15_io_Stationary_matrix_1_1),
    .io_Stationary_matrix_1_2(PathFinder_15_io_Stationary_matrix_1_2),
    .io_Stationary_matrix_1_3(PathFinder_15_io_Stationary_matrix_1_3),
    .io_Stationary_matrix_1_4(PathFinder_15_io_Stationary_matrix_1_4),
    .io_Stationary_matrix_1_5(PathFinder_15_io_Stationary_matrix_1_5),
    .io_Stationary_matrix_1_6(PathFinder_15_io_Stationary_matrix_1_6),
    .io_Stationary_matrix_1_7(PathFinder_15_io_Stationary_matrix_1_7),
    .io_Stationary_matrix_2_0(PathFinder_15_io_Stationary_matrix_2_0),
    .io_Stationary_matrix_2_1(PathFinder_15_io_Stationary_matrix_2_1),
    .io_Stationary_matrix_2_2(PathFinder_15_io_Stationary_matrix_2_2),
    .io_Stationary_matrix_2_3(PathFinder_15_io_Stationary_matrix_2_3),
    .io_Stationary_matrix_2_4(PathFinder_15_io_Stationary_matrix_2_4),
    .io_Stationary_matrix_2_5(PathFinder_15_io_Stationary_matrix_2_5),
    .io_Stationary_matrix_2_6(PathFinder_15_io_Stationary_matrix_2_6),
    .io_Stationary_matrix_2_7(PathFinder_15_io_Stationary_matrix_2_7),
    .io_Stationary_matrix_3_0(PathFinder_15_io_Stationary_matrix_3_0),
    .io_Stationary_matrix_3_1(PathFinder_15_io_Stationary_matrix_3_1),
    .io_Stationary_matrix_3_2(PathFinder_15_io_Stationary_matrix_3_2),
    .io_Stationary_matrix_3_3(PathFinder_15_io_Stationary_matrix_3_3),
    .io_Stationary_matrix_3_4(PathFinder_15_io_Stationary_matrix_3_4),
    .io_Stationary_matrix_3_5(PathFinder_15_io_Stationary_matrix_3_5),
    .io_Stationary_matrix_3_6(PathFinder_15_io_Stationary_matrix_3_6),
    .io_Stationary_matrix_3_7(PathFinder_15_io_Stationary_matrix_3_7),
    .io_Stationary_matrix_4_0(PathFinder_15_io_Stationary_matrix_4_0),
    .io_Stationary_matrix_4_1(PathFinder_15_io_Stationary_matrix_4_1),
    .io_Stationary_matrix_4_2(PathFinder_15_io_Stationary_matrix_4_2),
    .io_Stationary_matrix_4_3(PathFinder_15_io_Stationary_matrix_4_3),
    .io_Stationary_matrix_4_4(PathFinder_15_io_Stationary_matrix_4_4),
    .io_Stationary_matrix_4_5(PathFinder_15_io_Stationary_matrix_4_5),
    .io_Stationary_matrix_4_6(PathFinder_15_io_Stationary_matrix_4_6),
    .io_Stationary_matrix_4_7(PathFinder_15_io_Stationary_matrix_4_7),
    .io_Stationary_matrix_5_0(PathFinder_15_io_Stationary_matrix_5_0),
    .io_Stationary_matrix_5_1(PathFinder_15_io_Stationary_matrix_5_1),
    .io_Stationary_matrix_5_2(PathFinder_15_io_Stationary_matrix_5_2),
    .io_Stationary_matrix_5_3(PathFinder_15_io_Stationary_matrix_5_3),
    .io_Stationary_matrix_5_4(PathFinder_15_io_Stationary_matrix_5_4),
    .io_Stationary_matrix_5_5(PathFinder_15_io_Stationary_matrix_5_5),
    .io_Stationary_matrix_5_6(PathFinder_15_io_Stationary_matrix_5_6),
    .io_Stationary_matrix_5_7(PathFinder_15_io_Stationary_matrix_5_7),
    .io_Stationary_matrix_6_0(PathFinder_15_io_Stationary_matrix_6_0),
    .io_Stationary_matrix_6_1(PathFinder_15_io_Stationary_matrix_6_1),
    .io_Stationary_matrix_6_2(PathFinder_15_io_Stationary_matrix_6_2),
    .io_Stationary_matrix_6_3(PathFinder_15_io_Stationary_matrix_6_3),
    .io_Stationary_matrix_6_4(PathFinder_15_io_Stationary_matrix_6_4),
    .io_Stationary_matrix_6_5(PathFinder_15_io_Stationary_matrix_6_5),
    .io_Stationary_matrix_6_6(PathFinder_15_io_Stationary_matrix_6_6),
    .io_Stationary_matrix_6_7(PathFinder_15_io_Stationary_matrix_6_7),
    .io_Stationary_matrix_7_0(PathFinder_15_io_Stationary_matrix_7_0),
    .io_Stationary_matrix_7_1(PathFinder_15_io_Stationary_matrix_7_1),
    .io_Stationary_matrix_7_2(PathFinder_15_io_Stationary_matrix_7_2),
    .io_Stationary_matrix_7_3(PathFinder_15_io_Stationary_matrix_7_3),
    .io_Stationary_matrix_7_4(PathFinder_15_io_Stationary_matrix_7_4),
    .io_Stationary_matrix_7_5(PathFinder_15_io_Stationary_matrix_7_5),
    .io_Stationary_matrix_7_6(PathFinder_15_io_Stationary_matrix_7_6),
    .io_Stationary_matrix_7_7(PathFinder_15_io_Stationary_matrix_7_7),
    .io_Streaming_matrix_0(PathFinder_15_io_Streaming_matrix_0),
    .io_Streaming_matrix_1(PathFinder_15_io_Streaming_matrix_1),
    .io_Streaming_matrix_2(PathFinder_15_io_Streaming_matrix_2),
    .io_Streaming_matrix_3(PathFinder_15_io_Streaming_matrix_3),
    .io_Streaming_matrix_4(PathFinder_15_io_Streaming_matrix_4),
    .io_Streaming_matrix_5(PathFinder_15_io_Streaming_matrix_5),
    .io_Streaming_matrix_6(PathFinder_15_io_Streaming_matrix_6),
    .io_Streaming_matrix_7(PathFinder_15_io_Streaming_matrix_7),
    .io_i_mux_bus_0(PathFinder_15_io_i_mux_bus_0),
    .io_i_mux_bus_1(PathFinder_15_io_i_mux_bus_1),
    .io_i_mux_bus_2(PathFinder_15_io_i_mux_bus_2),
    .io_i_mux_bus_3(PathFinder_15_io_i_mux_bus_3),
    .io_Source_0(PathFinder_15_io_Source_0),
    .io_Source_1(PathFinder_15_io_Source_1),
    .io_Source_2(PathFinder_15_io_Source_2),
    .io_Source_3(PathFinder_15_io_Source_3),
    .io_PF_Valid(PathFinder_15_io_PF_Valid),
    .io_NoDPE(PathFinder_15_io_NoDPE),
    .io_DataValid(PathFinder_15_io_DataValid)
  );
  ivntop ivntop ( // @[FlexDPU.scala 87:21]
    .clock(ivntop_clock),
    .reset(ivntop_reset),
    .io_ProcessValid(ivntop_io_ProcessValid),
    .io_Stationary_matrix_0_0(ivntop_io_Stationary_matrix_0_0),
    .io_Stationary_matrix_0_1(ivntop_io_Stationary_matrix_0_1),
    .io_Stationary_matrix_0_2(ivntop_io_Stationary_matrix_0_2),
    .io_Stationary_matrix_0_3(ivntop_io_Stationary_matrix_0_3),
    .io_Stationary_matrix_0_4(ivntop_io_Stationary_matrix_0_4),
    .io_Stationary_matrix_0_5(ivntop_io_Stationary_matrix_0_5),
    .io_Stationary_matrix_0_6(ivntop_io_Stationary_matrix_0_6),
    .io_Stationary_matrix_0_7(ivntop_io_Stationary_matrix_0_7),
    .io_Stationary_matrix_1_0(ivntop_io_Stationary_matrix_1_0),
    .io_Stationary_matrix_1_1(ivntop_io_Stationary_matrix_1_1),
    .io_Stationary_matrix_1_2(ivntop_io_Stationary_matrix_1_2),
    .io_Stationary_matrix_1_3(ivntop_io_Stationary_matrix_1_3),
    .io_Stationary_matrix_1_4(ivntop_io_Stationary_matrix_1_4),
    .io_Stationary_matrix_1_5(ivntop_io_Stationary_matrix_1_5),
    .io_Stationary_matrix_1_6(ivntop_io_Stationary_matrix_1_6),
    .io_Stationary_matrix_1_7(ivntop_io_Stationary_matrix_1_7),
    .io_Stationary_matrix_2_0(ivntop_io_Stationary_matrix_2_0),
    .io_Stationary_matrix_2_1(ivntop_io_Stationary_matrix_2_1),
    .io_Stationary_matrix_2_2(ivntop_io_Stationary_matrix_2_2),
    .io_Stationary_matrix_2_3(ivntop_io_Stationary_matrix_2_3),
    .io_Stationary_matrix_2_4(ivntop_io_Stationary_matrix_2_4),
    .io_Stationary_matrix_2_5(ivntop_io_Stationary_matrix_2_5),
    .io_Stationary_matrix_2_6(ivntop_io_Stationary_matrix_2_6),
    .io_Stationary_matrix_2_7(ivntop_io_Stationary_matrix_2_7),
    .io_Stationary_matrix_3_0(ivntop_io_Stationary_matrix_3_0),
    .io_Stationary_matrix_3_1(ivntop_io_Stationary_matrix_3_1),
    .io_Stationary_matrix_3_2(ivntop_io_Stationary_matrix_3_2),
    .io_Stationary_matrix_3_3(ivntop_io_Stationary_matrix_3_3),
    .io_Stationary_matrix_3_4(ivntop_io_Stationary_matrix_3_4),
    .io_Stationary_matrix_3_5(ivntop_io_Stationary_matrix_3_5),
    .io_Stationary_matrix_3_6(ivntop_io_Stationary_matrix_3_6),
    .io_Stationary_matrix_3_7(ivntop_io_Stationary_matrix_3_7),
    .io_Stationary_matrix_4_0(ivntop_io_Stationary_matrix_4_0),
    .io_Stationary_matrix_4_1(ivntop_io_Stationary_matrix_4_1),
    .io_Stationary_matrix_4_2(ivntop_io_Stationary_matrix_4_2),
    .io_Stationary_matrix_4_3(ivntop_io_Stationary_matrix_4_3),
    .io_Stationary_matrix_4_4(ivntop_io_Stationary_matrix_4_4),
    .io_Stationary_matrix_4_5(ivntop_io_Stationary_matrix_4_5),
    .io_Stationary_matrix_4_6(ivntop_io_Stationary_matrix_4_6),
    .io_Stationary_matrix_4_7(ivntop_io_Stationary_matrix_4_7),
    .io_Stationary_matrix_5_0(ivntop_io_Stationary_matrix_5_0),
    .io_Stationary_matrix_5_1(ivntop_io_Stationary_matrix_5_1),
    .io_Stationary_matrix_5_2(ivntop_io_Stationary_matrix_5_2),
    .io_Stationary_matrix_5_3(ivntop_io_Stationary_matrix_5_3),
    .io_Stationary_matrix_5_4(ivntop_io_Stationary_matrix_5_4),
    .io_Stationary_matrix_5_5(ivntop_io_Stationary_matrix_5_5),
    .io_Stationary_matrix_5_6(ivntop_io_Stationary_matrix_5_6),
    .io_Stationary_matrix_5_7(ivntop_io_Stationary_matrix_5_7),
    .io_Stationary_matrix_6_0(ivntop_io_Stationary_matrix_6_0),
    .io_Stationary_matrix_6_1(ivntop_io_Stationary_matrix_6_1),
    .io_Stationary_matrix_6_2(ivntop_io_Stationary_matrix_6_2),
    .io_Stationary_matrix_6_3(ivntop_io_Stationary_matrix_6_3),
    .io_Stationary_matrix_6_4(ivntop_io_Stationary_matrix_6_4),
    .io_Stationary_matrix_6_5(ivntop_io_Stationary_matrix_6_5),
    .io_Stationary_matrix_6_6(ivntop_io_Stationary_matrix_6_6),
    .io_Stationary_matrix_6_7(ivntop_io_Stationary_matrix_6_7),
    .io_Stationary_matrix_7_0(ivntop_io_Stationary_matrix_7_0),
    .io_Stationary_matrix_7_1(ivntop_io_Stationary_matrix_7_1),
    .io_Stationary_matrix_7_2(ivntop_io_Stationary_matrix_7_2),
    .io_Stationary_matrix_7_3(ivntop_io_Stationary_matrix_7_3),
    .io_Stationary_matrix_7_4(ivntop_io_Stationary_matrix_7_4),
    .io_Stationary_matrix_7_5(ivntop_io_Stationary_matrix_7_5),
    .io_Stationary_matrix_7_6(ivntop_io_Stationary_matrix_7_6),
    .io_Stationary_matrix_7_7(ivntop_io_Stationary_matrix_7_7),
    .io_o_vn_0_0(ivntop_io_o_vn_0_0),
    .io_o_vn_0_1(ivntop_io_o_vn_0_1),
    .io_o_vn_0_2(ivntop_io_o_vn_0_2),
    .io_o_vn_0_3(ivntop_io_o_vn_0_3),
    .io_o_vn_1_0(ivntop_io_o_vn_1_0),
    .io_o_vn_1_1(ivntop_io_o_vn_1_1),
    .io_o_vn_1_2(ivntop_io_o_vn_1_2),
    .io_o_vn_1_3(ivntop_io_o_vn_1_3),
    .io_o_vn_2_0(ivntop_io_o_vn_2_0),
    .io_o_vn_2_1(ivntop_io_o_vn_2_1),
    .io_o_vn_2_2(ivntop_io_o_vn_2_2),
    .io_o_vn_2_3(ivntop_io_o_vn_2_3),
    .io_o_vn_3_0(ivntop_io_o_vn_3_0),
    .io_o_vn_3_1(ivntop_io_o_vn_3_1),
    .io_o_vn_3_2(ivntop_io_o_vn_3_2),
    .io_o_vn_3_3(ivntop_io_o_vn_3_3),
    .io_o_vn_4_0(ivntop_io_o_vn_4_0),
    .io_o_vn_4_1(ivntop_io_o_vn_4_1),
    .io_o_vn_4_2(ivntop_io_o_vn_4_2),
    .io_o_vn_4_3(ivntop_io_o_vn_4_3),
    .io_o_vn_5_0(ivntop_io_o_vn_5_0),
    .io_o_vn_5_1(ivntop_io_o_vn_5_1),
    .io_o_vn_5_2(ivntop_io_o_vn_5_2),
    .io_o_vn_5_3(ivntop_io_o_vn_5_3),
    .io_o_vn_6_0(ivntop_io_o_vn_6_0),
    .io_o_vn_6_1(ivntop_io_o_vn_6_1),
    .io_o_vn_6_2(ivntop_io_o_vn_6_2),
    .io_o_vn_6_3(ivntop_io_o_vn_6_3),
    .io_o_vn_7_0(ivntop_io_o_vn_7_0),
    .io_o_vn_7_1(ivntop_io_o_vn_7_1),
    .io_o_vn_7_2(ivntop_io_o_vn_7_2),
    .io_o_vn_7_3(ivntop_io_o_vn_7_3),
    .io_o_vn_8_0(ivntop_io_o_vn_8_0),
    .io_o_vn_8_1(ivntop_io_o_vn_8_1),
    .io_o_vn_8_2(ivntop_io_o_vn_8_2),
    .io_o_vn_8_3(ivntop_io_o_vn_8_3),
    .io_o_vn_9_0(ivntop_io_o_vn_9_0),
    .io_o_vn_9_1(ivntop_io_o_vn_9_1),
    .io_o_vn_9_2(ivntop_io_o_vn_9_2),
    .io_o_vn_9_3(ivntop_io_o_vn_9_3),
    .io_o_vn_10_0(ivntop_io_o_vn_10_0),
    .io_o_vn_10_1(ivntop_io_o_vn_10_1),
    .io_o_vn_10_2(ivntop_io_o_vn_10_2),
    .io_o_vn_10_3(ivntop_io_o_vn_10_3),
    .io_o_vn_11_0(ivntop_io_o_vn_11_0),
    .io_o_vn_11_1(ivntop_io_o_vn_11_1),
    .io_o_vn_11_2(ivntop_io_o_vn_11_2),
    .io_o_vn_11_3(ivntop_io_o_vn_11_3),
    .io_o_vn_12_0(ivntop_io_o_vn_12_0),
    .io_o_vn_12_1(ivntop_io_o_vn_12_1),
    .io_o_vn_12_2(ivntop_io_o_vn_12_2),
    .io_o_vn_12_3(ivntop_io_o_vn_12_3),
    .io_o_vn_13_0(ivntop_io_o_vn_13_0),
    .io_o_vn_13_1(ivntop_io_o_vn_13_1),
    .io_o_vn_13_2(ivntop_io_o_vn_13_2),
    .io_o_vn_13_3(ivntop_io_o_vn_13_3),
    .io_o_vn_14_0(ivntop_io_o_vn_14_0),
    .io_o_vn_14_1(ivntop_io_o_vn_14_1),
    .io_o_vn_14_2(ivntop_io_o_vn_14_2),
    .io_o_vn_14_3(ivntop_io_o_vn_14_3),
    .io_o_vn_15_0(ivntop_io_o_vn_15_0),
    .io_o_vn_15_1(ivntop_io_o_vn_15_1),
    .io_o_vn_15_2(ivntop_io_o_vn_15_2),
    .io_o_vn_15_3(ivntop_io_o_vn_15_3)
  );
  MuxesWrapper MuxesWrapper ( // @[FlexDPU.scala 124:53]
    .io_valid(MuxesWrapper_io_valid),
    .io_src_0(MuxesWrapper_io_src_0),
    .io_src_1(MuxesWrapper_io_src_1),
    .io_src_2(MuxesWrapper_io_src_2),
    .io_src_3(MuxesWrapper_io_src_3),
    .io_muxes_0(MuxesWrapper_io_muxes_0),
    .io_muxes_1(MuxesWrapper_io_muxes_1),
    .io_muxes_2(MuxesWrapper_io_muxes_2),
    .io_muxes_3(MuxesWrapper_io_muxes_3),
    .io_Osrc_0(MuxesWrapper_io_Osrc_0),
    .io_Osrc_1(MuxesWrapper_io_Osrc_1),
    .io_Osrc_2(MuxesWrapper_io_Osrc_2),
    .io_Osrc_3(MuxesWrapper_io_Osrc_3),
    .io_Omuxes_0_0(MuxesWrapper_io_Omuxes_0_0),
    .io_Omuxes_0_1(MuxesWrapper_io_Omuxes_0_1),
    .io_Omuxes_0_2(MuxesWrapper_io_Omuxes_0_2),
    .io_Omuxes_0_3(MuxesWrapper_io_Omuxes_0_3),
    .io_Omuxes_1_0(MuxesWrapper_io_Omuxes_1_0),
    .io_Omuxes_1_1(MuxesWrapper_io_Omuxes_1_1),
    .io_Omuxes_1_2(MuxesWrapper_io_Omuxes_1_2),
    .io_Omuxes_2_0(MuxesWrapper_io_Omuxes_2_0),
    .io_Omuxes_2_1(MuxesWrapper_io_Omuxes_2_1),
    .io_Omuxes_3_0(MuxesWrapper_io_Omuxes_3_0)
  );
  MuxesWrapper MuxesWrapper_1 ( // @[FlexDPU.scala 124:53]
    .io_valid(MuxesWrapper_1_io_valid),
    .io_src_0(MuxesWrapper_1_io_src_0),
    .io_src_1(MuxesWrapper_1_io_src_1),
    .io_src_2(MuxesWrapper_1_io_src_2),
    .io_src_3(MuxesWrapper_1_io_src_3),
    .io_muxes_0(MuxesWrapper_1_io_muxes_0),
    .io_muxes_1(MuxesWrapper_1_io_muxes_1),
    .io_muxes_2(MuxesWrapper_1_io_muxes_2),
    .io_muxes_3(MuxesWrapper_1_io_muxes_3),
    .io_Osrc_0(MuxesWrapper_1_io_Osrc_0),
    .io_Osrc_1(MuxesWrapper_1_io_Osrc_1),
    .io_Osrc_2(MuxesWrapper_1_io_Osrc_2),
    .io_Osrc_3(MuxesWrapper_1_io_Osrc_3),
    .io_Omuxes_0_0(MuxesWrapper_1_io_Omuxes_0_0),
    .io_Omuxes_0_1(MuxesWrapper_1_io_Omuxes_0_1),
    .io_Omuxes_0_2(MuxesWrapper_1_io_Omuxes_0_2),
    .io_Omuxes_0_3(MuxesWrapper_1_io_Omuxes_0_3),
    .io_Omuxes_1_0(MuxesWrapper_1_io_Omuxes_1_0),
    .io_Omuxes_1_1(MuxesWrapper_1_io_Omuxes_1_1),
    .io_Omuxes_1_2(MuxesWrapper_1_io_Omuxes_1_2),
    .io_Omuxes_2_0(MuxesWrapper_1_io_Omuxes_2_0),
    .io_Omuxes_2_1(MuxesWrapper_1_io_Omuxes_2_1),
    .io_Omuxes_3_0(MuxesWrapper_1_io_Omuxes_3_0)
  );
  MuxesWrapper MuxesWrapper_2 ( // @[FlexDPU.scala 124:53]
    .io_valid(MuxesWrapper_2_io_valid),
    .io_src_0(MuxesWrapper_2_io_src_0),
    .io_src_1(MuxesWrapper_2_io_src_1),
    .io_src_2(MuxesWrapper_2_io_src_2),
    .io_src_3(MuxesWrapper_2_io_src_3),
    .io_muxes_0(MuxesWrapper_2_io_muxes_0),
    .io_muxes_1(MuxesWrapper_2_io_muxes_1),
    .io_muxes_2(MuxesWrapper_2_io_muxes_2),
    .io_muxes_3(MuxesWrapper_2_io_muxes_3),
    .io_Osrc_0(MuxesWrapper_2_io_Osrc_0),
    .io_Osrc_1(MuxesWrapper_2_io_Osrc_1),
    .io_Osrc_2(MuxesWrapper_2_io_Osrc_2),
    .io_Osrc_3(MuxesWrapper_2_io_Osrc_3),
    .io_Omuxes_0_0(MuxesWrapper_2_io_Omuxes_0_0),
    .io_Omuxes_0_1(MuxesWrapper_2_io_Omuxes_0_1),
    .io_Omuxes_0_2(MuxesWrapper_2_io_Omuxes_0_2),
    .io_Omuxes_0_3(MuxesWrapper_2_io_Omuxes_0_3),
    .io_Omuxes_1_0(MuxesWrapper_2_io_Omuxes_1_0),
    .io_Omuxes_1_1(MuxesWrapper_2_io_Omuxes_1_1),
    .io_Omuxes_1_2(MuxesWrapper_2_io_Omuxes_1_2),
    .io_Omuxes_2_0(MuxesWrapper_2_io_Omuxes_2_0),
    .io_Omuxes_2_1(MuxesWrapper_2_io_Omuxes_2_1),
    .io_Omuxes_3_0(MuxesWrapper_2_io_Omuxes_3_0)
  );
  MuxesWrapper MuxesWrapper_3 ( // @[FlexDPU.scala 124:53]
    .io_valid(MuxesWrapper_3_io_valid),
    .io_src_0(MuxesWrapper_3_io_src_0),
    .io_src_1(MuxesWrapper_3_io_src_1),
    .io_src_2(MuxesWrapper_3_io_src_2),
    .io_src_3(MuxesWrapper_3_io_src_3),
    .io_muxes_0(MuxesWrapper_3_io_muxes_0),
    .io_muxes_1(MuxesWrapper_3_io_muxes_1),
    .io_muxes_2(MuxesWrapper_3_io_muxes_2),
    .io_muxes_3(MuxesWrapper_3_io_muxes_3),
    .io_Osrc_0(MuxesWrapper_3_io_Osrc_0),
    .io_Osrc_1(MuxesWrapper_3_io_Osrc_1),
    .io_Osrc_2(MuxesWrapper_3_io_Osrc_2),
    .io_Osrc_3(MuxesWrapper_3_io_Osrc_3),
    .io_Omuxes_0_0(MuxesWrapper_3_io_Omuxes_0_0),
    .io_Omuxes_0_1(MuxesWrapper_3_io_Omuxes_0_1),
    .io_Omuxes_0_2(MuxesWrapper_3_io_Omuxes_0_2),
    .io_Omuxes_0_3(MuxesWrapper_3_io_Omuxes_0_3),
    .io_Omuxes_1_0(MuxesWrapper_3_io_Omuxes_1_0),
    .io_Omuxes_1_1(MuxesWrapper_3_io_Omuxes_1_1),
    .io_Omuxes_1_2(MuxesWrapper_3_io_Omuxes_1_2),
    .io_Omuxes_2_0(MuxesWrapper_3_io_Omuxes_2_0),
    .io_Omuxes_2_1(MuxesWrapper_3_io_Omuxes_2_1),
    .io_Omuxes_3_0(MuxesWrapper_3_io_Omuxes_3_0)
  );
  MuxesWrapper MuxesWrapper_4 ( // @[FlexDPU.scala 124:53]
    .io_valid(MuxesWrapper_4_io_valid),
    .io_src_0(MuxesWrapper_4_io_src_0),
    .io_src_1(MuxesWrapper_4_io_src_1),
    .io_src_2(MuxesWrapper_4_io_src_2),
    .io_src_3(MuxesWrapper_4_io_src_3),
    .io_muxes_0(MuxesWrapper_4_io_muxes_0),
    .io_muxes_1(MuxesWrapper_4_io_muxes_1),
    .io_muxes_2(MuxesWrapper_4_io_muxes_2),
    .io_muxes_3(MuxesWrapper_4_io_muxes_3),
    .io_Osrc_0(MuxesWrapper_4_io_Osrc_0),
    .io_Osrc_1(MuxesWrapper_4_io_Osrc_1),
    .io_Osrc_2(MuxesWrapper_4_io_Osrc_2),
    .io_Osrc_3(MuxesWrapper_4_io_Osrc_3),
    .io_Omuxes_0_0(MuxesWrapper_4_io_Omuxes_0_0),
    .io_Omuxes_0_1(MuxesWrapper_4_io_Omuxes_0_1),
    .io_Omuxes_0_2(MuxesWrapper_4_io_Omuxes_0_2),
    .io_Omuxes_0_3(MuxesWrapper_4_io_Omuxes_0_3),
    .io_Omuxes_1_0(MuxesWrapper_4_io_Omuxes_1_0),
    .io_Omuxes_1_1(MuxesWrapper_4_io_Omuxes_1_1),
    .io_Omuxes_1_2(MuxesWrapper_4_io_Omuxes_1_2),
    .io_Omuxes_2_0(MuxesWrapper_4_io_Omuxes_2_0),
    .io_Omuxes_2_1(MuxesWrapper_4_io_Omuxes_2_1),
    .io_Omuxes_3_0(MuxesWrapper_4_io_Omuxes_3_0)
  );
  MuxesWrapper MuxesWrapper_5 ( // @[FlexDPU.scala 124:53]
    .io_valid(MuxesWrapper_5_io_valid),
    .io_src_0(MuxesWrapper_5_io_src_0),
    .io_src_1(MuxesWrapper_5_io_src_1),
    .io_src_2(MuxesWrapper_5_io_src_2),
    .io_src_3(MuxesWrapper_5_io_src_3),
    .io_muxes_0(MuxesWrapper_5_io_muxes_0),
    .io_muxes_1(MuxesWrapper_5_io_muxes_1),
    .io_muxes_2(MuxesWrapper_5_io_muxes_2),
    .io_muxes_3(MuxesWrapper_5_io_muxes_3),
    .io_Osrc_0(MuxesWrapper_5_io_Osrc_0),
    .io_Osrc_1(MuxesWrapper_5_io_Osrc_1),
    .io_Osrc_2(MuxesWrapper_5_io_Osrc_2),
    .io_Osrc_3(MuxesWrapper_5_io_Osrc_3),
    .io_Omuxes_0_0(MuxesWrapper_5_io_Omuxes_0_0),
    .io_Omuxes_0_1(MuxesWrapper_5_io_Omuxes_0_1),
    .io_Omuxes_0_2(MuxesWrapper_5_io_Omuxes_0_2),
    .io_Omuxes_0_3(MuxesWrapper_5_io_Omuxes_0_3),
    .io_Omuxes_1_0(MuxesWrapper_5_io_Omuxes_1_0),
    .io_Omuxes_1_1(MuxesWrapper_5_io_Omuxes_1_1),
    .io_Omuxes_1_2(MuxesWrapper_5_io_Omuxes_1_2),
    .io_Omuxes_2_0(MuxesWrapper_5_io_Omuxes_2_0),
    .io_Omuxes_2_1(MuxesWrapper_5_io_Omuxes_2_1),
    .io_Omuxes_3_0(MuxesWrapper_5_io_Omuxes_3_0)
  );
  MuxesWrapper MuxesWrapper_6 ( // @[FlexDPU.scala 124:53]
    .io_valid(MuxesWrapper_6_io_valid),
    .io_src_0(MuxesWrapper_6_io_src_0),
    .io_src_1(MuxesWrapper_6_io_src_1),
    .io_src_2(MuxesWrapper_6_io_src_2),
    .io_src_3(MuxesWrapper_6_io_src_3),
    .io_muxes_0(MuxesWrapper_6_io_muxes_0),
    .io_muxes_1(MuxesWrapper_6_io_muxes_1),
    .io_muxes_2(MuxesWrapper_6_io_muxes_2),
    .io_muxes_3(MuxesWrapper_6_io_muxes_3),
    .io_Osrc_0(MuxesWrapper_6_io_Osrc_0),
    .io_Osrc_1(MuxesWrapper_6_io_Osrc_1),
    .io_Osrc_2(MuxesWrapper_6_io_Osrc_2),
    .io_Osrc_3(MuxesWrapper_6_io_Osrc_3),
    .io_Omuxes_0_0(MuxesWrapper_6_io_Omuxes_0_0),
    .io_Omuxes_0_1(MuxesWrapper_6_io_Omuxes_0_1),
    .io_Omuxes_0_2(MuxesWrapper_6_io_Omuxes_0_2),
    .io_Omuxes_0_3(MuxesWrapper_6_io_Omuxes_0_3),
    .io_Omuxes_1_0(MuxesWrapper_6_io_Omuxes_1_0),
    .io_Omuxes_1_1(MuxesWrapper_6_io_Omuxes_1_1),
    .io_Omuxes_1_2(MuxesWrapper_6_io_Omuxes_1_2),
    .io_Omuxes_2_0(MuxesWrapper_6_io_Omuxes_2_0),
    .io_Omuxes_2_1(MuxesWrapper_6_io_Omuxes_2_1),
    .io_Omuxes_3_0(MuxesWrapper_6_io_Omuxes_3_0)
  );
  MuxesWrapper MuxesWrapper_7 ( // @[FlexDPU.scala 124:53]
    .io_valid(MuxesWrapper_7_io_valid),
    .io_src_0(MuxesWrapper_7_io_src_0),
    .io_src_1(MuxesWrapper_7_io_src_1),
    .io_src_2(MuxesWrapper_7_io_src_2),
    .io_src_3(MuxesWrapper_7_io_src_3),
    .io_muxes_0(MuxesWrapper_7_io_muxes_0),
    .io_muxes_1(MuxesWrapper_7_io_muxes_1),
    .io_muxes_2(MuxesWrapper_7_io_muxes_2),
    .io_muxes_3(MuxesWrapper_7_io_muxes_3),
    .io_Osrc_0(MuxesWrapper_7_io_Osrc_0),
    .io_Osrc_1(MuxesWrapper_7_io_Osrc_1),
    .io_Osrc_2(MuxesWrapper_7_io_Osrc_2),
    .io_Osrc_3(MuxesWrapper_7_io_Osrc_3),
    .io_Omuxes_0_0(MuxesWrapper_7_io_Omuxes_0_0),
    .io_Omuxes_0_1(MuxesWrapper_7_io_Omuxes_0_1),
    .io_Omuxes_0_2(MuxesWrapper_7_io_Omuxes_0_2),
    .io_Omuxes_0_3(MuxesWrapper_7_io_Omuxes_0_3),
    .io_Omuxes_1_0(MuxesWrapper_7_io_Omuxes_1_0),
    .io_Omuxes_1_1(MuxesWrapper_7_io_Omuxes_1_1),
    .io_Omuxes_1_2(MuxesWrapper_7_io_Omuxes_1_2),
    .io_Omuxes_2_0(MuxesWrapper_7_io_Omuxes_2_0),
    .io_Omuxes_2_1(MuxesWrapper_7_io_Omuxes_2_1),
    .io_Omuxes_3_0(MuxesWrapper_7_io_Omuxes_3_0)
  );
  MuxesWrapper MuxesWrapper_8 ( // @[FlexDPU.scala 124:53]
    .io_valid(MuxesWrapper_8_io_valid),
    .io_src_0(MuxesWrapper_8_io_src_0),
    .io_src_1(MuxesWrapper_8_io_src_1),
    .io_src_2(MuxesWrapper_8_io_src_2),
    .io_src_3(MuxesWrapper_8_io_src_3),
    .io_muxes_0(MuxesWrapper_8_io_muxes_0),
    .io_muxes_1(MuxesWrapper_8_io_muxes_1),
    .io_muxes_2(MuxesWrapper_8_io_muxes_2),
    .io_muxes_3(MuxesWrapper_8_io_muxes_3),
    .io_Osrc_0(MuxesWrapper_8_io_Osrc_0),
    .io_Osrc_1(MuxesWrapper_8_io_Osrc_1),
    .io_Osrc_2(MuxesWrapper_8_io_Osrc_2),
    .io_Osrc_3(MuxesWrapper_8_io_Osrc_3),
    .io_Omuxes_0_0(MuxesWrapper_8_io_Omuxes_0_0),
    .io_Omuxes_0_1(MuxesWrapper_8_io_Omuxes_0_1),
    .io_Omuxes_0_2(MuxesWrapper_8_io_Omuxes_0_2),
    .io_Omuxes_0_3(MuxesWrapper_8_io_Omuxes_0_3),
    .io_Omuxes_1_0(MuxesWrapper_8_io_Omuxes_1_0),
    .io_Omuxes_1_1(MuxesWrapper_8_io_Omuxes_1_1),
    .io_Omuxes_1_2(MuxesWrapper_8_io_Omuxes_1_2),
    .io_Omuxes_2_0(MuxesWrapper_8_io_Omuxes_2_0),
    .io_Omuxes_2_1(MuxesWrapper_8_io_Omuxes_2_1),
    .io_Omuxes_3_0(MuxesWrapper_8_io_Omuxes_3_0)
  );
  MuxesWrapper MuxesWrapper_9 ( // @[FlexDPU.scala 124:53]
    .io_valid(MuxesWrapper_9_io_valid),
    .io_src_0(MuxesWrapper_9_io_src_0),
    .io_src_1(MuxesWrapper_9_io_src_1),
    .io_src_2(MuxesWrapper_9_io_src_2),
    .io_src_3(MuxesWrapper_9_io_src_3),
    .io_muxes_0(MuxesWrapper_9_io_muxes_0),
    .io_muxes_1(MuxesWrapper_9_io_muxes_1),
    .io_muxes_2(MuxesWrapper_9_io_muxes_2),
    .io_muxes_3(MuxesWrapper_9_io_muxes_3),
    .io_Osrc_0(MuxesWrapper_9_io_Osrc_0),
    .io_Osrc_1(MuxesWrapper_9_io_Osrc_1),
    .io_Osrc_2(MuxesWrapper_9_io_Osrc_2),
    .io_Osrc_3(MuxesWrapper_9_io_Osrc_3),
    .io_Omuxes_0_0(MuxesWrapper_9_io_Omuxes_0_0),
    .io_Omuxes_0_1(MuxesWrapper_9_io_Omuxes_0_1),
    .io_Omuxes_0_2(MuxesWrapper_9_io_Omuxes_0_2),
    .io_Omuxes_0_3(MuxesWrapper_9_io_Omuxes_0_3),
    .io_Omuxes_1_0(MuxesWrapper_9_io_Omuxes_1_0),
    .io_Omuxes_1_1(MuxesWrapper_9_io_Omuxes_1_1),
    .io_Omuxes_1_2(MuxesWrapper_9_io_Omuxes_1_2),
    .io_Omuxes_2_0(MuxesWrapper_9_io_Omuxes_2_0),
    .io_Omuxes_2_1(MuxesWrapper_9_io_Omuxes_2_1),
    .io_Omuxes_3_0(MuxesWrapper_9_io_Omuxes_3_0)
  );
  MuxesWrapper MuxesWrapper_10 ( // @[FlexDPU.scala 124:53]
    .io_valid(MuxesWrapper_10_io_valid),
    .io_src_0(MuxesWrapper_10_io_src_0),
    .io_src_1(MuxesWrapper_10_io_src_1),
    .io_src_2(MuxesWrapper_10_io_src_2),
    .io_src_3(MuxesWrapper_10_io_src_3),
    .io_muxes_0(MuxesWrapper_10_io_muxes_0),
    .io_muxes_1(MuxesWrapper_10_io_muxes_1),
    .io_muxes_2(MuxesWrapper_10_io_muxes_2),
    .io_muxes_3(MuxesWrapper_10_io_muxes_3),
    .io_Osrc_0(MuxesWrapper_10_io_Osrc_0),
    .io_Osrc_1(MuxesWrapper_10_io_Osrc_1),
    .io_Osrc_2(MuxesWrapper_10_io_Osrc_2),
    .io_Osrc_3(MuxesWrapper_10_io_Osrc_3),
    .io_Omuxes_0_0(MuxesWrapper_10_io_Omuxes_0_0),
    .io_Omuxes_0_1(MuxesWrapper_10_io_Omuxes_0_1),
    .io_Omuxes_0_2(MuxesWrapper_10_io_Omuxes_0_2),
    .io_Omuxes_0_3(MuxesWrapper_10_io_Omuxes_0_3),
    .io_Omuxes_1_0(MuxesWrapper_10_io_Omuxes_1_0),
    .io_Omuxes_1_1(MuxesWrapper_10_io_Omuxes_1_1),
    .io_Omuxes_1_2(MuxesWrapper_10_io_Omuxes_1_2),
    .io_Omuxes_2_0(MuxesWrapper_10_io_Omuxes_2_0),
    .io_Omuxes_2_1(MuxesWrapper_10_io_Omuxes_2_1),
    .io_Omuxes_3_0(MuxesWrapper_10_io_Omuxes_3_0)
  );
  MuxesWrapper MuxesWrapper_11 ( // @[FlexDPU.scala 124:53]
    .io_valid(MuxesWrapper_11_io_valid),
    .io_src_0(MuxesWrapper_11_io_src_0),
    .io_src_1(MuxesWrapper_11_io_src_1),
    .io_src_2(MuxesWrapper_11_io_src_2),
    .io_src_3(MuxesWrapper_11_io_src_3),
    .io_muxes_0(MuxesWrapper_11_io_muxes_0),
    .io_muxes_1(MuxesWrapper_11_io_muxes_1),
    .io_muxes_2(MuxesWrapper_11_io_muxes_2),
    .io_muxes_3(MuxesWrapper_11_io_muxes_3),
    .io_Osrc_0(MuxesWrapper_11_io_Osrc_0),
    .io_Osrc_1(MuxesWrapper_11_io_Osrc_1),
    .io_Osrc_2(MuxesWrapper_11_io_Osrc_2),
    .io_Osrc_3(MuxesWrapper_11_io_Osrc_3),
    .io_Omuxes_0_0(MuxesWrapper_11_io_Omuxes_0_0),
    .io_Omuxes_0_1(MuxesWrapper_11_io_Omuxes_0_1),
    .io_Omuxes_0_2(MuxesWrapper_11_io_Omuxes_0_2),
    .io_Omuxes_0_3(MuxesWrapper_11_io_Omuxes_0_3),
    .io_Omuxes_1_0(MuxesWrapper_11_io_Omuxes_1_0),
    .io_Omuxes_1_1(MuxesWrapper_11_io_Omuxes_1_1),
    .io_Omuxes_1_2(MuxesWrapper_11_io_Omuxes_1_2),
    .io_Omuxes_2_0(MuxesWrapper_11_io_Omuxes_2_0),
    .io_Omuxes_2_1(MuxesWrapper_11_io_Omuxes_2_1),
    .io_Omuxes_3_0(MuxesWrapper_11_io_Omuxes_3_0)
  );
  MuxesWrapper MuxesWrapper_12 ( // @[FlexDPU.scala 124:53]
    .io_valid(MuxesWrapper_12_io_valid),
    .io_src_0(MuxesWrapper_12_io_src_0),
    .io_src_1(MuxesWrapper_12_io_src_1),
    .io_src_2(MuxesWrapper_12_io_src_2),
    .io_src_3(MuxesWrapper_12_io_src_3),
    .io_muxes_0(MuxesWrapper_12_io_muxes_0),
    .io_muxes_1(MuxesWrapper_12_io_muxes_1),
    .io_muxes_2(MuxesWrapper_12_io_muxes_2),
    .io_muxes_3(MuxesWrapper_12_io_muxes_3),
    .io_Osrc_0(MuxesWrapper_12_io_Osrc_0),
    .io_Osrc_1(MuxesWrapper_12_io_Osrc_1),
    .io_Osrc_2(MuxesWrapper_12_io_Osrc_2),
    .io_Osrc_3(MuxesWrapper_12_io_Osrc_3),
    .io_Omuxes_0_0(MuxesWrapper_12_io_Omuxes_0_0),
    .io_Omuxes_0_1(MuxesWrapper_12_io_Omuxes_0_1),
    .io_Omuxes_0_2(MuxesWrapper_12_io_Omuxes_0_2),
    .io_Omuxes_0_3(MuxesWrapper_12_io_Omuxes_0_3),
    .io_Omuxes_1_0(MuxesWrapper_12_io_Omuxes_1_0),
    .io_Omuxes_1_1(MuxesWrapper_12_io_Omuxes_1_1),
    .io_Omuxes_1_2(MuxesWrapper_12_io_Omuxes_1_2),
    .io_Omuxes_2_0(MuxesWrapper_12_io_Omuxes_2_0),
    .io_Omuxes_2_1(MuxesWrapper_12_io_Omuxes_2_1),
    .io_Omuxes_3_0(MuxesWrapper_12_io_Omuxes_3_0)
  );
  MuxesWrapper MuxesWrapper_13 ( // @[FlexDPU.scala 124:53]
    .io_valid(MuxesWrapper_13_io_valid),
    .io_src_0(MuxesWrapper_13_io_src_0),
    .io_src_1(MuxesWrapper_13_io_src_1),
    .io_src_2(MuxesWrapper_13_io_src_2),
    .io_src_3(MuxesWrapper_13_io_src_3),
    .io_muxes_0(MuxesWrapper_13_io_muxes_0),
    .io_muxes_1(MuxesWrapper_13_io_muxes_1),
    .io_muxes_2(MuxesWrapper_13_io_muxes_2),
    .io_muxes_3(MuxesWrapper_13_io_muxes_3),
    .io_Osrc_0(MuxesWrapper_13_io_Osrc_0),
    .io_Osrc_1(MuxesWrapper_13_io_Osrc_1),
    .io_Osrc_2(MuxesWrapper_13_io_Osrc_2),
    .io_Osrc_3(MuxesWrapper_13_io_Osrc_3),
    .io_Omuxes_0_0(MuxesWrapper_13_io_Omuxes_0_0),
    .io_Omuxes_0_1(MuxesWrapper_13_io_Omuxes_0_1),
    .io_Omuxes_0_2(MuxesWrapper_13_io_Omuxes_0_2),
    .io_Omuxes_0_3(MuxesWrapper_13_io_Omuxes_0_3),
    .io_Omuxes_1_0(MuxesWrapper_13_io_Omuxes_1_0),
    .io_Omuxes_1_1(MuxesWrapper_13_io_Omuxes_1_1),
    .io_Omuxes_1_2(MuxesWrapper_13_io_Omuxes_1_2),
    .io_Omuxes_2_0(MuxesWrapper_13_io_Omuxes_2_0),
    .io_Omuxes_2_1(MuxesWrapper_13_io_Omuxes_2_1),
    .io_Omuxes_3_0(MuxesWrapper_13_io_Omuxes_3_0)
  );
  MuxesWrapper MuxesWrapper_14 ( // @[FlexDPU.scala 124:53]
    .io_valid(MuxesWrapper_14_io_valid),
    .io_src_0(MuxesWrapper_14_io_src_0),
    .io_src_1(MuxesWrapper_14_io_src_1),
    .io_src_2(MuxesWrapper_14_io_src_2),
    .io_src_3(MuxesWrapper_14_io_src_3),
    .io_muxes_0(MuxesWrapper_14_io_muxes_0),
    .io_muxes_1(MuxesWrapper_14_io_muxes_1),
    .io_muxes_2(MuxesWrapper_14_io_muxes_2),
    .io_muxes_3(MuxesWrapper_14_io_muxes_3),
    .io_Osrc_0(MuxesWrapper_14_io_Osrc_0),
    .io_Osrc_1(MuxesWrapper_14_io_Osrc_1),
    .io_Osrc_2(MuxesWrapper_14_io_Osrc_2),
    .io_Osrc_3(MuxesWrapper_14_io_Osrc_3),
    .io_Omuxes_0_0(MuxesWrapper_14_io_Omuxes_0_0),
    .io_Omuxes_0_1(MuxesWrapper_14_io_Omuxes_0_1),
    .io_Omuxes_0_2(MuxesWrapper_14_io_Omuxes_0_2),
    .io_Omuxes_0_3(MuxesWrapper_14_io_Omuxes_0_3),
    .io_Omuxes_1_0(MuxesWrapper_14_io_Omuxes_1_0),
    .io_Omuxes_1_1(MuxesWrapper_14_io_Omuxes_1_1),
    .io_Omuxes_1_2(MuxesWrapper_14_io_Omuxes_1_2),
    .io_Omuxes_2_0(MuxesWrapper_14_io_Omuxes_2_0),
    .io_Omuxes_2_1(MuxesWrapper_14_io_Omuxes_2_1),
    .io_Omuxes_3_0(MuxesWrapper_14_io_Omuxes_3_0)
  );
  MuxesWrapper MuxesWrapper_15 ( // @[FlexDPU.scala 124:53]
    .io_valid(MuxesWrapper_15_io_valid),
    .io_src_0(MuxesWrapper_15_io_src_0),
    .io_src_1(MuxesWrapper_15_io_src_1),
    .io_src_2(MuxesWrapper_15_io_src_2),
    .io_src_3(MuxesWrapper_15_io_src_3),
    .io_muxes_0(MuxesWrapper_15_io_muxes_0),
    .io_muxes_1(MuxesWrapper_15_io_muxes_1),
    .io_muxes_2(MuxesWrapper_15_io_muxes_2),
    .io_muxes_3(MuxesWrapper_15_io_muxes_3),
    .io_Osrc_0(MuxesWrapper_15_io_Osrc_0),
    .io_Osrc_1(MuxesWrapper_15_io_Osrc_1),
    .io_Osrc_2(MuxesWrapper_15_io_Osrc_2),
    .io_Osrc_3(MuxesWrapper_15_io_Osrc_3),
    .io_Omuxes_0_0(MuxesWrapper_15_io_Omuxes_0_0),
    .io_Omuxes_0_1(MuxesWrapper_15_io_Omuxes_0_1),
    .io_Omuxes_0_2(MuxesWrapper_15_io_Omuxes_0_2),
    .io_Omuxes_0_3(MuxesWrapper_15_io_Omuxes_0_3),
    .io_Omuxes_1_0(MuxesWrapper_15_io_Omuxes_1_0),
    .io_Omuxes_1_1(MuxesWrapper_15_io_Omuxes_1_1),
    .io_Omuxes_1_2(MuxesWrapper_15_io_Omuxes_1_2),
    .io_Omuxes_2_0(MuxesWrapper_15_io_Omuxes_2_0),
    .io_Omuxes_2_1(MuxesWrapper_15_io_Omuxes_2_1),
    .io_Omuxes_3_0(MuxesWrapper_15_io_Omuxes_3_0)
  );
  flexdpecom4 flexdpecom4 ( // @[FlexDPU.scala 132:47]
    .clock(flexdpecom4_clock),
    .reset(flexdpecom4_reset),
    .io_i_data_valid(flexdpecom4_io_i_data_valid),
    .io_i_data_bus_0(flexdpecom4_io_i_data_bus_0),
    .io_i_data_bus_1(flexdpecom4_io_i_data_bus_1),
    .io_i_data_bus_2(flexdpecom4_io_i_data_bus_2),
    .io_i_data_bus_3(flexdpecom4_io_i_data_bus_3),
    .io_i_data_bus2_0(flexdpecom4_io_i_data_bus2_0),
    .io_i_data_bus2_1(flexdpecom4_io_i_data_bus2_1),
    .io_i_data_bus2_2(flexdpecom4_io_i_data_bus2_2),
    .io_i_data_bus2_3(flexdpecom4_io_i_data_bus2_3),
    .io_i_vn_0(flexdpecom4_io_i_vn_0),
    .io_i_vn_1(flexdpecom4_io_i_vn_1),
    .io_i_vn_2(flexdpecom4_io_i_vn_2),
    .io_i_vn_3(flexdpecom4_io_i_vn_3),
    .io_o_adder_0(flexdpecom4_io_o_adder_0),
    .io_o_adder_1(flexdpecom4_io_o_adder_1),
    .io_o_adder_2(flexdpecom4_io_o_adder_2),
    .io_i_mux_bus_0_0(flexdpecom4_io_i_mux_bus_0_0),
    .io_i_mux_bus_0_1(flexdpecom4_io_i_mux_bus_0_1),
    .io_i_mux_bus_0_2(flexdpecom4_io_i_mux_bus_0_2),
    .io_i_mux_bus_0_3(flexdpecom4_io_i_mux_bus_0_3),
    .io_i_mux_bus_1_0(flexdpecom4_io_i_mux_bus_1_0),
    .io_i_mux_bus_1_1(flexdpecom4_io_i_mux_bus_1_1),
    .io_i_mux_bus_1_2(flexdpecom4_io_i_mux_bus_1_2),
    .io_i_mux_bus_2_0(flexdpecom4_io_i_mux_bus_2_0),
    .io_i_mux_bus_2_1(flexdpecom4_io_i_mux_bus_2_1),
    .io_i_mux_bus_3_0(flexdpecom4_io_i_mux_bus_3_0)
  );
  flexdpecom4 flexdpecom4_1 ( // @[FlexDPU.scala 132:47]
    .clock(flexdpecom4_1_clock),
    .reset(flexdpecom4_1_reset),
    .io_i_data_valid(flexdpecom4_1_io_i_data_valid),
    .io_i_data_bus_0(flexdpecom4_1_io_i_data_bus_0),
    .io_i_data_bus_1(flexdpecom4_1_io_i_data_bus_1),
    .io_i_data_bus_2(flexdpecom4_1_io_i_data_bus_2),
    .io_i_data_bus_3(flexdpecom4_1_io_i_data_bus_3),
    .io_i_data_bus2_0(flexdpecom4_1_io_i_data_bus2_0),
    .io_i_data_bus2_1(flexdpecom4_1_io_i_data_bus2_1),
    .io_i_data_bus2_2(flexdpecom4_1_io_i_data_bus2_2),
    .io_i_data_bus2_3(flexdpecom4_1_io_i_data_bus2_3),
    .io_i_vn_0(flexdpecom4_1_io_i_vn_0),
    .io_i_vn_1(flexdpecom4_1_io_i_vn_1),
    .io_i_vn_2(flexdpecom4_1_io_i_vn_2),
    .io_i_vn_3(flexdpecom4_1_io_i_vn_3),
    .io_o_adder_0(flexdpecom4_1_io_o_adder_0),
    .io_o_adder_1(flexdpecom4_1_io_o_adder_1),
    .io_o_adder_2(flexdpecom4_1_io_o_adder_2),
    .io_i_mux_bus_0_0(flexdpecom4_1_io_i_mux_bus_0_0),
    .io_i_mux_bus_0_1(flexdpecom4_1_io_i_mux_bus_0_1),
    .io_i_mux_bus_0_2(flexdpecom4_1_io_i_mux_bus_0_2),
    .io_i_mux_bus_0_3(flexdpecom4_1_io_i_mux_bus_0_3),
    .io_i_mux_bus_1_0(flexdpecom4_1_io_i_mux_bus_1_0),
    .io_i_mux_bus_1_1(flexdpecom4_1_io_i_mux_bus_1_1),
    .io_i_mux_bus_1_2(flexdpecom4_1_io_i_mux_bus_1_2),
    .io_i_mux_bus_2_0(flexdpecom4_1_io_i_mux_bus_2_0),
    .io_i_mux_bus_2_1(flexdpecom4_1_io_i_mux_bus_2_1),
    .io_i_mux_bus_3_0(flexdpecom4_1_io_i_mux_bus_3_0)
  );
  flexdpecom4 flexdpecom4_2 ( // @[FlexDPU.scala 132:47]
    .clock(flexdpecom4_2_clock),
    .reset(flexdpecom4_2_reset),
    .io_i_data_valid(flexdpecom4_2_io_i_data_valid),
    .io_i_data_bus_0(flexdpecom4_2_io_i_data_bus_0),
    .io_i_data_bus_1(flexdpecom4_2_io_i_data_bus_1),
    .io_i_data_bus_2(flexdpecom4_2_io_i_data_bus_2),
    .io_i_data_bus_3(flexdpecom4_2_io_i_data_bus_3),
    .io_i_data_bus2_0(flexdpecom4_2_io_i_data_bus2_0),
    .io_i_data_bus2_1(flexdpecom4_2_io_i_data_bus2_1),
    .io_i_data_bus2_2(flexdpecom4_2_io_i_data_bus2_2),
    .io_i_data_bus2_3(flexdpecom4_2_io_i_data_bus2_3),
    .io_i_vn_0(flexdpecom4_2_io_i_vn_0),
    .io_i_vn_1(flexdpecom4_2_io_i_vn_1),
    .io_i_vn_2(flexdpecom4_2_io_i_vn_2),
    .io_i_vn_3(flexdpecom4_2_io_i_vn_3),
    .io_o_adder_0(flexdpecom4_2_io_o_adder_0),
    .io_o_adder_1(flexdpecom4_2_io_o_adder_1),
    .io_o_adder_2(flexdpecom4_2_io_o_adder_2),
    .io_i_mux_bus_0_0(flexdpecom4_2_io_i_mux_bus_0_0),
    .io_i_mux_bus_0_1(flexdpecom4_2_io_i_mux_bus_0_1),
    .io_i_mux_bus_0_2(flexdpecom4_2_io_i_mux_bus_0_2),
    .io_i_mux_bus_0_3(flexdpecom4_2_io_i_mux_bus_0_3),
    .io_i_mux_bus_1_0(flexdpecom4_2_io_i_mux_bus_1_0),
    .io_i_mux_bus_1_1(flexdpecom4_2_io_i_mux_bus_1_1),
    .io_i_mux_bus_1_2(flexdpecom4_2_io_i_mux_bus_1_2),
    .io_i_mux_bus_2_0(flexdpecom4_2_io_i_mux_bus_2_0),
    .io_i_mux_bus_2_1(flexdpecom4_2_io_i_mux_bus_2_1),
    .io_i_mux_bus_3_0(flexdpecom4_2_io_i_mux_bus_3_0)
  );
  flexdpecom4 flexdpecom4_3 ( // @[FlexDPU.scala 132:47]
    .clock(flexdpecom4_3_clock),
    .reset(flexdpecom4_3_reset),
    .io_i_data_valid(flexdpecom4_3_io_i_data_valid),
    .io_i_data_bus_0(flexdpecom4_3_io_i_data_bus_0),
    .io_i_data_bus_1(flexdpecom4_3_io_i_data_bus_1),
    .io_i_data_bus_2(flexdpecom4_3_io_i_data_bus_2),
    .io_i_data_bus_3(flexdpecom4_3_io_i_data_bus_3),
    .io_i_data_bus2_0(flexdpecom4_3_io_i_data_bus2_0),
    .io_i_data_bus2_1(flexdpecom4_3_io_i_data_bus2_1),
    .io_i_data_bus2_2(flexdpecom4_3_io_i_data_bus2_2),
    .io_i_data_bus2_3(flexdpecom4_3_io_i_data_bus2_3),
    .io_i_vn_0(flexdpecom4_3_io_i_vn_0),
    .io_i_vn_1(flexdpecom4_3_io_i_vn_1),
    .io_i_vn_2(flexdpecom4_3_io_i_vn_2),
    .io_i_vn_3(flexdpecom4_3_io_i_vn_3),
    .io_o_adder_0(flexdpecom4_3_io_o_adder_0),
    .io_o_adder_1(flexdpecom4_3_io_o_adder_1),
    .io_o_adder_2(flexdpecom4_3_io_o_adder_2),
    .io_i_mux_bus_0_0(flexdpecom4_3_io_i_mux_bus_0_0),
    .io_i_mux_bus_0_1(flexdpecom4_3_io_i_mux_bus_0_1),
    .io_i_mux_bus_0_2(flexdpecom4_3_io_i_mux_bus_0_2),
    .io_i_mux_bus_0_3(flexdpecom4_3_io_i_mux_bus_0_3),
    .io_i_mux_bus_1_0(flexdpecom4_3_io_i_mux_bus_1_0),
    .io_i_mux_bus_1_1(flexdpecom4_3_io_i_mux_bus_1_1),
    .io_i_mux_bus_1_2(flexdpecom4_3_io_i_mux_bus_1_2),
    .io_i_mux_bus_2_0(flexdpecom4_3_io_i_mux_bus_2_0),
    .io_i_mux_bus_2_1(flexdpecom4_3_io_i_mux_bus_2_1),
    .io_i_mux_bus_3_0(flexdpecom4_3_io_i_mux_bus_3_0)
  );
  flexdpecom4 flexdpecom4_4 ( // @[FlexDPU.scala 132:47]
    .clock(flexdpecom4_4_clock),
    .reset(flexdpecom4_4_reset),
    .io_i_data_valid(flexdpecom4_4_io_i_data_valid),
    .io_i_data_bus_0(flexdpecom4_4_io_i_data_bus_0),
    .io_i_data_bus_1(flexdpecom4_4_io_i_data_bus_1),
    .io_i_data_bus_2(flexdpecom4_4_io_i_data_bus_2),
    .io_i_data_bus_3(flexdpecom4_4_io_i_data_bus_3),
    .io_i_data_bus2_0(flexdpecom4_4_io_i_data_bus2_0),
    .io_i_data_bus2_1(flexdpecom4_4_io_i_data_bus2_1),
    .io_i_data_bus2_2(flexdpecom4_4_io_i_data_bus2_2),
    .io_i_data_bus2_3(flexdpecom4_4_io_i_data_bus2_3),
    .io_i_vn_0(flexdpecom4_4_io_i_vn_0),
    .io_i_vn_1(flexdpecom4_4_io_i_vn_1),
    .io_i_vn_2(flexdpecom4_4_io_i_vn_2),
    .io_i_vn_3(flexdpecom4_4_io_i_vn_3),
    .io_o_adder_0(flexdpecom4_4_io_o_adder_0),
    .io_o_adder_1(flexdpecom4_4_io_o_adder_1),
    .io_o_adder_2(flexdpecom4_4_io_o_adder_2),
    .io_i_mux_bus_0_0(flexdpecom4_4_io_i_mux_bus_0_0),
    .io_i_mux_bus_0_1(flexdpecom4_4_io_i_mux_bus_0_1),
    .io_i_mux_bus_0_2(flexdpecom4_4_io_i_mux_bus_0_2),
    .io_i_mux_bus_0_3(flexdpecom4_4_io_i_mux_bus_0_3),
    .io_i_mux_bus_1_0(flexdpecom4_4_io_i_mux_bus_1_0),
    .io_i_mux_bus_1_1(flexdpecom4_4_io_i_mux_bus_1_1),
    .io_i_mux_bus_1_2(flexdpecom4_4_io_i_mux_bus_1_2),
    .io_i_mux_bus_2_0(flexdpecom4_4_io_i_mux_bus_2_0),
    .io_i_mux_bus_2_1(flexdpecom4_4_io_i_mux_bus_2_1),
    .io_i_mux_bus_3_0(flexdpecom4_4_io_i_mux_bus_3_0)
  );
  flexdpecom4 flexdpecom4_5 ( // @[FlexDPU.scala 132:47]
    .clock(flexdpecom4_5_clock),
    .reset(flexdpecom4_5_reset),
    .io_i_data_valid(flexdpecom4_5_io_i_data_valid),
    .io_i_data_bus_0(flexdpecom4_5_io_i_data_bus_0),
    .io_i_data_bus_1(flexdpecom4_5_io_i_data_bus_1),
    .io_i_data_bus_2(flexdpecom4_5_io_i_data_bus_2),
    .io_i_data_bus_3(flexdpecom4_5_io_i_data_bus_3),
    .io_i_data_bus2_0(flexdpecom4_5_io_i_data_bus2_0),
    .io_i_data_bus2_1(flexdpecom4_5_io_i_data_bus2_1),
    .io_i_data_bus2_2(flexdpecom4_5_io_i_data_bus2_2),
    .io_i_data_bus2_3(flexdpecom4_5_io_i_data_bus2_3),
    .io_i_vn_0(flexdpecom4_5_io_i_vn_0),
    .io_i_vn_1(flexdpecom4_5_io_i_vn_1),
    .io_i_vn_2(flexdpecom4_5_io_i_vn_2),
    .io_i_vn_3(flexdpecom4_5_io_i_vn_3),
    .io_o_adder_0(flexdpecom4_5_io_o_adder_0),
    .io_o_adder_1(flexdpecom4_5_io_o_adder_1),
    .io_o_adder_2(flexdpecom4_5_io_o_adder_2),
    .io_i_mux_bus_0_0(flexdpecom4_5_io_i_mux_bus_0_0),
    .io_i_mux_bus_0_1(flexdpecom4_5_io_i_mux_bus_0_1),
    .io_i_mux_bus_0_2(flexdpecom4_5_io_i_mux_bus_0_2),
    .io_i_mux_bus_0_3(flexdpecom4_5_io_i_mux_bus_0_3),
    .io_i_mux_bus_1_0(flexdpecom4_5_io_i_mux_bus_1_0),
    .io_i_mux_bus_1_1(flexdpecom4_5_io_i_mux_bus_1_1),
    .io_i_mux_bus_1_2(flexdpecom4_5_io_i_mux_bus_1_2),
    .io_i_mux_bus_2_0(flexdpecom4_5_io_i_mux_bus_2_0),
    .io_i_mux_bus_2_1(flexdpecom4_5_io_i_mux_bus_2_1),
    .io_i_mux_bus_3_0(flexdpecom4_5_io_i_mux_bus_3_0)
  );
  flexdpecom4 flexdpecom4_6 ( // @[FlexDPU.scala 132:47]
    .clock(flexdpecom4_6_clock),
    .reset(flexdpecom4_6_reset),
    .io_i_data_valid(flexdpecom4_6_io_i_data_valid),
    .io_i_data_bus_0(flexdpecom4_6_io_i_data_bus_0),
    .io_i_data_bus_1(flexdpecom4_6_io_i_data_bus_1),
    .io_i_data_bus_2(flexdpecom4_6_io_i_data_bus_2),
    .io_i_data_bus_3(flexdpecom4_6_io_i_data_bus_3),
    .io_i_data_bus2_0(flexdpecom4_6_io_i_data_bus2_0),
    .io_i_data_bus2_1(flexdpecom4_6_io_i_data_bus2_1),
    .io_i_data_bus2_2(flexdpecom4_6_io_i_data_bus2_2),
    .io_i_data_bus2_3(flexdpecom4_6_io_i_data_bus2_3),
    .io_i_vn_0(flexdpecom4_6_io_i_vn_0),
    .io_i_vn_1(flexdpecom4_6_io_i_vn_1),
    .io_i_vn_2(flexdpecom4_6_io_i_vn_2),
    .io_i_vn_3(flexdpecom4_6_io_i_vn_3),
    .io_o_adder_0(flexdpecom4_6_io_o_adder_0),
    .io_o_adder_1(flexdpecom4_6_io_o_adder_1),
    .io_o_adder_2(flexdpecom4_6_io_o_adder_2),
    .io_i_mux_bus_0_0(flexdpecom4_6_io_i_mux_bus_0_0),
    .io_i_mux_bus_0_1(flexdpecom4_6_io_i_mux_bus_0_1),
    .io_i_mux_bus_0_2(flexdpecom4_6_io_i_mux_bus_0_2),
    .io_i_mux_bus_0_3(flexdpecom4_6_io_i_mux_bus_0_3),
    .io_i_mux_bus_1_0(flexdpecom4_6_io_i_mux_bus_1_0),
    .io_i_mux_bus_1_1(flexdpecom4_6_io_i_mux_bus_1_1),
    .io_i_mux_bus_1_2(flexdpecom4_6_io_i_mux_bus_1_2),
    .io_i_mux_bus_2_0(flexdpecom4_6_io_i_mux_bus_2_0),
    .io_i_mux_bus_2_1(flexdpecom4_6_io_i_mux_bus_2_1),
    .io_i_mux_bus_3_0(flexdpecom4_6_io_i_mux_bus_3_0)
  );
  flexdpecom4 flexdpecom4_7 ( // @[FlexDPU.scala 132:47]
    .clock(flexdpecom4_7_clock),
    .reset(flexdpecom4_7_reset),
    .io_i_data_valid(flexdpecom4_7_io_i_data_valid),
    .io_i_data_bus_0(flexdpecom4_7_io_i_data_bus_0),
    .io_i_data_bus_1(flexdpecom4_7_io_i_data_bus_1),
    .io_i_data_bus_2(flexdpecom4_7_io_i_data_bus_2),
    .io_i_data_bus_3(flexdpecom4_7_io_i_data_bus_3),
    .io_i_data_bus2_0(flexdpecom4_7_io_i_data_bus2_0),
    .io_i_data_bus2_1(flexdpecom4_7_io_i_data_bus2_1),
    .io_i_data_bus2_2(flexdpecom4_7_io_i_data_bus2_2),
    .io_i_data_bus2_3(flexdpecom4_7_io_i_data_bus2_3),
    .io_i_vn_0(flexdpecom4_7_io_i_vn_0),
    .io_i_vn_1(flexdpecom4_7_io_i_vn_1),
    .io_i_vn_2(flexdpecom4_7_io_i_vn_2),
    .io_i_vn_3(flexdpecom4_7_io_i_vn_3),
    .io_o_adder_0(flexdpecom4_7_io_o_adder_0),
    .io_o_adder_1(flexdpecom4_7_io_o_adder_1),
    .io_o_adder_2(flexdpecom4_7_io_o_adder_2),
    .io_i_mux_bus_0_0(flexdpecom4_7_io_i_mux_bus_0_0),
    .io_i_mux_bus_0_1(flexdpecom4_7_io_i_mux_bus_0_1),
    .io_i_mux_bus_0_2(flexdpecom4_7_io_i_mux_bus_0_2),
    .io_i_mux_bus_0_3(flexdpecom4_7_io_i_mux_bus_0_3),
    .io_i_mux_bus_1_0(flexdpecom4_7_io_i_mux_bus_1_0),
    .io_i_mux_bus_1_1(flexdpecom4_7_io_i_mux_bus_1_1),
    .io_i_mux_bus_1_2(flexdpecom4_7_io_i_mux_bus_1_2),
    .io_i_mux_bus_2_0(flexdpecom4_7_io_i_mux_bus_2_0),
    .io_i_mux_bus_2_1(flexdpecom4_7_io_i_mux_bus_2_1),
    .io_i_mux_bus_3_0(flexdpecom4_7_io_i_mux_bus_3_0)
  );
  flexdpecom4 flexdpecom4_8 ( // @[FlexDPU.scala 132:47]
    .clock(flexdpecom4_8_clock),
    .reset(flexdpecom4_8_reset),
    .io_i_data_valid(flexdpecom4_8_io_i_data_valid),
    .io_i_data_bus_0(flexdpecom4_8_io_i_data_bus_0),
    .io_i_data_bus_1(flexdpecom4_8_io_i_data_bus_1),
    .io_i_data_bus_2(flexdpecom4_8_io_i_data_bus_2),
    .io_i_data_bus_3(flexdpecom4_8_io_i_data_bus_3),
    .io_i_data_bus2_0(flexdpecom4_8_io_i_data_bus2_0),
    .io_i_data_bus2_1(flexdpecom4_8_io_i_data_bus2_1),
    .io_i_data_bus2_2(flexdpecom4_8_io_i_data_bus2_2),
    .io_i_data_bus2_3(flexdpecom4_8_io_i_data_bus2_3),
    .io_i_vn_0(flexdpecom4_8_io_i_vn_0),
    .io_i_vn_1(flexdpecom4_8_io_i_vn_1),
    .io_i_vn_2(flexdpecom4_8_io_i_vn_2),
    .io_i_vn_3(flexdpecom4_8_io_i_vn_3),
    .io_o_adder_0(flexdpecom4_8_io_o_adder_0),
    .io_o_adder_1(flexdpecom4_8_io_o_adder_1),
    .io_o_adder_2(flexdpecom4_8_io_o_adder_2),
    .io_i_mux_bus_0_0(flexdpecom4_8_io_i_mux_bus_0_0),
    .io_i_mux_bus_0_1(flexdpecom4_8_io_i_mux_bus_0_1),
    .io_i_mux_bus_0_2(flexdpecom4_8_io_i_mux_bus_0_2),
    .io_i_mux_bus_0_3(flexdpecom4_8_io_i_mux_bus_0_3),
    .io_i_mux_bus_1_0(flexdpecom4_8_io_i_mux_bus_1_0),
    .io_i_mux_bus_1_1(flexdpecom4_8_io_i_mux_bus_1_1),
    .io_i_mux_bus_1_2(flexdpecom4_8_io_i_mux_bus_1_2),
    .io_i_mux_bus_2_0(flexdpecom4_8_io_i_mux_bus_2_0),
    .io_i_mux_bus_2_1(flexdpecom4_8_io_i_mux_bus_2_1),
    .io_i_mux_bus_3_0(flexdpecom4_8_io_i_mux_bus_3_0)
  );
  flexdpecom4 flexdpecom4_9 ( // @[FlexDPU.scala 132:47]
    .clock(flexdpecom4_9_clock),
    .reset(flexdpecom4_9_reset),
    .io_i_data_valid(flexdpecom4_9_io_i_data_valid),
    .io_i_data_bus_0(flexdpecom4_9_io_i_data_bus_0),
    .io_i_data_bus_1(flexdpecom4_9_io_i_data_bus_1),
    .io_i_data_bus_2(flexdpecom4_9_io_i_data_bus_2),
    .io_i_data_bus_3(flexdpecom4_9_io_i_data_bus_3),
    .io_i_data_bus2_0(flexdpecom4_9_io_i_data_bus2_0),
    .io_i_data_bus2_1(flexdpecom4_9_io_i_data_bus2_1),
    .io_i_data_bus2_2(flexdpecom4_9_io_i_data_bus2_2),
    .io_i_data_bus2_3(flexdpecom4_9_io_i_data_bus2_3),
    .io_i_vn_0(flexdpecom4_9_io_i_vn_0),
    .io_i_vn_1(flexdpecom4_9_io_i_vn_1),
    .io_i_vn_2(flexdpecom4_9_io_i_vn_2),
    .io_i_vn_3(flexdpecom4_9_io_i_vn_3),
    .io_o_adder_0(flexdpecom4_9_io_o_adder_0),
    .io_o_adder_1(flexdpecom4_9_io_o_adder_1),
    .io_o_adder_2(flexdpecom4_9_io_o_adder_2),
    .io_i_mux_bus_0_0(flexdpecom4_9_io_i_mux_bus_0_0),
    .io_i_mux_bus_0_1(flexdpecom4_9_io_i_mux_bus_0_1),
    .io_i_mux_bus_0_2(flexdpecom4_9_io_i_mux_bus_0_2),
    .io_i_mux_bus_0_3(flexdpecom4_9_io_i_mux_bus_0_3),
    .io_i_mux_bus_1_0(flexdpecom4_9_io_i_mux_bus_1_0),
    .io_i_mux_bus_1_1(flexdpecom4_9_io_i_mux_bus_1_1),
    .io_i_mux_bus_1_2(flexdpecom4_9_io_i_mux_bus_1_2),
    .io_i_mux_bus_2_0(flexdpecom4_9_io_i_mux_bus_2_0),
    .io_i_mux_bus_2_1(flexdpecom4_9_io_i_mux_bus_2_1),
    .io_i_mux_bus_3_0(flexdpecom4_9_io_i_mux_bus_3_0)
  );
  flexdpecom4 flexdpecom4_10 ( // @[FlexDPU.scala 132:47]
    .clock(flexdpecom4_10_clock),
    .reset(flexdpecom4_10_reset),
    .io_i_data_valid(flexdpecom4_10_io_i_data_valid),
    .io_i_data_bus_0(flexdpecom4_10_io_i_data_bus_0),
    .io_i_data_bus_1(flexdpecom4_10_io_i_data_bus_1),
    .io_i_data_bus_2(flexdpecom4_10_io_i_data_bus_2),
    .io_i_data_bus_3(flexdpecom4_10_io_i_data_bus_3),
    .io_i_data_bus2_0(flexdpecom4_10_io_i_data_bus2_0),
    .io_i_data_bus2_1(flexdpecom4_10_io_i_data_bus2_1),
    .io_i_data_bus2_2(flexdpecom4_10_io_i_data_bus2_2),
    .io_i_data_bus2_3(flexdpecom4_10_io_i_data_bus2_3),
    .io_i_vn_0(flexdpecom4_10_io_i_vn_0),
    .io_i_vn_1(flexdpecom4_10_io_i_vn_1),
    .io_i_vn_2(flexdpecom4_10_io_i_vn_2),
    .io_i_vn_3(flexdpecom4_10_io_i_vn_3),
    .io_o_adder_0(flexdpecom4_10_io_o_adder_0),
    .io_o_adder_1(flexdpecom4_10_io_o_adder_1),
    .io_o_adder_2(flexdpecom4_10_io_o_adder_2),
    .io_i_mux_bus_0_0(flexdpecom4_10_io_i_mux_bus_0_0),
    .io_i_mux_bus_0_1(flexdpecom4_10_io_i_mux_bus_0_1),
    .io_i_mux_bus_0_2(flexdpecom4_10_io_i_mux_bus_0_2),
    .io_i_mux_bus_0_3(flexdpecom4_10_io_i_mux_bus_0_3),
    .io_i_mux_bus_1_0(flexdpecom4_10_io_i_mux_bus_1_0),
    .io_i_mux_bus_1_1(flexdpecom4_10_io_i_mux_bus_1_1),
    .io_i_mux_bus_1_2(flexdpecom4_10_io_i_mux_bus_1_2),
    .io_i_mux_bus_2_0(flexdpecom4_10_io_i_mux_bus_2_0),
    .io_i_mux_bus_2_1(flexdpecom4_10_io_i_mux_bus_2_1),
    .io_i_mux_bus_3_0(flexdpecom4_10_io_i_mux_bus_3_0)
  );
  flexdpecom4 flexdpecom4_11 ( // @[FlexDPU.scala 132:47]
    .clock(flexdpecom4_11_clock),
    .reset(flexdpecom4_11_reset),
    .io_i_data_valid(flexdpecom4_11_io_i_data_valid),
    .io_i_data_bus_0(flexdpecom4_11_io_i_data_bus_0),
    .io_i_data_bus_1(flexdpecom4_11_io_i_data_bus_1),
    .io_i_data_bus_2(flexdpecom4_11_io_i_data_bus_2),
    .io_i_data_bus_3(flexdpecom4_11_io_i_data_bus_3),
    .io_i_data_bus2_0(flexdpecom4_11_io_i_data_bus2_0),
    .io_i_data_bus2_1(flexdpecom4_11_io_i_data_bus2_1),
    .io_i_data_bus2_2(flexdpecom4_11_io_i_data_bus2_2),
    .io_i_data_bus2_3(flexdpecom4_11_io_i_data_bus2_3),
    .io_i_vn_0(flexdpecom4_11_io_i_vn_0),
    .io_i_vn_1(flexdpecom4_11_io_i_vn_1),
    .io_i_vn_2(flexdpecom4_11_io_i_vn_2),
    .io_i_vn_3(flexdpecom4_11_io_i_vn_3),
    .io_o_adder_0(flexdpecom4_11_io_o_adder_0),
    .io_o_adder_1(flexdpecom4_11_io_o_adder_1),
    .io_o_adder_2(flexdpecom4_11_io_o_adder_2),
    .io_i_mux_bus_0_0(flexdpecom4_11_io_i_mux_bus_0_0),
    .io_i_mux_bus_0_1(flexdpecom4_11_io_i_mux_bus_0_1),
    .io_i_mux_bus_0_2(flexdpecom4_11_io_i_mux_bus_0_2),
    .io_i_mux_bus_0_3(flexdpecom4_11_io_i_mux_bus_0_3),
    .io_i_mux_bus_1_0(flexdpecom4_11_io_i_mux_bus_1_0),
    .io_i_mux_bus_1_1(flexdpecom4_11_io_i_mux_bus_1_1),
    .io_i_mux_bus_1_2(flexdpecom4_11_io_i_mux_bus_1_2),
    .io_i_mux_bus_2_0(flexdpecom4_11_io_i_mux_bus_2_0),
    .io_i_mux_bus_2_1(flexdpecom4_11_io_i_mux_bus_2_1),
    .io_i_mux_bus_3_0(flexdpecom4_11_io_i_mux_bus_3_0)
  );
  flexdpecom4 flexdpecom4_12 ( // @[FlexDPU.scala 132:47]
    .clock(flexdpecom4_12_clock),
    .reset(flexdpecom4_12_reset),
    .io_i_data_valid(flexdpecom4_12_io_i_data_valid),
    .io_i_data_bus_0(flexdpecom4_12_io_i_data_bus_0),
    .io_i_data_bus_1(flexdpecom4_12_io_i_data_bus_1),
    .io_i_data_bus_2(flexdpecom4_12_io_i_data_bus_2),
    .io_i_data_bus_3(flexdpecom4_12_io_i_data_bus_3),
    .io_i_data_bus2_0(flexdpecom4_12_io_i_data_bus2_0),
    .io_i_data_bus2_1(flexdpecom4_12_io_i_data_bus2_1),
    .io_i_data_bus2_2(flexdpecom4_12_io_i_data_bus2_2),
    .io_i_data_bus2_3(flexdpecom4_12_io_i_data_bus2_3),
    .io_i_vn_0(flexdpecom4_12_io_i_vn_0),
    .io_i_vn_1(flexdpecom4_12_io_i_vn_1),
    .io_i_vn_2(flexdpecom4_12_io_i_vn_2),
    .io_i_vn_3(flexdpecom4_12_io_i_vn_3),
    .io_o_adder_0(flexdpecom4_12_io_o_adder_0),
    .io_o_adder_1(flexdpecom4_12_io_o_adder_1),
    .io_o_adder_2(flexdpecom4_12_io_o_adder_2),
    .io_i_mux_bus_0_0(flexdpecom4_12_io_i_mux_bus_0_0),
    .io_i_mux_bus_0_1(flexdpecom4_12_io_i_mux_bus_0_1),
    .io_i_mux_bus_0_2(flexdpecom4_12_io_i_mux_bus_0_2),
    .io_i_mux_bus_0_3(flexdpecom4_12_io_i_mux_bus_0_3),
    .io_i_mux_bus_1_0(flexdpecom4_12_io_i_mux_bus_1_0),
    .io_i_mux_bus_1_1(flexdpecom4_12_io_i_mux_bus_1_1),
    .io_i_mux_bus_1_2(flexdpecom4_12_io_i_mux_bus_1_2),
    .io_i_mux_bus_2_0(flexdpecom4_12_io_i_mux_bus_2_0),
    .io_i_mux_bus_2_1(flexdpecom4_12_io_i_mux_bus_2_1),
    .io_i_mux_bus_3_0(flexdpecom4_12_io_i_mux_bus_3_0)
  );
  flexdpecom4 flexdpecom4_13 ( // @[FlexDPU.scala 132:47]
    .clock(flexdpecom4_13_clock),
    .reset(flexdpecom4_13_reset),
    .io_i_data_valid(flexdpecom4_13_io_i_data_valid),
    .io_i_data_bus_0(flexdpecom4_13_io_i_data_bus_0),
    .io_i_data_bus_1(flexdpecom4_13_io_i_data_bus_1),
    .io_i_data_bus_2(flexdpecom4_13_io_i_data_bus_2),
    .io_i_data_bus_3(flexdpecom4_13_io_i_data_bus_3),
    .io_i_data_bus2_0(flexdpecom4_13_io_i_data_bus2_0),
    .io_i_data_bus2_1(flexdpecom4_13_io_i_data_bus2_1),
    .io_i_data_bus2_2(flexdpecom4_13_io_i_data_bus2_2),
    .io_i_data_bus2_3(flexdpecom4_13_io_i_data_bus2_3),
    .io_i_vn_0(flexdpecom4_13_io_i_vn_0),
    .io_i_vn_1(flexdpecom4_13_io_i_vn_1),
    .io_i_vn_2(flexdpecom4_13_io_i_vn_2),
    .io_i_vn_3(flexdpecom4_13_io_i_vn_3),
    .io_o_adder_0(flexdpecom4_13_io_o_adder_0),
    .io_o_adder_1(flexdpecom4_13_io_o_adder_1),
    .io_o_adder_2(flexdpecom4_13_io_o_adder_2),
    .io_i_mux_bus_0_0(flexdpecom4_13_io_i_mux_bus_0_0),
    .io_i_mux_bus_0_1(flexdpecom4_13_io_i_mux_bus_0_1),
    .io_i_mux_bus_0_2(flexdpecom4_13_io_i_mux_bus_0_2),
    .io_i_mux_bus_0_3(flexdpecom4_13_io_i_mux_bus_0_3),
    .io_i_mux_bus_1_0(flexdpecom4_13_io_i_mux_bus_1_0),
    .io_i_mux_bus_1_1(flexdpecom4_13_io_i_mux_bus_1_1),
    .io_i_mux_bus_1_2(flexdpecom4_13_io_i_mux_bus_1_2),
    .io_i_mux_bus_2_0(flexdpecom4_13_io_i_mux_bus_2_0),
    .io_i_mux_bus_2_1(flexdpecom4_13_io_i_mux_bus_2_1),
    .io_i_mux_bus_3_0(flexdpecom4_13_io_i_mux_bus_3_0)
  );
  flexdpecom4 flexdpecom4_14 ( // @[FlexDPU.scala 132:47]
    .clock(flexdpecom4_14_clock),
    .reset(flexdpecom4_14_reset),
    .io_i_data_valid(flexdpecom4_14_io_i_data_valid),
    .io_i_data_bus_0(flexdpecom4_14_io_i_data_bus_0),
    .io_i_data_bus_1(flexdpecom4_14_io_i_data_bus_1),
    .io_i_data_bus_2(flexdpecom4_14_io_i_data_bus_2),
    .io_i_data_bus_3(flexdpecom4_14_io_i_data_bus_3),
    .io_i_data_bus2_0(flexdpecom4_14_io_i_data_bus2_0),
    .io_i_data_bus2_1(flexdpecom4_14_io_i_data_bus2_1),
    .io_i_data_bus2_2(flexdpecom4_14_io_i_data_bus2_2),
    .io_i_data_bus2_3(flexdpecom4_14_io_i_data_bus2_3),
    .io_i_vn_0(flexdpecom4_14_io_i_vn_0),
    .io_i_vn_1(flexdpecom4_14_io_i_vn_1),
    .io_i_vn_2(flexdpecom4_14_io_i_vn_2),
    .io_i_vn_3(flexdpecom4_14_io_i_vn_3),
    .io_o_adder_0(flexdpecom4_14_io_o_adder_0),
    .io_o_adder_1(flexdpecom4_14_io_o_adder_1),
    .io_o_adder_2(flexdpecom4_14_io_o_adder_2),
    .io_i_mux_bus_0_0(flexdpecom4_14_io_i_mux_bus_0_0),
    .io_i_mux_bus_0_1(flexdpecom4_14_io_i_mux_bus_0_1),
    .io_i_mux_bus_0_2(flexdpecom4_14_io_i_mux_bus_0_2),
    .io_i_mux_bus_0_3(flexdpecom4_14_io_i_mux_bus_0_3),
    .io_i_mux_bus_1_0(flexdpecom4_14_io_i_mux_bus_1_0),
    .io_i_mux_bus_1_1(flexdpecom4_14_io_i_mux_bus_1_1),
    .io_i_mux_bus_1_2(flexdpecom4_14_io_i_mux_bus_1_2),
    .io_i_mux_bus_2_0(flexdpecom4_14_io_i_mux_bus_2_0),
    .io_i_mux_bus_2_1(flexdpecom4_14_io_i_mux_bus_2_1),
    .io_i_mux_bus_3_0(flexdpecom4_14_io_i_mux_bus_3_0)
  );
  flexdpecom4 flexdpecom4_15 ( // @[FlexDPU.scala 132:47]
    .clock(flexdpecom4_15_clock),
    .reset(flexdpecom4_15_reset),
    .io_i_data_valid(flexdpecom4_15_io_i_data_valid),
    .io_i_data_bus_0(flexdpecom4_15_io_i_data_bus_0),
    .io_i_data_bus_1(flexdpecom4_15_io_i_data_bus_1),
    .io_i_data_bus_2(flexdpecom4_15_io_i_data_bus_2),
    .io_i_data_bus_3(flexdpecom4_15_io_i_data_bus_3),
    .io_i_data_bus2_0(flexdpecom4_15_io_i_data_bus2_0),
    .io_i_data_bus2_1(flexdpecom4_15_io_i_data_bus2_1),
    .io_i_data_bus2_2(flexdpecom4_15_io_i_data_bus2_2),
    .io_i_data_bus2_3(flexdpecom4_15_io_i_data_bus2_3),
    .io_i_vn_0(flexdpecom4_15_io_i_vn_0),
    .io_i_vn_1(flexdpecom4_15_io_i_vn_1),
    .io_i_vn_2(flexdpecom4_15_io_i_vn_2),
    .io_i_vn_3(flexdpecom4_15_io_i_vn_3),
    .io_o_adder_0(flexdpecom4_15_io_o_adder_0),
    .io_o_adder_1(flexdpecom4_15_io_o_adder_1),
    .io_o_adder_2(flexdpecom4_15_io_o_adder_2),
    .io_i_mux_bus_0_0(flexdpecom4_15_io_i_mux_bus_0_0),
    .io_i_mux_bus_0_1(flexdpecom4_15_io_i_mux_bus_0_1),
    .io_i_mux_bus_0_2(flexdpecom4_15_io_i_mux_bus_0_2),
    .io_i_mux_bus_0_3(flexdpecom4_15_io_i_mux_bus_0_3),
    .io_i_mux_bus_1_0(flexdpecom4_15_io_i_mux_bus_1_0),
    .io_i_mux_bus_1_1(flexdpecom4_15_io_i_mux_bus_1_1),
    .io_i_mux_bus_1_2(flexdpecom4_15_io_i_mux_bus_1_2),
    .io_i_mux_bus_2_0(flexdpecom4_15_io_i_mux_bus_2_0),
    .io_i_mux_bus_2_1(flexdpecom4_15_io_i_mux_bus_2_1),
    .io_i_mux_bus_3_0(flexdpecom4_15_io_i_mux_bus_3_0)
  );
  assign PathFinder_clock = clock;
  assign PathFinder_reset = reset;
  assign PathFinder_io_Stationary_matrix_0_0 = Statvalid & check ? io_Stationary_matrix_0_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_0_1 = Statvalid & check ? io_Stationary_matrix_0_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_0_2 = Statvalid & check ? io_Stationary_matrix_0_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_0_3 = Statvalid & check ? io_Stationary_matrix_0_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_0_4 = Statvalid & check ? io_Stationary_matrix_0_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_0_5 = Statvalid & check ? io_Stationary_matrix_0_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_0_6 = Statvalid & check ? io_Stationary_matrix_0_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_0_7 = Statvalid & check ? io_Stationary_matrix_0_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_1_0 = Statvalid & check ? io_Stationary_matrix_1_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_1_1 = Statvalid & check ? io_Stationary_matrix_1_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_1_2 = Statvalid & check ? io_Stationary_matrix_1_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_1_3 = Statvalid & check ? io_Stationary_matrix_1_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_1_4 = Statvalid & check ? io_Stationary_matrix_1_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_1_5 = Statvalid & check ? io_Stationary_matrix_1_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_1_6 = Statvalid & check ? io_Stationary_matrix_1_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_1_7 = Statvalid & check ? io_Stationary_matrix_1_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_2_0 = Statvalid & check ? io_Stationary_matrix_2_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_2_1 = Statvalid & check ? io_Stationary_matrix_2_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_2_2 = Statvalid & check ? io_Stationary_matrix_2_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_2_3 = Statvalid & check ? io_Stationary_matrix_2_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_2_4 = Statvalid & check ? io_Stationary_matrix_2_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_2_5 = Statvalid & check ? io_Stationary_matrix_2_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_2_6 = Statvalid & check ? io_Stationary_matrix_2_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_2_7 = Statvalid & check ? io_Stationary_matrix_2_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_3_0 = Statvalid & check ? io_Stationary_matrix_3_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_3_1 = Statvalid & check ? io_Stationary_matrix_3_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_3_2 = Statvalid & check ? io_Stationary_matrix_3_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_3_3 = Statvalid & check ? io_Stationary_matrix_3_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_3_4 = Statvalid & check ? io_Stationary_matrix_3_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_3_5 = Statvalid & check ? io_Stationary_matrix_3_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_3_6 = Statvalid & check ? io_Stationary_matrix_3_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_3_7 = Statvalid & check ? io_Stationary_matrix_3_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_4_0 = Statvalid & check ? io_Stationary_matrix_4_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_4_1 = Statvalid & check ? io_Stationary_matrix_4_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_4_2 = Statvalid & check ? io_Stationary_matrix_4_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_4_3 = Statvalid & check ? io_Stationary_matrix_4_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_4_4 = Statvalid & check ? io_Stationary_matrix_4_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_4_5 = Statvalid & check ? io_Stationary_matrix_4_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_4_6 = Statvalid & check ? io_Stationary_matrix_4_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_4_7 = Statvalid & check ? io_Stationary_matrix_4_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_5_0 = Statvalid & check ? io_Stationary_matrix_5_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_5_1 = Statvalid & check ? io_Stationary_matrix_5_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_5_2 = Statvalid & check ? io_Stationary_matrix_5_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_5_3 = Statvalid & check ? io_Stationary_matrix_5_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_5_4 = Statvalid & check ? io_Stationary_matrix_5_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_5_5 = Statvalid & check ? io_Stationary_matrix_5_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_5_6 = Statvalid & check ? io_Stationary_matrix_5_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_5_7 = Statvalid & check ? io_Stationary_matrix_5_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_6_0 = Statvalid & check ? io_Stationary_matrix_6_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_6_1 = Statvalid & check ? io_Stationary_matrix_6_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_6_2 = Statvalid & check ? io_Stationary_matrix_6_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_6_3 = Statvalid & check ? io_Stationary_matrix_6_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_6_4 = Statvalid & check ? io_Stationary_matrix_6_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_6_5 = Statvalid & check ? io_Stationary_matrix_6_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_6_6 = Statvalid & check ? io_Stationary_matrix_6_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_6_7 = Statvalid & check ? io_Stationary_matrix_6_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_7_0 = Statvalid & check ? io_Stationary_matrix_7_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_7_1 = Statvalid & check ? io_Stationary_matrix_7_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_7_2 = Statvalid & check ? io_Stationary_matrix_7_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_7_3 = Statvalid & check ? io_Stationary_matrix_7_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_7_4 = Statvalid & check ? io_Stationary_matrix_7_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_7_5 = Statvalid & check ? io_Stationary_matrix_7_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_7_6 = Statvalid & check ? io_Stationary_matrix_7_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Stationary_matrix_7_7 = Statvalid & check ? io_Stationary_matrix_7_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_io_Streaming_matrix_0 = _GEN_397[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_io_Streaming_matrix_1 = _GEN_398[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_io_Streaming_matrix_2 = _GEN_399[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_io_Streaming_matrix_3 = _GEN_400[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_io_Streaming_matrix_4 = _GEN_401[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_io_Streaming_matrix_5 = _GEN_402[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_io_Streaming_matrix_6 = _GEN_403[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_io_Streaming_matrix_7 = _GEN_404[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_io_NoDPE = 32'h0; // @[FlexDPU.scala 77:21]
  assign PathFinder_io_DataValid = Statvalid & check & Statvalid; // @[FlexDPU.scala 112:29 115:25 81:25]
  assign PathFinder_1_clock = clock;
  assign PathFinder_1_reset = reset;
  assign PathFinder_1_io_Stationary_matrix_0_0 = Statvalid & check ? io_Stationary_matrix_0_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_0_1 = Statvalid & check ? io_Stationary_matrix_0_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_0_2 = Statvalid & check ? io_Stationary_matrix_0_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_0_3 = Statvalid & check ? io_Stationary_matrix_0_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_0_4 = Statvalid & check ? io_Stationary_matrix_0_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_0_5 = Statvalid & check ? io_Stationary_matrix_0_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_0_6 = Statvalid & check ? io_Stationary_matrix_0_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_0_7 = Statvalid & check ? io_Stationary_matrix_0_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_1_0 = Statvalid & check ? io_Stationary_matrix_1_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_1_1 = Statvalid & check ? io_Stationary_matrix_1_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_1_2 = Statvalid & check ? io_Stationary_matrix_1_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_1_3 = Statvalid & check ? io_Stationary_matrix_1_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_1_4 = Statvalid & check ? io_Stationary_matrix_1_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_1_5 = Statvalid & check ? io_Stationary_matrix_1_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_1_6 = Statvalid & check ? io_Stationary_matrix_1_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_1_7 = Statvalid & check ? io_Stationary_matrix_1_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_2_0 = Statvalid & check ? io_Stationary_matrix_2_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_2_1 = Statvalid & check ? io_Stationary_matrix_2_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_2_2 = Statvalid & check ? io_Stationary_matrix_2_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_2_3 = Statvalid & check ? io_Stationary_matrix_2_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_2_4 = Statvalid & check ? io_Stationary_matrix_2_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_2_5 = Statvalid & check ? io_Stationary_matrix_2_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_2_6 = Statvalid & check ? io_Stationary_matrix_2_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_2_7 = Statvalid & check ? io_Stationary_matrix_2_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_3_0 = Statvalid & check ? io_Stationary_matrix_3_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_3_1 = Statvalid & check ? io_Stationary_matrix_3_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_3_2 = Statvalid & check ? io_Stationary_matrix_3_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_3_3 = Statvalid & check ? io_Stationary_matrix_3_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_3_4 = Statvalid & check ? io_Stationary_matrix_3_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_3_5 = Statvalid & check ? io_Stationary_matrix_3_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_3_6 = Statvalid & check ? io_Stationary_matrix_3_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_3_7 = Statvalid & check ? io_Stationary_matrix_3_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_4_0 = Statvalid & check ? io_Stationary_matrix_4_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_4_1 = Statvalid & check ? io_Stationary_matrix_4_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_4_2 = Statvalid & check ? io_Stationary_matrix_4_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_4_3 = Statvalid & check ? io_Stationary_matrix_4_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_4_4 = Statvalid & check ? io_Stationary_matrix_4_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_4_5 = Statvalid & check ? io_Stationary_matrix_4_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_4_6 = Statvalid & check ? io_Stationary_matrix_4_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_4_7 = Statvalid & check ? io_Stationary_matrix_4_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_5_0 = Statvalid & check ? io_Stationary_matrix_5_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_5_1 = Statvalid & check ? io_Stationary_matrix_5_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_5_2 = Statvalid & check ? io_Stationary_matrix_5_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_5_3 = Statvalid & check ? io_Stationary_matrix_5_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_5_4 = Statvalid & check ? io_Stationary_matrix_5_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_5_5 = Statvalid & check ? io_Stationary_matrix_5_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_5_6 = Statvalid & check ? io_Stationary_matrix_5_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_5_7 = Statvalid & check ? io_Stationary_matrix_5_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_6_0 = Statvalid & check ? io_Stationary_matrix_6_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_6_1 = Statvalid & check ? io_Stationary_matrix_6_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_6_2 = Statvalid & check ? io_Stationary_matrix_6_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_6_3 = Statvalid & check ? io_Stationary_matrix_6_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_6_4 = Statvalid & check ? io_Stationary_matrix_6_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_6_5 = Statvalid & check ? io_Stationary_matrix_6_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_6_6 = Statvalid & check ? io_Stationary_matrix_6_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_6_7 = Statvalid & check ? io_Stationary_matrix_6_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_7_0 = Statvalid & check ? io_Stationary_matrix_7_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_7_1 = Statvalid & check ? io_Stationary_matrix_7_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_7_2 = Statvalid & check ? io_Stationary_matrix_7_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_7_3 = Statvalid & check ? io_Stationary_matrix_7_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_7_4 = Statvalid & check ? io_Stationary_matrix_7_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_7_5 = Statvalid & check ? io_Stationary_matrix_7_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_7_6 = Statvalid & check ? io_Stationary_matrix_7_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Stationary_matrix_7_7 = Statvalid & check ? io_Stationary_matrix_7_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_1_io_Streaming_matrix_0 = _GEN_397[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_1_io_Streaming_matrix_1 = _GEN_398[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_1_io_Streaming_matrix_2 = _GEN_399[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_1_io_Streaming_matrix_3 = _GEN_400[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_1_io_Streaming_matrix_4 = _GEN_401[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_1_io_Streaming_matrix_5 = _GEN_402[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_1_io_Streaming_matrix_6 = _GEN_403[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_1_io_Streaming_matrix_7 = _GEN_404[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_1_io_NoDPE = {{31'd0}, _T_14}; // @[FlexDPU.scala 77:21]
  assign PathFinder_1_io_DataValid = Statvalid & check & Statvalid; // @[FlexDPU.scala 112:29 115:25 81:25]
  assign PathFinder_2_clock = clock;
  assign PathFinder_2_reset = reset;
  assign PathFinder_2_io_Stationary_matrix_0_0 = Statvalid & check ? io_Stationary_matrix_0_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_0_1 = Statvalid & check ? io_Stationary_matrix_0_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_0_2 = Statvalid & check ? io_Stationary_matrix_0_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_0_3 = Statvalid & check ? io_Stationary_matrix_0_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_0_4 = Statvalid & check ? io_Stationary_matrix_0_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_0_5 = Statvalid & check ? io_Stationary_matrix_0_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_0_6 = Statvalid & check ? io_Stationary_matrix_0_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_0_7 = Statvalid & check ? io_Stationary_matrix_0_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_1_0 = Statvalid & check ? io_Stationary_matrix_1_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_1_1 = Statvalid & check ? io_Stationary_matrix_1_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_1_2 = Statvalid & check ? io_Stationary_matrix_1_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_1_3 = Statvalid & check ? io_Stationary_matrix_1_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_1_4 = Statvalid & check ? io_Stationary_matrix_1_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_1_5 = Statvalid & check ? io_Stationary_matrix_1_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_1_6 = Statvalid & check ? io_Stationary_matrix_1_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_1_7 = Statvalid & check ? io_Stationary_matrix_1_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_2_0 = Statvalid & check ? io_Stationary_matrix_2_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_2_1 = Statvalid & check ? io_Stationary_matrix_2_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_2_2 = Statvalid & check ? io_Stationary_matrix_2_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_2_3 = Statvalid & check ? io_Stationary_matrix_2_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_2_4 = Statvalid & check ? io_Stationary_matrix_2_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_2_5 = Statvalid & check ? io_Stationary_matrix_2_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_2_6 = Statvalid & check ? io_Stationary_matrix_2_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_2_7 = Statvalid & check ? io_Stationary_matrix_2_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_3_0 = Statvalid & check ? io_Stationary_matrix_3_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_3_1 = Statvalid & check ? io_Stationary_matrix_3_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_3_2 = Statvalid & check ? io_Stationary_matrix_3_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_3_3 = Statvalid & check ? io_Stationary_matrix_3_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_3_4 = Statvalid & check ? io_Stationary_matrix_3_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_3_5 = Statvalid & check ? io_Stationary_matrix_3_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_3_6 = Statvalid & check ? io_Stationary_matrix_3_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_3_7 = Statvalid & check ? io_Stationary_matrix_3_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_4_0 = Statvalid & check ? io_Stationary_matrix_4_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_4_1 = Statvalid & check ? io_Stationary_matrix_4_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_4_2 = Statvalid & check ? io_Stationary_matrix_4_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_4_3 = Statvalid & check ? io_Stationary_matrix_4_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_4_4 = Statvalid & check ? io_Stationary_matrix_4_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_4_5 = Statvalid & check ? io_Stationary_matrix_4_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_4_6 = Statvalid & check ? io_Stationary_matrix_4_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_4_7 = Statvalid & check ? io_Stationary_matrix_4_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_5_0 = Statvalid & check ? io_Stationary_matrix_5_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_5_1 = Statvalid & check ? io_Stationary_matrix_5_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_5_2 = Statvalid & check ? io_Stationary_matrix_5_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_5_3 = Statvalid & check ? io_Stationary_matrix_5_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_5_4 = Statvalid & check ? io_Stationary_matrix_5_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_5_5 = Statvalid & check ? io_Stationary_matrix_5_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_5_6 = Statvalid & check ? io_Stationary_matrix_5_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_5_7 = Statvalid & check ? io_Stationary_matrix_5_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_6_0 = Statvalid & check ? io_Stationary_matrix_6_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_6_1 = Statvalid & check ? io_Stationary_matrix_6_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_6_2 = Statvalid & check ? io_Stationary_matrix_6_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_6_3 = Statvalid & check ? io_Stationary_matrix_6_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_6_4 = Statvalid & check ? io_Stationary_matrix_6_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_6_5 = Statvalid & check ? io_Stationary_matrix_6_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_6_6 = Statvalid & check ? io_Stationary_matrix_6_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_6_7 = Statvalid & check ? io_Stationary_matrix_6_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_7_0 = Statvalid & check ? io_Stationary_matrix_7_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_7_1 = Statvalid & check ? io_Stationary_matrix_7_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_7_2 = Statvalid & check ? io_Stationary_matrix_7_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_7_3 = Statvalid & check ? io_Stationary_matrix_7_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_7_4 = Statvalid & check ? io_Stationary_matrix_7_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_7_5 = Statvalid & check ? io_Stationary_matrix_7_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_7_6 = Statvalid & check ? io_Stationary_matrix_7_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Stationary_matrix_7_7 = Statvalid & check ? io_Stationary_matrix_7_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_2_io_Streaming_matrix_0 = _GEN_397[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_2_io_Streaming_matrix_1 = _GEN_398[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_2_io_Streaming_matrix_2 = _GEN_399[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_2_io_Streaming_matrix_3 = _GEN_400[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_2_io_Streaming_matrix_4 = _GEN_401[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_2_io_Streaming_matrix_5 = _GEN_402[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_2_io_Streaming_matrix_6 = _GEN_403[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_2_io_Streaming_matrix_7 = _GEN_404[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_2_io_NoDPE = {{30'd0}, _GEN_554}; // @[FlexDPU.scala 77:21]
  assign PathFinder_2_io_DataValid = Statvalid & check & Statvalid; // @[FlexDPU.scala 112:29 115:25 81:25]
  assign PathFinder_3_clock = clock;
  assign PathFinder_3_reset = reset;
  assign PathFinder_3_io_Stationary_matrix_0_0 = Statvalid & check ? io_Stationary_matrix_0_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_0_1 = Statvalid & check ? io_Stationary_matrix_0_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_0_2 = Statvalid & check ? io_Stationary_matrix_0_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_0_3 = Statvalid & check ? io_Stationary_matrix_0_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_0_4 = Statvalid & check ? io_Stationary_matrix_0_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_0_5 = Statvalid & check ? io_Stationary_matrix_0_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_0_6 = Statvalid & check ? io_Stationary_matrix_0_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_0_7 = Statvalid & check ? io_Stationary_matrix_0_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_1_0 = Statvalid & check ? io_Stationary_matrix_1_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_1_1 = Statvalid & check ? io_Stationary_matrix_1_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_1_2 = Statvalid & check ? io_Stationary_matrix_1_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_1_3 = Statvalid & check ? io_Stationary_matrix_1_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_1_4 = Statvalid & check ? io_Stationary_matrix_1_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_1_5 = Statvalid & check ? io_Stationary_matrix_1_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_1_6 = Statvalid & check ? io_Stationary_matrix_1_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_1_7 = Statvalid & check ? io_Stationary_matrix_1_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_2_0 = Statvalid & check ? io_Stationary_matrix_2_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_2_1 = Statvalid & check ? io_Stationary_matrix_2_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_2_2 = Statvalid & check ? io_Stationary_matrix_2_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_2_3 = Statvalid & check ? io_Stationary_matrix_2_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_2_4 = Statvalid & check ? io_Stationary_matrix_2_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_2_5 = Statvalid & check ? io_Stationary_matrix_2_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_2_6 = Statvalid & check ? io_Stationary_matrix_2_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_2_7 = Statvalid & check ? io_Stationary_matrix_2_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_3_0 = Statvalid & check ? io_Stationary_matrix_3_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_3_1 = Statvalid & check ? io_Stationary_matrix_3_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_3_2 = Statvalid & check ? io_Stationary_matrix_3_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_3_3 = Statvalid & check ? io_Stationary_matrix_3_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_3_4 = Statvalid & check ? io_Stationary_matrix_3_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_3_5 = Statvalid & check ? io_Stationary_matrix_3_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_3_6 = Statvalid & check ? io_Stationary_matrix_3_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_3_7 = Statvalid & check ? io_Stationary_matrix_3_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_4_0 = Statvalid & check ? io_Stationary_matrix_4_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_4_1 = Statvalid & check ? io_Stationary_matrix_4_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_4_2 = Statvalid & check ? io_Stationary_matrix_4_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_4_3 = Statvalid & check ? io_Stationary_matrix_4_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_4_4 = Statvalid & check ? io_Stationary_matrix_4_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_4_5 = Statvalid & check ? io_Stationary_matrix_4_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_4_6 = Statvalid & check ? io_Stationary_matrix_4_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_4_7 = Statvalid & check ? io_Stationary_matrix_4_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_5_0 = Statvalid & check ? io_Stationary_matrix_5_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_5_1 = Statvalid & check ? io_Stationary_matrix_5_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_5_2 = Statvalid & check ? io_Stationary_matrix_5_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_5_3 = Statvalid & check ? io_Stationary_matrix_5_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_5_4 = Statvalid & check ? io_Stationary_matrix_5_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_5_5 = Statvalid & check ? io_Stationary_matrix_5_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_5_6 = Statvalid & check ? io_Stationary_matrix_5_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_5_7 = Statvalid & check ? io_Stationary_matrix_5_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_6_0 = Statvalid & check ? io_Stationary_matrix_6_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_6_1 = Statvalid & check ? io_Stationary_matrix_6_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_6_2 = Statvalid & check ? io_Stationary_matrix_6_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_6_3 = Statvalid & check ? io_Stationary_matrix_6_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_6_4 = Statvalid & check ? io_Stationary_matrix_6_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_6_5 = Statvalid & check ? io_Stationary_matrix_6_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_6_6 = Statvalid & check ? io_Stationary_matrix_6_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_6_7 = Statvalid & check ? io_Stationary_matrix_6_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_7_0 = Statvalid & check ? io_Stationary_matrix_7_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_7_1 = Statvalid & check ? io_Stationary_matrix_7_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_7_2 = Statvalid & check ? io_Stationary_matrix_7_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_7_3 = Statvalid & check ? io_Stationary_matrix_7_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_7_4 = Statvalid & check ? io_Stationary_matrix_7_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_7_5 = Statvalid & check ? io_Stationary_matrix_7_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_7_6 = Statvalid & check ? io_Stationary_matrix_7_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Stationary_matrix_7_7 = Statvalid & check ? io_Stationary_matrix_7_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_3_io_Streaming_matrix_0 = _GEN_397[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_3_io_Streaming_matrix_1 = _GEN_398[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_3_io_Streaming_matrix_2 = _GEN_399[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_3_io_Streaming_matrix_3 = _GEN_400[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_3_io_Streaming_matrix_4 = _GEN_401[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_3_io_Streaming_matrix_5 = _GEN_402[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_3_io_Streaming_matrix_6 = _GEN_403[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_3_io_Streaming_matrix_7 = _GEN_404[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_3_io_NoDPE = {{30'd0}, _GEN_627}; // @[FlexDPU.scala 77:21]
  assign PathFinder_3_io_DataValid = Statvalid & check & Statvalid; // @[FlexDPU.scala 112:29 115:25 81:25]
  assign PathFinder_4_clock = clock;
  assign PathFinder_4_reset = reset;
  assign PathFinder_4_io_Stationary_matrix_0_0 = Statvalid & check ? io_Stationary_matrix_0_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_0_1 = Statvalid & check ? io_Stationary_matrix_0_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_0_2 = Statvalid & check ? io_Stationary_matrix_0_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_0_3 = Statvalid & check ? io_Stationary_matrix_0_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_0_4 = Statvalid & check ? io_Stationary_matrix_0_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_0_5 = Statvalid & check ? io_Stationary_matrix_0_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_0_6 = Statvalid & check ? io_Stationary_matrix_0_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_0_7 = Statvalid & check ? io_Stationary_matrix_0_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_1_0 = Statvalid & check ? io_Stationary_matrix_1_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_1_1 = Statvalid & check ? io_Stationary_matrix_1_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_1_2 = Statvalid & check ? io_Stationary_matrix_1_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_1_3 = Statvalid & check ? io_Stationary_matrix_1_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_1_4 = Statvalid & check ? io_Stationary_matrix_1_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_1_5 = Statvalid & check ? io_Stationary_matrix_1_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_1_6 = Statvalid & check ? io_Stationary_matrix_1_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_1_7 = Statvalid & check ? io_Stationary_matrix_1_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_2_0 = Statvalid & check ? io_Stationary_matrix_2_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_2_1 = Statvalid & check ? io_Stationary_matrix_2_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_2_2 = Statvalid & check ? io_Stationary_matrix_2_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_2_3 = Statvalid & check ? io_Stationary_matrix_2_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_2_4 = Statvalid & check ? io_Stationary_matrix_2_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_2_5 = Statvalid & check ? io_Stationary_matrix_2_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_2_6 = Statvalid & check ? io_Stationary_matrix_2_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_2_7 = Statvalid & check ? io_Stationary_matrix_2_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_3_0 = Statvalid & check ? io_Stationary_matrix_3_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_3_1 = Statvalid & check ? io_Stationary_matrix_3_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_3_2 = Statvalid & check ? io_Stationary_matrix_3_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_3_3 = Statvalid & check ? io_Stationary_matrix_3_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_3_4 = Statvalid & check ? io_Stationary_matrix_3_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_3_5 = Statvalid & check ? io_Stationary_matrix_3_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_3_6 = Statvalid & check ? io_Stationary_matrix_3_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_3_7 = Statvalid & check ? io_Stationary_matrix_3_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_4_0 = Statvalid & check ? io_Stationary_matrix_4_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_4_1 = Statvalid & check ? io_Stationary_matrix_4_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_4_2 = Statvalid & check ? io_Stationary_matrix_4_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_4_3 = Statvalid & check ? io_Stationary_matrix_4_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_4_4 = Statvalid & check ? io_Stationary_matrix_4_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_4_5 = Statvalid & check ? io_Stationary_matrix_4_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_4_6 = Statvalid & check ? io_Stationary_matrix_4_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_4_7 = Statvalid & check ? io_Stationary_matrix_4_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_5_0 = Statvalid & check ? io_Stationary_matrix_5_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_5_1 = Statvalid & check ? io_Stationary_matrix_5_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_5_2 = Statvalid & check ? io_Stationary_matrix_5_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_5_3 = Statvalid & check ? io_Stationary_matrix_5_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_5_4 = Statvalid & check ? io_Stationary_matrix_5_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_5_5 = Statvalid & check ? io_Stationary_matrix_5_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_5_6 = Statvalid & check ? io_Stationary_matrix_5_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_5_7 = Statvalid & check ? io_Stationary_matrix_5_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_6_0 = Statvalid & check ? io_Stationary_matrix_6_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_6_1 = Statvalid & check ? io_Stationary_matrix_6_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_6_2 = Statvalid & check ? io_Stationary_matrix_6_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_6_3 = Statvalid & check ? io_Stationary_matrix_6_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_6_4 = Statvalid & check ? io_Stationary_matrix_6_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_6_5 = Statvalid & check ? io_Stationary_matrix_6_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_6_6 = Statvalid & check ? io_Stationary_matrix_6_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_6_7 = Statvalid & check ? io_Stationary_matrix_6_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_7_0 = Statvalid & check ? io_Stationary_matrix_7_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_7_1 = Statvalid & check ? io_Stationary_matrix_7_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_7_2 = Statvalid & check ? io_Stationary_matrix_7_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_7_3 = Statvalid & check ? io_Stationary_matrix_7_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_7_4 = Statvalid & check ? io_Stationary_matrix_7_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_7_5 = Statvalid & check ? io_Stationary_matrix_7_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_7_6 = Statvalid & check ? io_Stationary_matrix_7_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Stationary_matrix_7_7 = Statvalid & check ? io_Stationary_matrix_7_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_4_io_Streaming_matrix_0 = _GEN_397[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_4_io_Streaming_matrix_1 = _GEN_398[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_4_io_Streaming_matrix_2 = _GEN_399[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_4_io_Streaming_matrix_3 = _GEN_400[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_4_io_Streaming_matrix_4 = _GEN_401[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_4_io_Streaming_matrix_5 = _GEN_402[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_4_io_Streaming_matrix_6 = _GEN_403[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_4_io_Streaming_matrix_7 = _GEN_404[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_4_io_NoDPE = {{29'd0}, _GEN_700}; // @[FlexDPU.scala 77:21]
  assign PathFinder_4_io_DataValid = Statvalid & check & Statvalid; // @[FlexDPU.scala 112:29 115:25 81:25]
  assign PathFinder_5_clock = clock;
  assign PathFinder_5_reset = reset;
  assign PathFinder_5_io_Stationary_matrix_0_0 = Statvalid & check ? io_Stationary_matrix_0_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_0_1 = Statvalid & check ? io_Stationary_matrix_0_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_0_2 = Statvalid & check ? io_Stationary_matrix_0_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_0_3 = Statvalid & check ? io_Stationary_matrix_0_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_0_4 = Statvalid & check ? io_Stationary_matrix_0_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_0_5 = Statvalid & check ? io_Stationary_matrix_0_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_0_6 = Statvalid & check ? io_Stationary_matrix_0_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_0_7 = Statvalid & check ? io_Stationary_matrix_0_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_1_0 = Statvalid & check ? io_Stationary_matrix_1_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_1_1 = Statvalid & check ? io_Stationary_matrix_1_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_1_2 = Statvalid & check ? io_Stationary_matrix_1_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_1_3 = Statvalid & check ? io_Stationary_matrix_1_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_1_4 = Statvalid & check ? io_Stationary_matrix_1_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_1_5 = Statvalid & check ? io_Stationary_matrix_1_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_1_6 = Statvalid & check ? io_Stationary_matrix_1_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_1_7 = Statvalid & check ? io_Stationary_matrix_1_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_2_0 = Statvalid & check ? io_Stationary_matrix_2_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_2_1 = Statvalid & check ? io_Stationary_matrix_2_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_2_2 = Statvalid & check ? io_Stationary_matrix_2_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_2_3 = Statvalid & check ? io_Stationary_matrix_2_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_2_4 = Statvalid & check ? io_Stationary_matrix_2_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_2_5 = Statvalid & check ? io_Stationary_matrix_2_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_2_6 = Statvalid & check ? io_Stationary_matrix_2_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_2_7 = Statvalid & check ? io_Stationary_matrix_2_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_3_0 = Statvalid & check ? io_Stationary_matrix_3_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_3_1 = Statvalid & check ? io_Stationary_matrix_3_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_3_2 = Statvalid & check ? io_Stationary_matrix_3_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_3_3 = Statvalid & check ? io_Stationary_matrix_3_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_3_4 = Statvalid & check ? io_Stationary_matrix_3_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_3_5 = Statvalid & check ? io_Stationary_matrix_3_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_3_6 = Statvalid & check ? io_Stationary_matrix_3_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_3_7 = Statvalid & check ? io_Stationary_matrix_3_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_4_0 = Statvalid & check ? io_Stationary_matrix_4_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_4_1 = Statvalid & check ? io_Stationary_matrix_4_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_4_2 = Statvalid & check ? io_Stationary_matrix_4_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_4_3 = Statvalid & check ? io_Stationary_matrix_4_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_4_4 = Statvalid & check ? io_Stationary_matrix_4_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_4_5 = Statvalid & check ? io_Stationary_matrix_4_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_4_6 = Statvalid & check ? io_Stationary_matrix_4_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_4_7 = Statvalid & check ? io_Stationary_matrix_4_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_5_0 = Statvalid & check ? io_Stationary_matrix_5_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_5_1 = Statvalid & check ? io_Stationary_matrix_5_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_5_2 = Statvalid & check ? io_Stationary_matrix_5_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_5_3 = Statvalid & check ? io_Stationary_matrix_5_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_5_4 = Statvalid & check ? io_Stationary_matrix_5_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_5_5 = Statvalid & check ? io_Stationary_matrix_5_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_5_6 = Statvalid & check ? io_Stationary_matrix_5_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_5_7 = Statvalid & check ? io_Stationary_matrix_5_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_6_0 = Statvalid & check ? io_Stationary_matrix_6_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_6_1 = Statvalid & check ? io_Stationary_matrix_6_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_6_2 = Statvalid & check ? io_Stationary_matrix_6_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_6_3 = Statvalid & check ? io_Stationary_matrix_6_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_6_4 = Statvalid & check ? io_Stationary_matrix_6_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_6_5 = Statvalid & check ? io_Stationary_matrix_6_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_6_6 = Statvalid & check ? io_Stationary_matrix_6_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_6_7 = Statvalid & check ? io_Stationary_matrix_6_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_7_0 = Statvalid & check ? io_Stationary_matrix_7_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_7_1 = Statvalid & check ? io_Stationary_matrix_7_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_7_2 = Statvalid & check ? io_Stationary_matrix_7_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_7_3 = Statvalid & check ? io_Stationary_matrix_7_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_7_4 = Statvalid & check ? io_Stationary_matrix_7_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_7_5 = Statvalid & check ? io_Stationary_matrix_7_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_7_6 = Statvalid & check ? io_Stationary_matrix_7_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Stationary_matrix_7_7 = Statvalid & check ? io_Stationary_matrix_7_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_5_io_Streaming_matrix_0 = _GEN_397[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_5_io_Streaming_matrix_1 = _GEN_398[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_5_io_Streaming_matrix_2 = _GEN_399[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_5_io_Streaming_matrix_3 = _GEN_400[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_5_io_Streaming_matrix_4 = _GEN_401[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_5_io_Streaming_matrix_5 = _GEN_402[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_5_io_Streaming_matrix_6 = _GEN_403[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_5_io_Streaming_matrix_7 = _GEN_404[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_5_io_NoDPE = {{29'd0}, _GEN_773}; // @[FlexDPU.scala 77:21]
  assign PathFinder_5_io_DataValid = Statvalid & check & Statvalid; // @[FlexDPU.scala 112:29 115:25 81:25]
  assign PathFinder_6_clock = clock;
  assign PathFinder_6_reset = reset;
  assign PathFinder_6_io_Stationary_matrix_0_0 = Statvalid & check ? io_Stationary_matrix_0_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_0_1 = Statvalid & check ? io_Stationary_matrix_0_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_0_2 = Statvalid & check ? io_Stationary_matrix_0_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_0_3 = Statvalid & check ? io_Stationary_matrix_0_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_0_4 = Statvalid & check ? io_Stationary_matrix_0_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_0_5 = Statvalid & check ? io_Stationary_matrix_0_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_0_6 = Statvalid & check ? io_Stationary_matrix_0_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_0_7 = Statvalid & check ? io_Stationary_matrix_0_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_1_0 = Statvalid & check ? io_Stationary_matrix_1_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_1_1 = Statvalid & check ? io_Stationary_matrix_1_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_1_2 = Statvalid & check ? io_Stationary_matrix_1_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_1_3 = Statvalid & check ? io_Stationary_matrix_1_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_1_4 = Statvalid & check ? io_Stationary_matrix_1_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_1_5 = Statvalid & check ? io_Stationary_matrix_1_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_1_6 = Statvalid & check ? io_Stationary_matrix_1_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_1_7 = Statvalid & check ? io_Stationary_matrix_1_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_2_0 = Statvalid & check ? io_Stationary_matrix_2_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_2_1 = Statvalid & check ? io_Stationary_matrix_2_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_2_2 = Statvalid & check ? io_Stationary_matrix_2_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_2_3 = Statvalid & check ? io_Stationary_matrix_2_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_2_4 = Statvalid & check ? io_Stationary_matrix_2_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_2_5 = Statvalid & check ? io_Stationary_matrix_2_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_2_6 = Statvalid & check ? io_Stationary_matrix_2_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_2_7 = Statvalid & check ? io_Stationary_matrix_2_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_3_0 = Statvalid & check ? io_Stationary_matrix_3_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_3_1 = Statvalid & check ? io_Stationary_matrix_3_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_3_2 = Statvalid & check ? io_Stationary_matrix_3_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_3_3 = Statvalid & check ? io_Stationary_matrix_3_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_3_4 = Statvalid & check ? io_Stationary_matrix_3_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_3_5 = Statvalid & check ? io_Stationary_matrix_3_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_3_6 = Statvalid & check ? io_Stationary_matrix_3_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_3_7 = Statvalid & check ? io_Stationary_matrix_3_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_4_0 = Statvalid & check ? io_Stationary_matrix_4_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_4_1 = Statvalid & check ? io_Stationary_matrix_4_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_4_2 = Statvalid & check ? io_Stationary_matrix_4_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_4_3 = Statvalid & check ? io_Stationary_matrix_4_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_4_4 = Statvalid & check ? io_Stationary_matrix_4_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_4_5 = Statvalid & check ? io_Stationary_matrix_4_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_4_6 = Statvalid & check ? io_Stationary_matrix_4_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_4_7 = Statvalid & check ? io_Stationary_matrix_4_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_5_0 = Statvalid & check ? io_Stationary_matrix_5_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_5_1 = Statvalid & check ? io_Stationary_matrix_5_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_5_2 = Statvalid & check ? io_Stationary_matrix_5_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_5_3 = Statvalid & check ? io_Stationary_matrix_5_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_5_4 = Statvalid & check ? io_Stationary_matrix_5_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_5_5 = Statvalid & check ? io_Stationary_matrix_5_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_5_6 = Statvalid & check ? io_Stationary_matrix_5_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_5_7 = Statvalid & check ? io_Stationary_matrix_5_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_6_0 = Statvalid & check ? io_Stationary_matrix_6_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_6_1 = Statvalid & check ? io_Stationary_matrix_6_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_6_2 = Statvalid & check ? io_Stationary_matrix_6_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_6_3 = Statvalid & check ? io_Stationary_matrix_6_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_6_4 = Statvalid & check ? io_Stationary_matrix_6_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_6_5 = Statvalid & check ? io_Stationary_matrix_6_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_6_6 = Statvalid & check ? io_Stationary_matrix_6_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_6_7 = Statvalid & check ? io_Stationary_matrix_6_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_7_0 = Statvalid & check ? io_Stationary_matrix_7_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_7_1 = Statvalid & check ? io_Stationary_matrix_7_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_7_2 = Statvalid & check ? io_Stationary_matrix_7_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_7_3 = Statvalid & check ? io_Stationary_matrix_7_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_7_4 = Statvalid & check ? io_Stationary_matrix_7_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_7_5 = Statvalid & check ? io_Stationary_matrix_7_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_7_6 = Statvalid & check ? io_Stationary_matrix_7_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Stationary_matrix_7_7 = Statvalid & check ? io_Stationary_matrix_7_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_6_io_Streaming_matrix_0 = _GEN_397[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_6_io_Streaming_matrix_1 = _GEN_398[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_6_io_Streaming_matrix_2 = _GEN_399[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_6_io_Streaming_matrix_3 = _GEN_400[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_6_io_Streaming_matrix_4 = _GEN_401[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_6_io_Streaming_matrix_5 = _GEN_402[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_6_io_Streaming_matrix_6 = _GEN_403[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_6_io_Streaming_matrix_7 = _GEN_404[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_6_io_NoDPE = {{29'd0}, _GEN_846}; // @[FlexDPU.scala 77:21]
  assign PathFinder_6_io_DataValid = Statvalid & check & Statvalid; // @[FlexDPU.scala 112:29 115:25 81:25]
  assign PathFinder_7_clock = clock;
  assign PathFinder_7_reset = reset;
  assign PathFinder_7_io_Stationary_matrix_0_0 = Statvalid & check ? io_Stationary_matrix_0_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_0_1 = Statvalid & check ? io_Stationary_matrix_0_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_0_2 = Statvalid & check ? io_Stationary_matrix_0_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_0_3 = Statvalid & check ? io_Stationary_matrix_0_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_0_4 = Statvalid & check ? io_Stationary_matrix_0_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_0_5 = Statvalid & check ? io_Stationary_matrix_0_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_0_6 = Statvalid & check ? io_Stationary_matrix_0_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_0_7 = Statvalid & check ? io_Stationary_matrix_0_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_1_0 = Statvalid & check ? io_Stationary_matrix_1_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_1_1 = Statvalid & check ? io_Stationary_matrix_1_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_1_2 = Statvalid & check ? io_Stationary_matrix_1_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_1_3 = Statvalid & check ? io_Stationary_matrix_1_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_1_4 = Statvalid & check ? io_Stationary_matrix_1_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_1_5 = Statvalid & check ? io_Stationary_matrix_1_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_1_6 = Statvalid & check ? io_Stationary_matrix_1_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_1_7 = Statvalid & check ? io_Stationary_matrix_1_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_2_0 = Statvalid & check ? io_Stationary_matrix_2_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_2_1 = Statvalid & check ? io_Stationary_matrix_2_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_2_2 = Statvalid & check ? io_Stationary_matrix_2_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_2_3 = Statvalid & check ? io_Stationary_matrix_2_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_2_4 = Statvalid & check ? io_Stationary_matrix_2_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_2_5 = Statvalid & check ? io_Stationary_matrix_2_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_2_6 = Statvalid & check ? io_Stationary_matrix_2_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_2_7 = Statvalid & check ? io_Stationary_matrix_2_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_3_0 = Statvalid & check ? io_Stationary_matrix_3_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_3_1 = Statvalid & check ? io_Stationary_matrix_3_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_3_2 = Statvalid & check ? io_Stationary_matrix_3_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_3_3 = Statvalid & check ? io_Stationary_matrix_3_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_3_4 = Statvalid & check ? io_Stationary_matrix_3_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_3_5 = Statvalid & check ? io_Stationary_matrix_3_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_3_6 = Statvalid & check ? io_Stationary_matrix_3_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_3_7 = Statvalid & check ? io_Stationary_matrix_3_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_4_0 = Statvalid & check ? io_Stationary_matrix_4_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_4_1 = Statvalid & check ? io_Stationary_matrix_4_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_4_2 = Statvalid & check ? io_Stationary_matrix_4_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_4_3 = Statvalid & check ? io_Stationary_matrix_4_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_4_4 = Statvalid & check ? io_Stationary_matrix_4_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_4_5 = Statvalid & check ? io_Stationary_matrix_4_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_4_6 = Statvalid & check ? io_Stationary_matrix_4_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_4_7 = Statvalid & check ? io_Stationary_matrix_4_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_5_0 = Statvalid & check ? io_Stationary_matrix_5_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_5_1 = Statvalid & check ? io_Stationary_matrix_5_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_5_2 = Statvalid & check ? io_Stationary_matrix_5_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_5_3 = Statvalid & check ? io_Stationary_matrix_5_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_5_4 = Statvalid & check ? io_Stationary_matrix_5_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_5_5 = Statvalid & check ? io_Stationary_matrix_5_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_5_6 = Statvalid & check ? io_Stationary_matrix_5_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_5_7 = Statvalid & check ? io_Stationary_matrix_5_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_6_0 = Statvalid & check ? io_Stationary_matrix_6_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_6_1 = Statvalid & check ? io_Stationary_matrix_6_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_6_2 = Statvalid & check ? io_Stationary_matrix_6_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_6_3 = Statvalid & check ? io_Stationary_matrix_6_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_6_4 = Statvalid & check ? io_Stationary_matrix_6_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_6_5 = Statvalid & check ? io_Stationary_matrix_6_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_6_6 = Statvalid & check ? io_Stationary_matrix_6_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_6_7 = Statvalid & check ? io_Stationary_matrix_6_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_7_0 = Statvalid & check ? io_Stationary_matrix_7_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_7_1 = Statvalid & check ? io_Stationary_matrix_7_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_7_2 = Statvalid & check ? io_Stationary_matrix_7_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_7_3 = Statvalid & check ? io_Stationary_matrix_7_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_7_4 = Statvalid & check ? io_Stationary_matrix_7_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_7_5 = Statvalid & check ? io_Stationary_matrix_7_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_7_6 = Statvalid & check ? io_Stationary_matrix_7_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Stationary_matrix_7_7 = Statvalid & check ? io_Stationary_matrix_7_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_7_io_Streaming_matrix_0 = _GEN_397[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_7_io_Streaming_matrix_1 = _GEN_398[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_7_io_Streaming_matrix_2 = _GEN_399[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_7_io_Streaming_matrix_3 = _GEN_400[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_7_io_Streaming_matrix_4 = _GEN_401[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_7_io_Streaming_matrix_5 = _GEN_402[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_7_io_Streaming_matrix_6 = _GEN_403[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_7_io_Streaming_matrix_7 = _GEN_404[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_7_io_NoDPE = {{29'd0}, _GEN_919}; // @[FlexDPU.scala 77:21]
  assign PathFinder_7_io_DataValid = Statvalid & check & Statvalid; // @[FlexDPU.scala 112:29 115:25 81:25]
  assign PathFinder_8_clock = clock;
  assign PathFinder_8_reset = reset;
  assign PathFinder_8_io_Stationary_matrix_0_0 = Statvalid & check ? io_Stationary_matrix_0_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_0_1 = Statvalid & check ? io_Stationary_matrix_0_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_0_2 = Statvalid & check ? io_Stationary_matrix_0_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_0_3 = Statvalid & check ? io_Stationary_matrix_0_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_0_4 = Statvalid & check ? io_Stationary_matrix_0_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_0_5 = Statvalid & check ? io_Stationary_matrix_0_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_0_6 = Statvalid & check ? io_Stationary_matrix_0_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_0_7 = Statvalid & check ? io_Stationary_matrix_0_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_1_0 = Statvalid & check ? io_Stationary_matrix_1_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_1_1 = Statvalid & check ? io_Stationary_matrix_1_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_1_2 = Statvalid & check ? io_Stationary_matrix_1_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_1_3 = Statvalid & check ? io_Stationary_matrix_1_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_1_4 = Statvalid & check ? io_Stationary_matrix_1_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_1_5 = Statvalid & check ? io_Stationary_matrix_1_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_1_6 = Statvalid & check ? io_Stationary_matrix_1_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_1_7 = Statvalid & check ? io_Stationary_matrix_1_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_2_0 = Statvalid & check ? io_Stationary_matrix_2_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_2_1 = Statvalid & check ? io_Stationary_matrix_2_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_2_2 = Statvalid & check ? io_Stationary_matrix_2_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_2_3 = Statvalid & check ? io_Stationary_matrix_2_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_2_4 = Statvalid & check ? io_Stationary_matrix_2_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_2_5 = Statvalid & check ? io_Stationary_matrix_2_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_2_6 = Statvalid & check ? io_Stationary_matrix_2_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_2_7 = Statvalid & check ? io_Stationary_matrix_2_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_3_0 = Statvalid & check ? io_Stationary_matrix_3_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_3_1 = Statvalid & check ? io_Stationary_matrix_3_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_3_2 = Statvalid & check ? io_Stationary_matrix_3_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_3_3 = Statvalid & check ? io_Stationary_matrix_3_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_3_4 = Statvalid & check ? io_Stationary_matrix_3_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_3_5 = Statvalid & check ? io_Stationary_matrix_3_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_3_6 = Statvalid & check ? io_Stationary_matrix_3_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_3_7 = Statvalid & check ? io_Stationary_matrix_3_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_4_0 = Statvalid & check ? io_Stationary_matrix_4_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_4_1 = Statvalid & check ? io_Stationary_matrix_4_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_4_2 = Statvalid & check ? io_Stationary_matrix_4_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_4_3 = Statvalid & check ? io_Stationary_matrix_4_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_4_4 = Statvalid & check ? io_Stationary_matrix_4_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_4_5 = Statvalid & check ? io_Stationary_matrix_4_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_4_6 = Statvalid & check ? io_Stationary_matrix_4_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_4_7 = Statvalid & check ? io_Stationary_matrix_4_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_5_0 = Statvalid & check ? io_Stationary_matrix_5_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_5_1 = Statvalid & check ? io_Stationary_matrix_5_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_5_2 = Statvalid & check ? io_Stationary_matrix_5_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_5_3 = Statvalid & check ? io_Stationary_matrix_5_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_5_4 = Statvalid & check ? io_Stationary_matrix_5_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_5_5 = Statvalid & check ? io_Stationary_matrix_5_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_5_6 = Statvalid & check ? io_Stationary_matrix_5_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_5_7 = Statvalid & check ? io_Stationary_matrix_5_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_6_0 = Statvalid & check ? io_Stationary_matrix_6_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_6_1 = Statvalid & check ? io_Stationary_matrix_6_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_6_2 = Statvalid & check ? io_Stationary_matrix_6_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_6_3 = Statvalid & check ? io_Stationary_matrix_6_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_6_4 = Statvalid & check ? io_Stationary_matrix_6_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_6_5 = Statvalid & check ? io_Stationary_matrix_6_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_6_6 = Statvalid & check ? io_Stationary_matrix_6_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_6_7 = Statvalid & check ? io_Stationary_matrix_6_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_7_0 = Statvalid & check ? io_Stationary_matrix_7_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_7_1 = Statvalid & check ? io_Stationary_matrix_7_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_7_2 = Statvalid & check ? io_Stationary_matrix_7_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_7_3 = Statvalid & check ? io_Stationary_matrix_7_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_7_4 = Statvalid & check ? io_Stationary_matrix_7_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_7_5 = Statvalid & check ? io_Stationary_matrix_7_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_7_6 = Statvalid & check ? io_Stationary_matrix_7_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Stationary_matrix_7_7 = Statvalid & check ? io_Stationary_matrix_7_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_8_io_Streaming_matrix_0 = _GEN_397[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_8_io_Streaming_matrix_1 = _GEN_398[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_8_io_Streaming_matrix_2 = _GEN_399[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_8_io_Streaming_matrix_3 = _GEN_400[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_8_io_Streaming_matrix_4 = _GEN_401[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_8_io_Streaming_matrix_5 = _GEN_402[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_8_io_Streaming_matrix_6 = _GEN_403[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_8_io_Streaming_matrix_7 = _GEN_404[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_8_io_NoDPE = {{28'd0}, _GEN_992}; // @[FlexDPU.scala 77:21]
  assign PathFinder_8_io_DataValid = Statvalid & check & Statvalid; // @[FlexDPU.scala 112:29 115:25 81:25]
  assign PathFinder_9_clock = clock;
  assign PathFinder_9_reset = reset;
  assign PathFinder_9_io_Stationary_matrix_0_0 = Statvalid & check ? io_Stationary_matrix_0_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_0_1 = Statvalid & check ? io_Stationary_matrix_0_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_0_2 = Statvalid & check ? io_Stationary_matrix_0_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_0_3 = Statvalid & check ? io_Stationary_matrix_0_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_0_4 = Statvalid & check ? io_Stationary_matrix_0_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_0_5 = Statvalid & check ? io_Stationary_matrix_0_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_0_6 = Statvalid & check ? io_Stationary_matrix_0_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_0_7 = Statvalid & check ? io_Stationary_matrix_0_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_1_0 = Statvalid & check ? io_Stationary_matrix_1_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_1_1 = Statvalid & check ? io_Stationary_matrix_1_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_1_2 = Statvalid & check ? io_Stationary_matrix_1_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_1_3 = Statvalid & check ? io_Stationary_matrix_1_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_1_4 = Statvalid & check ? io_Stationary_matrix_1_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_1_5 = Statvalid & check ? io_Stationary_matrix_1_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_1_6 = Statvalid & check ? io_Stationary_matrix_1_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_1_7 = Statvalid & check ? io_Stationary_matrix_1_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_2_0 = Statvalid & check ? io_Stationary_matrix_2_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_2_1 = Statvalid & check ? io_Stationary_matrix_2_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_2_2 = Statvalid & check ? io_Stationary_matrix_2_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_2_3 = Statvalid & check ? io_Stationary_matrix_2_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_2_4 = Statvalid & check ? io_Stationary_matrix_2_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_2_5 = Statvalid & check ? io_Stationary_matrix_2_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_2_6 = Statvalid & check ? io_Stationary_matrix_2_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_2_7 = Statvalid & check ? io_Stationary_matrix_2_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_3_0 = Statvalid & check ? io_Stationary_matrix_3_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_3_1 = Statvalid & check ? io_Stationary_matrix_3_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_3_2 = Statvalid & check ? io_Stationary_matrix_3_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_3_3 = Statvalid & check ? io_Stationary_matrix_3_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_3_4 = Statvalid & check ? io_Stationary_matrix_3_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_3_5 = Statvalid & check ? io_Stationary_matrix_3_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_3_6 = Statvalid & check ? io_Stationary_matrix_3_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_3_7 = Statvalid & check ? io_Stationary_matrix_3_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_4_0 = Statvalid & check ? io_Stationary_matrix_4_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_4_1 = Statvalid & check ? io_Stationary_matrix_4_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_4_2 = Statvalid & check ? io_Stationary_matrix_4_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_4_3 = Statvalid & check ? io_Stationary_matrix_4_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_4_4 = Statvalid & check ? io_Stationary_matrix_4_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_4_5 = Statvalid & check ? io_Stationary_matrix_4_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_4_6 = Statvalid & check ? io_Stationary_matrix_4_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_4_7 = Statvalid & check ? io_Stationary_matrix_4_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_5_0 = Statvalid & check ? io_Stationary_matrix_5_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_5_1 = Statvalid & check ? io_Stationary_matrix_5_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_5_2 = Statvalid & check ? io_Stationary_matrix_5_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_5_3 = Statvalid & check ? io_Stationary_matrix_5_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_5_4 = Statvalid & check ? io_Stationary_matrix_5_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_5_5 = Statvalid & check ? io_Stationary_matrix_5_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_5_6 = Statvalid & check ? io_Stationary_matrix_5_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_5_7 = Statvalid & check ? io_Stationary_matrix_5_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_6_0 = Statvalid & check ? io_Stationary_matrix_6_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_6_1 = Statvalid & check ? io_Stationary_matrix_6_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_6_2 = Statvalid & check ? io_Stationary_matrix_6_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_6_3 = Statvalid & check ? io_Stationary_matrix_6_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_6_4 = Statvalid & check ? io_Stationary_matrix_6_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_6_5 = Statvalid & check ? io_Stationary_matrix_6_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_6_6 = Statvalid & check ? io_Stationary_matrix_6_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_6_7 = Statvalid & check ? io_Stationary_matrix_6_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_7_0 = Statvalid & check ? io_Stationary_matrix_7_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_7_1 = Statvalid & check ? io_Stationary_matrix_7_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_7_2 = Statvalid & check ? io_Stationary_matrix_7_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_7_3 = Statvalid & check ? io_Stationary_matrix_7_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_7_4 = Statvalid & check ? io_Stationary_matrix_7_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_7_5 = Statvalid & check ? io_Stationary_matrix_7_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_7_6 = Statvalid & check ? io_Stationary_matrix_7_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Stationary_matrix_7_7 = Statvalid & check ? io_Stationary_matrix_7_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_9_io_Streaming_matrix_0 = _GEN_397[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_9_io_Streaming_matrix_1 = _GEN_398[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_9_io_Streaming_matrix_2 = _GEN_399[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_9_io_Streaming_matrix_3 = _GEN_400[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_9_io_Streaming_matrix_4 = _GEN_401[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_9_io_Streaming_matrix_5 = _GEN_402[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_9_io_Streaming_matrix_6 = _GEN_403[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_9_io_Streaming_matrix_7 = _GEN_404[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_9_io_NoDPE = {{28'd0}, _GEN_1065}; // @[FlexDPU.scala 77:21]
  assign PathFinder_9_io_DataValid = Statvalid & check & Statvalid; // @[FlexDPU.scala 112:29 115:25 81:25]
  assign PathFinder_10_clock = clock;
  assign PathFinder_10_reset = reset;
  assign PathFinder_10_io_Stationary_matrix_0_0 = Statvalid & check ? io_Stationary_matrix_0_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_0_1 = Statvalid & check ? io_Stationary_matrix_0_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_0_2 = Statvalid & check ? io_Stationary_matrix_0_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_0_3 = Statvalid & check ? io_Stationary_matrix_0_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_0_4 = Statvalid & check ? io_Stationary_matrix_0_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_0_5 = Statvalid & check ? io_Stationary_matrix_0_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_0_6 = Statvalid & check ? io_Stationary_matrix_0_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_0_7 = Statvalid & check ? io_Stationary_matrix_0_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_1_0 = Statvalid & check ? io_Stationary_matrix_1_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_1_1 = Statvalid & check ? io_Stationary_matrix_1_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_1_2 = Statvalid & check ? io_Stationary_matrix_1_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_1_3 = Statvalid & check ? io_Stationary_matrix_1_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_1_4 = Statvalid & check ? io_Stationary_matrix_1_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_1_5 = Statvalid & check ? io_Stationary_matrix_1_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_1_6 = Statvalid & check ? io_Stationary_matrix_1_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_1_7 = Statvalid & check ? io_Stationary_matrix_1_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_2_0 = Statvalid & check ? io_Stationary_matrix_2_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_2_1 = Statvalid & check ? io_Stationary_matrix_2_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_2_2 = Statvalid & check ? io_Stationary_matrix_2_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_2_3 = Statvalid & check ? io_Stationary_matrix_2_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_2_4 = Statvalid & check ? io_Stationary_matrix_2_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_2_5 = Statvalid & check ? io_Stationary_matrix_2_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_2_6 = Statvalid & check ? io_Stationary_matrix_2_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_2_7 = Statvalid & check ? io_Stationary_matrix_2_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_3_0 = Statvalid & check ? io_Stationary_matrix_3_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_3_1 = Statvalid & check ? io_Stationary_matrix_3_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_3_2 = Statvalid & check ? io_Stationary_matrix_3_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_3_3 = Statvalid & check ? io_Stationary_matrix_3_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_3_4 = Statvalid & check ? io_Stationary_matrix_3_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_3_5 = Statvalid & check ? io_Stationary_matrix_3_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_3_6 = Statvalid & check ? io_Stationary_matrix_3_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_3_7 = Statvalid & check ? io_Stationary_matrix_3_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_4_0 = Statvalid & check ? io_Stationary_matrix_4_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_4_1 = Statvalid & check ? io_Stationary_matrix_4_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_4_2 = Statvalid & check ? io_Stationary_matrix_4_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_4_3 = Statvalid & check ? io_Stationary_matrix_4_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_4_4 = Statvalid & check ? io_Stationary_matrix_4_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_4_5 = Statvalid & check ? io_Stationary_matrix_4_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_4_6 = Statvalid & check ? io_Stationary_matrix_4_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_4_7 = Statvalid & check ? io_Stationary_matrix_4_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_5_0 = Statvalid & check ? io_Stationary_matrix_5_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_5_1 = Statvalid & check ? io_Stationary_matrix_5_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_5_2 = Statvalid & check ? io_Stationary_matrix_5_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_5_3 = Statvalid & check ? io_Stationary_matrix_5_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_5_4 = Statvalid & check ? io_Stationary_matrix_5_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_5_5 = Statvalid & check ? io_Stationary_matrix_5_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_5_6 = Statvalid & check ? io_Stationary_matrix_5_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_5_7 = Statvalid & check ? io_Stationary_matrix_5_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_6_0 = Statvalid & check ? io_Stationary_matrix_6_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_6_1 = Statvalid & check ? io_Stationary_matrix_6_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_6_2 = Statvalid & check ? io_Stationary_matrix_6_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_6_3 = Statvalid & check ? io_Stationary_matrix_6_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_6_4 = Statvalid & check ? io_Stationary_matrix_6_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_6_5 = Statvalid & check ? io_Stationary_matrix_6_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_6_6 = Statvalid & check ? io_Stationary_matrix_6_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_6_7 = Statvalid & check ? io_Stationary_matrix_6_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_7_0 = Statvalid & check ? io_Stationary_matrix_7_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_7_1 = Statvalid & check ? io_Stationary_matrix_7_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_7_2 = Statvalid & check ? io_Stationary_matrix_7_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_7_3 = Statvalid & check ? io_Stationary_matrix_7_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_7_4 = Statvalid & check ? io_Stationary_matrix_7_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_7_5 = Statvalid & check ? io_Stationary_matrix_7_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_7_6 = Statvalid & check ? io_Stationary_matrix_7_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Stationary_matrix_7_7 = Statvalid & check ? io_Stationary_matrix_7_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_10_io_Streaming_matrix_0 = _GEN_397[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_10_io_Streaming_matrix_1 = _GEN_398[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_10_io_Streaming_matrix_2 = _GEN_399[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_10_io_Streaming_matrix_3 = _GEN_400[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_10_io_Streaming_matrix_4 = _GEN_401[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_10_io_Streaming_matrix_5 = _GEN_402[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_10_io_Streaming_matrix_6 = _GEN_403[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_10_io_Streaming_matrix_7 = _GEN_404[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_10_io_NoDPE = {{28'd0}, _GEN_1138}; // @[FlexDPU.scala 77:21]
  assign PathFinder_10_io_DataValid = Statvalid & check & Statvalid; // @[FlexDPU.scala 112:29 115:25 81:25]
  assign PathFinder_11_clock = clock;
  assign PathFinder_11_reset = reset;
  assign PathFinder_11_io_Stationary_matrix_0_0 = Statvalid & check ? io_Stationary_matrix_0_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_0_1 = Statvalid & check ? io_Stationary_matrix_0_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_0_2 = Statvalid & check ? io_Stationary_matrix_0_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_0_3 = Statvalid & check ? io_Stationary_matrix_0_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_0_4 = Statvalid & check ? io_Stationary_matrix_0_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_0_5 = Statvalid & check ? io_Stationary_matrix_0_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_0_6 = Statvalid & check ? io_Stationary_matrix_0_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_0_7 = Statvalid & check ? io_Stationary_matrix_0_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_1_0 = Statvalid & check ? io_Stationary_matrix_1_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_1_1 = Statvalid & check ? io_Stationary_matrix_1_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_1_2 = Statvalid & check ? io_Stationary_matrix_1_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_1_3 = Statvalid & check ? io_Stationary_matrix_1_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_1_4 = Statvalid & check ? io_Stationary_matrix_1_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_1_5 = Statvalid & check ? io_Stationary_matrix_1_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_1_6 = Statvalid & check ? io_Stationary_matrix_1_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_1_7 = Statvalid & check ? io_Stationary_matrix_1_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_2_0 = Statvalid & check ? io_Stationary_matrix_2_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_2_1 = Statvalid & check ? io_Stationary_matrix_2_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_2_2 = Statvalid & check ? io_Stationary_matrix_2_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_2_3 = Statvalid & check ? io_Stationary_matrix_2_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_2_4 = Statvalid & check ? io_Stationary_matrix_2_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_2_5 = Statvalid & check ? io_Stationary_matrix_2_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_2_6 = Statvalid & check ? io_Stationary_matrix_2_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_2_7 = Statvalid & check ? io_Stationary_matrix_2_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_3_0 = Statvalid & check ? io_Stationary_matrix_3_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_3_1 = Statvalid & check ? io_Stationary_matrix_3_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_3_2 = Statvalid & check ? io_Stationary_matrix_3_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_3_3 = Statvalid & check ? io_Stationary_matrix_3_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_3_4 = Statvalid & check ? io_Stationary_matrix_3_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_3_5 = Statvalid & check ? io_Stationary_matrix_3_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_3_6 = Statvalid & check ? io_Stationary_matrix_3_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_3_7 = Statvalid & check ? io_Stationary_matrix_3_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_4_0 = Statvalid & check ? io_Stationary_matrix_4_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_4_1 = Statvalid & check ? io_Stationary_matrix_4_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_4_2 = Statvalid & check ? io_Stationary_matrix_4_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_4_3 = Statvalid & check ? io_Stationary_matrix_4_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_4_4 = Statvalid & check ? io_Stationary_matrix_4_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_4_5 = Statvalid & check ? io_Stationary_matrix_4_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_4_6 = Statvalid & check ? io_Stationary_matrix_4_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_4_7 = Statvalid & check ? io_Stationary_matrix_4_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_5_0 = Statvalid & check ? io_Stationary_matrix_5_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_5_1 = Statvalid & check ? io_Stationary_matrix_5_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_5_2 = Statvalid & check ? io_Stationary_matrix_5_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_5_3 = Statvalid & check ? io_Stationary_matrix_5_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_5_4 = Statvalid & check ? io_Stationary_matrix_5_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_5_5 = Statvalid & check ? io_Stationary_matrix_5_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_5_6 = Statvalid & check ? io_Stationary_matrix_5_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_5_7 = Statvalid & check ? io_Stationary_matrix_5_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_6_0 = Statvalid & check ? io_Stationary_matrix_6_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_6_1 = Statvalid & check ? io_Stationary_matrix_6_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_6_2 = Statvalid & check ? io_Stationary_matrix_6_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_6_3 = Statvalid & check ? io_Stationary_matrix_6_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_6_4 = Statvalid & check ? io_Stationary_matrix_6_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_6_5 = Statvalid & check ? io_Stationary_matrix_6_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_6_6 = Statvalid & check ? io_Stationary_matrix_6_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_6_7 = Statvalid & check ? io_Stationary_matrix_6_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_7_0 = Statvalid & check ? io_Stationary_matrix_7_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_7_1 = Statvalid & check ? io_Stationary_matrix_7_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_7_2 = Statvalid & check ? io_Stationary_matrix_7_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_7_3 = Statvalid & check ? io_Stationary_matrix_7_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_7_4 = Statvalid & check ? io_Stationary_matrix_7_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_7_5 = Statvalid & check ? io_Stationary_matrix_7_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_7_6 = Statvalid & check ? io_Stationary_matrix_7_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Stationary_matrix_7_7 = Statvalid & check ? io_Stationary_matrix_7_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_11_io_Streaming_matrix_0 = _GEN_397[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_11_io_Streaming_matrix_1 = _GEN_398[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_11_io_Streaming_matrix_2 = _GEN_399[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_11_io_Streaming_matrix_3 = _GEN_400[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_11_io_Streaming_matrix_4 = _GEN_401[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_11_io_Streaming_matrix_5 = _GEN_402[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_11_io_Streaming_matrix_6 = _GEN_403[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_11_io_Streaming_matrix_7 = _GEN_404[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_11_io_NoDPE = {{28'd0}, _GEN_1211}; // @[FlexDPU.scala 77:21]
  assign PathFinder_11_io_DataValid = Statvalid & check & Statvalid; // @[FlexDPU.scala 112:29 115:25 81:25]
  assign PathFinder_12_clock = clock;
  assign PathFinder_12_reset = reset;
  assign PathFinder_12_io_Stationary_matrix_0_0 = Statvalid & check ? io_Stationary_matrix_0_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_0_1 = Statvalid & check ? io_Stationary_matrix_0_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_0_2 = Statvalid & check ? io_Stationary_matrix_0_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_0_3 = Statvalid & check ? io_Stationary_matrix_0_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_0_4 = Statvalid & check ? io_Stationary_matrix_0_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_0_5 = Statvalid & check ? io_Stationary_matrix_0_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_0_6 = Statvalid & check ? io_Stationary_matrix_0_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_0_7 = Statvalid & check ? io_Stationary_matrix_0_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_1_0 = Statvalid & check ? io_Stationary_matrix_1_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_1_1 = Statvalid & check ? io_Stationary_matrix_1_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_1_2 = Statvalid & check ? io_Stationary_matrix_1_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_1_3 = Statvalid & check ? io_Stationary_matrix_1_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_1_4 = Statvalid & check ? io_Stationary_matrix_1_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_1_5 = Statvalid & check ? io_Stationary_matrix_1_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_1_6 = Statvalid & check ? io_Stationary_matrix_1_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_1_7 = Statvalid & check ? io_Stationary_matrix_1_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_2_0 = Statvalid & check ? io_Stationary_matrix_2_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_2_1 = Statvalid & check ? io_Stationary_matrix_2_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_2_2 = Statvalid & check ? io_Stationary_matrix_2_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_2_3 = Statvalid & check ? io_Stationary_matrix_2_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_2_4 = Statvalid & check ? io_Stationary_matrix_2_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_2_5 = Statvalid & check ? io_Stationary_matrix_2_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_2_6 = Statvalid & check ? io_Stationary_matrix_2_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_2_7 = Statvalid & check ? io_Stationary_matrix_2_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_3_0 = Statvalid & check ? io_Stationary_matrix_3_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_3_1 = Statvalid & check ? io_Stationary_matrix_3_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_3_2 = Statvalid & check ? io_Stationary_matrix_3_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_3_3 = Statvalid & check ? io_Stationary_matrix_3_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_3_4 = Statvalid & check ? io_Stationary_matrix_3_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_3_5 = Statvalid & check ? io_Stationary_matrix_3_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_3_6 = Statvalid & check ? io_Stationary_matrix_3_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_3_7 = Statvalid & check ? io_Stationary_matrix_3_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_4_0 = Statvalid & check ? io_Stationary_matrix_4_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_4_1 = Statvalid & check ? io_Stationary_matrix_4_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_4_2 = Statvalid & check ? io_Stationary_matrix_4_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_4_3 = Statvalid & check ? io_Stationary_matrix_4_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_4_4 = Statvalid & check ? io_Stationary_matrix_4_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_4_5 = Statvalid & check ? io_Stationary_matrix_4_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_4_6 = Statvalid & check ? io_Stationary_matrix_4_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_4_7 = Statvalid & check ? io_Stationary_matrix_4_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_5_0 = Statvalid & check ? io_Stationary_matrix_5_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_5_1 = Statvalid & check ? io_Stationary_matrix_5_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_5_2 = Statvalid & check ? io_Stationary_matrix_5_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_5_3 = Statvalid & check ? io_Stationary_matrix_5_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_5_4 = Statvalid & check ? io_Stationary_matrix_5_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_5_5 = Statvalid & check ? io_Stationary_matrix_5_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_5_6 = Statvalid & check ? io_Stationary_matrix_5_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_5_7 = Statvalid & check ? io_Stationary_matrix_5_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_6_0 = Statvalid & check ? io_Stationary_matrix_6_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_6_1 = Statvalid & check ? io_Stationary_matrix_6_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_6_2 = Statvalid & check ? io_Stationary_matrix_6_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_6_3 = Statvalid & check ? io_Stationary_matrix_6_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_6_4 = Statvalid & check ? io_Stationary_matrix_6_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_6_5 = Statvalid & check ? io_Stationary_matrix_6_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_6_6 = Statvalid & check ? io_Stationary_matrix_6_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_6_7 = Statvalid & check ? io_Stationary_matrix_6_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_7_0 = Statvalid & check ? io_Stationary_matrix_7_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_7_1 = Statvalid & check ? io_Stationary_matrix_7_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_7_2 = Statvalid & check ? io_Stationary_matrix_7_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_7_3 = Statvalid & check ? io_Stationary_matrix_7_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_7_4 = Statvalid & check ? io_Stationary_matrix_7_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_7_5 = Statvalid & check ? io_Stationary_matrix_7_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_7_6 = Statvalid & check ? io_Stationary_matrix_7_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Stationary_matrix_7_7 = Statvalid & check ? io_Stationary_matrix_7_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_12_io_Streaming_matrix_0 = _GEN_397[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_12_io_Streaming_matrix_1 = _GEN_398[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_12_io_Streaming_matrix_2 = _GEN_399[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_12_io_Streaming_matrix_3 = _GEN_400[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_12_io_Streaming_matrix_4 = _GEN_401[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_12_io_Streaming_matrix_5 = _GEN_402[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_12_io_Streaming_matrix_6 = _GEN_403[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_12_io_Streaming_matrix_7 = _GEN_404[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_12_io_NoDPE = {{28'd0}, _GEN_1284}; // @[FlexDPU.scala 77:21]
  assign PathFinder_12_io_DataValid = Statvalid & check & Statvalid; // @[FlexDPU.scala 112:29 115:25 81:25]
  assign PathFinder_13_clock = clock;
  assign PathFinder_13_reset = reset;
  assign PathFinder_13_io_Stationary_matrix_0_0 = Statvalid & check ? io_Stationary_matrix_0_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_0_1 = Statvalid & check ? io_Stationary_matrix_0_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_0_2 = Statvalid & check ? io_Stationary_matrix_0_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_0_3 = Statvalid & check ? io_Stationary_matrix_0_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_0_4 = Statvalid & check ? io_Stationary_matrix_0_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_0_5 = Statvalid & check ? io_Stationary_matrix_0_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_0_6 = Statvalid & check ? io_Stationary_matrix_0_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_0_7 = Statvalid & check ? io_Stationary_matrix_0_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_1_0 = Statvalid & check ? io_Stationary_matrix_1_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_1_1 = Statvalid & check ? io_Stationary_matrix_1_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_1_2 = Statvalid & check ? io_Stationary_matrix_1_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_1_3 = Statvalid & check ? io_Stationary_matrix_1_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_1_4 = Statvalid & check ? io_Stationary_matrix_1_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_1_5 = Statvalid & check ? io_Stationary_matrix_1_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_1_6 = Statvalid & check ? io_Stationary_matrix_1_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_1_7 = Statvalid & check ? io_Stationary_matrix_1_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_2_0 = Statvalid & check ? io_Stationary_matrix_2_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_2_1 = Statvalid & check ? io_Stationary_matrix_2_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_2_2 = Statvalid & check ? io_Stationary_matrix_2_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_2_3 = Statvalid & check ? io_Stationary_matrix_2_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_2_4 = Statvalid & check ? io_Stationary_matrix_2_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_2_5 = Statvalid & check ? io_Stationary_matrix_2_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_2_6 = Statvalid & check ? io_Stationary_matrix_2_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_2_7 = Statvalid & check ? io_Stationary_matrix_2_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_3_0 = Statvalid & check ? io_Stationary_matrix_3_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_3_1 = Statvalid & check ? io_Stationary_matrix_3_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_3_2 = Statvalid & check ? io_Stationary_matrix_3_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_3_3 = Statvalid & check ? io_Stationary_matrix_3_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_3_4 = Statvalid & check ? io_Stationary_matrix_3_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_3_5 = Statvalid & check ? io_Stationary_matrix_3_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_3_6 = Statvalid & check ? io_Stationary_matrix_3_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_3_7 = Statvalid & check ? io_Stationary_matrix_3_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_4_0 = Statvalid & check ? io_Stationary_matrix_4_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_4_1 = Statvalid & check ? io_Stationary_matrix_4_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_4_2 = Statvalid & check ? io_Stationary_matrix_4_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_4_3 = Statvalid & check ? io_Stationary_matrix_4_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_4_4 = Statvalid & check ? io_Stationary_matrix_4_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_4_5 = Statvalid & check ? io_Stationary_matrix_4_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_4_6 = Statvalid & check ? io_Stationary_matrix_4_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_4_7 = Statvalid & check ? io_Stationary_matrix_4_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_5_0 = Statvalid & check ? io_Stationary_matrix_5_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_5_1 = Statvalid & check ? io_Stationary_matrix_5_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_5_2 = Statvalid & check ? io_Stationary_matrix_5_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_5_3 = Statvalid & check ? io_Stationary_matrix_5_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_5_4 = Statvalid & check ? io_Stationary_matrix_5_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_5_5 = Statvalid & check ? io_Stationary_matrix_5_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_5_6 = Statvalid & check ? io_Stationary_matrix_5_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_5_7 = Statvalid & check ? io_Stationary_matrix_5_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_6_0 = Statvalid & check ? io_Stationary_matrix_6_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_6_1 = Statvalid & check ? io_Stationary_matrix_6_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_6_2 = Statvalid & check ? io_Stationary_matrix_6_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_6_3 = Statvalid & check ? io_Stationary_matrix_6_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_6_4 = Statvalid & check ? io_Stationary_matrix_6_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_6_5 = Statvalid & check ? io_Stationary_matrix_6_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_6_6 = Statvalid & check ? io_Stationary_matrix_6_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_6_7 = Statvalid & check ? io_Stationary_matrix_6_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_7_0 = Statvalid & check ? io_Stationary_matrix_7_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_7_1 = Statvalid & check ? io_Stationary_matrix_7_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_7_2 = Statvalid & check ? io_Stationary_matrix_7_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_7_3 = Statvalid & check ? io_Stationary_matrix_7_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_7_4 = Statvalid & check ? io_Stationary_matrix_7_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_7_5 = Statvalid & check ? io_Stationary_matrix_7_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_7_6 = Statvalid & check ? io_Stationary_matrix_7_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Stationary_matrix_7_7 = Statvalid & check ? io_Stationary_matrix_7_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_13_io_Streaming_matrix_0 = _GEN_397[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_13_io_Streaming_matrix_1 = _GEN_398[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_13_io_Streaming_matrix_2 = _GEN_399[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_13_io_Streaming_matrix_3 = _GEN_400[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_13_io_Streaming_matrix_4 = _GEN_401[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_13_io_Streaming_matrix_5 = _GEN_402[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_13_io_Streaming_matrix_6 = _GEN_403[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_13_io_Streaming_matrix_7 = _GEN_404[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_13_io_NoDPE = {{28'd0}, _GEN_1357}; // @[FlexDPU.scala 77:21]
  assign PathFinder_13_io_DataValid = Statvalid & check & Statvalid; // @[FlexDPU.scala 112:29 115:25 81:25]
  assign PathFinder_14_clock = clock;
  assign PathFinder_14_reset = reset;
  assign PathFinder_14_io_Stationary_matrix_0_0 = Statvalid & check ? io_Stationary_matrix_0_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_0_1 = Statvalid & check ? io_Stationary_matrix_0_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_0_2 = Statvalid & check ? io_Stationary_matrix_0_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_0_3 = Statvalid & check ? io_Stationary_matrix_0_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_0_4 = Statvalid & check ? io_Stationary_matrix_0_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_0_5 = Statvalid & check ? io_Stationary_matrix_0_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_0_6 = Statvalid & check ? io_Stationary_matrix_0_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_0_7 = Statvalid & check ? io_Stationary_matrix_0_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_1_0 = Statvalid & check ? io_Stationary_matrix_1_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_1_1 = Statvalid & check ? io_Stationary_matrix_1_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_1_2 = Statvalid & check ? io_Stationary_matrix_1_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_1_3 = Statvalid & check ? io_Stationary_matrix_1_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_1_4 = Statvalid & check ? io_Stationary_matrix_1_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_1_5 = Statvalid & check ? io_Stationary_matrix_1_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_1_6 = Statvalid & check ? io_Stationary_matrix_1_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_1_7 = Statvalid & check ? io_Stationary_matrix_1_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_2_0 = Statvalid & check ? io_Stationary_matrix_2_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_2_1 = Statvalid & check ? io_Stationary_matrix_2_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_2_2 = Statvalid & check ? io_Stationary_matrix_2_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_2_3 = Statvalid & check ? io_Stationary_matrix_2_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_2_4 = Statvalid & check ? io_Stationary_matrix_2_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_2_5 = Statvalid & check ? io_Stationary_matrix_2_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_2_6 = Statvalid & check ? io_Stationary_matrix_2_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_2_7 = Statvalid & check ? io_Stationary_matrix_2_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_3_0 = Statvalid & check ? io_Stationary_matrix_3_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_3_1 = Statvalid & check ? io_Stationary_matrix_3_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_3_2 = Statvalid & check ? io_Stationary_matrix_3_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_3_3 = Statvalid & check ? io_Stationary_matrix_3_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_3_4 = Statvalid & check ? io_Stationary_matrix_3_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_3_5 = Statvalid & check ? io_Stationary_matrix_3_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_3_6 = Statvalid & check ? io_Stationary_matrix_3_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_3_7 = Statvalid & check ? io_Stationary_matrix_3_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_4_0 = Statvalid & check ? io_Stationary_matrix_4_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_4_1 = Statvalid & check ? io_Stationary_matrix_4_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_4_2 = Statvalid & check ? io_Stationary_matrix_4_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_4_3 = Statvalid & check ? io_Stationary_matrix_4_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_4_4 = Statvalid & check ? io_Stationary_matrix_4_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_4_5 = Statvalid & check ? io_Stationary_matrix_4_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_4_6 = Statvalid & check ? io_Stationary_matrix_4_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_4_7 = Statvalid & check ? io_Stationary_matrix_4_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_5_0 = Statvalid & check ? io_Stationary_matrix_5_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_5_1 = Statvalid & check ? io_Stationary_matrix_5_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_5_2 = Statvalid & check ? io_Stationary_matrix_5_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_5_3 = Statvalid & check ? io_Stationary_matrix_5_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_5_4 = Statvalid & check ? io_Stationary_matrix_5_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_5_5 = Statvalid & check ? io_Stationary_matrix_5_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_5_6 = Statvalid & check ? io_Stationary_matrix_5_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_5_7 = Statvalid & check ? io_Stationary_matrix_5_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_6_0 = Statvalid & check ? io_Stationary_matrix_6_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_6_1 = Statvalid & check ? io_Stationary_matrix_6_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_6_2 = Statvalid & check ? io_Stationary_matrix_6_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_6_3 = Statvalid & check ? io_Stationary_matrix_6_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_6_4 = Statvalid & check ? io_Stationary_matrix_6_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_6_5 = Statvalid & check ? io_Stationary_matrix_6_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_6_6 = Statvalid & check ? io_Stationary_matrix_6_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_6_7 = Statvalid & check ? io_Stationary_matrix_6_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_7_0 = Statvalid & check ? io_Stationary_matrix_7_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_7_1 = Statvalid & check ? io_Stationary_matrix_7_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_7_2 = Statvalid & check ? io_Stationary_matrix_7_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_7_3 = Statvalid & check ? io_Stationary_matrix_7_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_7_4 = Statvalid & check ? io_Stationary_matrix_7_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_7_5 = Statvalid & check ? io_Stationary_matrix_7_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_7_6 = Statvalid & check ? io_Stationary_matrix_7_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Stationary_matrix_7_7 = Statvalid & check ? io_Stationary_matrix_7_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_14_io_Streaming_matrix_0 = _GEN_397[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_14_io_Streaming_matrix_1 = _GEN_398[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_14_io_Streaming_matrix_2 = _GEN_399[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_14_io_Streaming_matrix_3 = _GEN_400[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_14_io_Streaming_matrix_4 = _GEN_401[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_14_io_Streaming_matrix_5 = _GEN_402[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_14_io_Streaming_matrix_6 = _GEN_403[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_14_io_Streaming_matrix_7 = _GEN_404[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_14_io_NoDPE = {{28'd0}, _GEN_1430}; // @[FlexDPU.scala 77:21]
  assign PathFinder_14_io_DataValid = Statvalid & check & Statvalid; // @[FlexDPU.scala 112:29 115:25 81:25]
  assign PathFinder_15_clock = clock;
  assign PathFinder_15_reset = reset;
  assign PathFinder_15_io_Stationary_matrix_0_0 = Statvalid & check ? io_Stationary_matrix_0_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_0_1 = Statvalid & check ? io_Stationary_matrix_0_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_0_2 = Statvalid & check ? io_Stationary_matrix_0_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_0_3 = Statvalid & check ? io_Stationary_matrix_0_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_0_4 = Statvalid & check ? io_Stationary_matrix_0_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_0_5 = Statvalid & check ? io_Stationary_matrix_0_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_0_6 = Statvalid & check ? io_Stationary_matrix_0_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_0_7 = Statvalid & check ? io_Stationary_matrix_0_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_1_0 = Statvalid & check ? io_Stationary_matrix_1_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_1_1 = Statvalid & check ? io_Stationary_matrix_1_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_1_2 = Statvalid & check ? io_Stationary_matrix_1_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_1_3 = Statvalid & check ? io_Stationary_matrix_1_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_1_4 = Statvalid & check ? io_Stationary_matrix_1_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_1_5 = Statvalid & check ? io_Stationary_matrix_1_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_1_6 = Statvalid & check ? io_Stationary_matrix_1_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_1_7 = Statvalid & check ? io_Stationary_matrix_1_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_2_0 = Statvalid & check ? io_Stationary_matrix_2_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_2_1 = Statvalid & check ? io_Stationary_matrix_2_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_2_2 = Statvalid & check ? io_Stationary_matrix_2_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_2_3 = Statvalid & check ? io_Stationary_matrix_2_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_2_4 = Statvalid & check ? io_Stationary_matrix_2_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_2_5 = Statvalid & check ? io_Stationary_matrix_2_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_2_6 = Statvalid & check ? io_Stationary_matrix_2_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_2_7 = Statvalid & check ? io_Stationary_matrix_2_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_3_0 = Statvalid & check ? io_Stationary_matrix_3_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_3_1 = Statvalid & check ? io_Stationary_matrix_3_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_3_2 = Statvalid & check ? io_Stationary_matrix_3_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_3_3 = Statvalid & check ? io_Stationary_matrix_3_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_3_4 = Statvalid & check ? io_Stationary_matrix_3_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_3_5 = Statvalid & check ? io_Stationary_matrix_3_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_3_6 = Statvalid & check ? io_Stationary_matrix_3_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_3_7 = Statvalid & check ? io_Stationary_matrix_3_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_4_0 = Statvalid & check ? io_Stationary_matrix_4_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_4_1 = Statvalid & check ? io_Stationary_matrix_4_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_4_2 = Statvalid & check ? io_Stationary_matrix_4_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_4_3 = Statvalid & check ? io_Stationary_matrix_4_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_4_4 = Statvalid & check ? io_Stationary_matrix_4_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_4_5 = Statvalid & check ? io_Stationary_matrix_4_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_4_6 = Statvalid & check ? io_Stationary_matrix_4_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_4_7 = Statvalid & check ? io_Stationary_matrix_4_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_5_0 = Statvalid & check ? io_Stationary_matrix_5_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_5_1 = Statvalid & check ? io_Stationary_matrix_5_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_5_2 = Statvalid & check ? io_Stationary_matrix_5_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_5_3 = Statvalid & check ? io_Stationary_matrix_5_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_5_4 = Statvalid & check ? io_Stationary_matrix_5_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_5_5 = Statvalid & check ? io_Stationary_matrix_5_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_5_6 = Statvalid & check ? io_Stationary_matrix_5_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_5_7 = Statvalid & check ? io_Stationary_matrix_5_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_6_0 = Statvalid & check ? io_Stationary_matrix_6_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_6_1 = Statvalid & check ? io_Stationary_matrix_6_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_6_2 = Statvalid & check ? io_Stationary_matrix_6_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_6_3 = Statvalid & check ? io_Stationary_matrix_6_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_6_4 = Statvalid & check ? io_Stationary_matrix_6_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_6_5 = Statvalid & check ? io_Stationary_matrix_6_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_6_6 = Statvalid & check ? io_Stationary_matrix_6_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_6_7 = Statvalid & check ? io_Stationary_matrix_6_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_7_0 = Statvalid & check ? io_Stationary_matrix_7_0 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_7_1 = Statvalid & check ? io_Stationary_matrix_7_1 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_7_2 = Statvalid & check ? io_Stationary_matrix_7_2 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_7_3 = Statvalid & check ? io_Stationary_matrix_7_3 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_7_4 = Statvalid & check ? io_Stationary_matrix_7_4 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_7_5 = Statvalid & check ? io_Stationary_matrix_7_5 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_7_6 = Statvalid & check ? io_Stationary_matrix_7_6 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Stationary_matrix_7_7 = Statvalid & check ? io_Stationary_matrix_7_7 : 16'h0; // @[FlexDPU.scala 112:29 116:33 82:33]
  assign PathFinder_15_io_Streaming_matrix_0 = _GEN_397[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_15_io_Streaming_matrix_1 = _GEN_398[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_15_io_Streaming_matrix_2 = _GEN_399[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_15_io_Streaming_matrix_3 = _GEN_400[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_15_io_Streaming_matrix_4 = _GEN_401[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_15_io_Streaming_matrix_5 = _GEN_402[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_15_io_Streaming_matrix_6 = _GEN_403[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_15_io_Streaming_matrix_7 = _GEN_404[15:0]; // @[FlexDPU.scala 77:21]
  assign PathFinder_15_io_NoDPE = {{28'd0}, _GEN_1503}; // @[FlexDPU.scala 77:21]
  assign PathFinder_15_io_DataValid = Statvalid & check & Statvalid; // @[FlexDPU.scala 112:29 115:25 81:25]
  assign ivntop_clock = clock;
  assign ivntop_reset = reset;
  assign ivntop_io_Stationary_matrix_0_0 = io_Stationary_matrix_0_0; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_0_1 = io_Stationary_matrix_0_1; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_0_2 = io_Stationary_matrix_0_2; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_0_3 = io_Stationary_matrix_0_3; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_0_4 = io_Stationary_matrix_0_4; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_0_5 = io_Stationary_matrix_0_5; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_0_6 = io_Stationary_matrix_0_6; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_0_7 = io_Stationary_matrix_0_7; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_1_0 = io_Stationary_matrix_1_0; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_1_1 = io_Stationary_matrix_1_1; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_1_2 = io_Stationary_matrix_1_2; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_1_3 = io_Stationary_matrix_1_3; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_1_4 = io_Stationary_matrix_1_4; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_1_5 = io_Stationary_matrix_1_5; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_1_6 = io_Stationary_matrix_1_6; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_1_7 = io_Stationary_matrix_1_7; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_2_0 = io_Stationary_matrix_2_0; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_2_1 = io_Stationary_matrix_2_1; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_2_2 = io_Stationary_matrix_2_2; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_2_3 = io_Stationary_matrix_2_3; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_2_4 = io_Stationary_matrix_2_4; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_2_5 = io_Stationary_matrix_2_5; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_2_6 = io_Stationary_matrix_2_6; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_2_7 = io_Stationary_matrix_2_7; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_3_0 = io_Stationary_matrix_3_0; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_3_1 = io_Stationary_matrix_3_1; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_3_2 = io_Stationary_matrix_3_2; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_3_3 = io_Stationary_matrix_3_3; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_3_4 = io_Stationary_matrix_3_4; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_3_5 = io_Stationary_matrix_3_5; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_3_6 = io_Stationary_matrix_3_6; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_3_7 = io_Stationary_matrix_3_7; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_4_0 = io_Stationary_matrix_4_0; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_4_1 = io_Stationary_matrix_4_1; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_4_2 = io_Stationary_matrix_4_2; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_4_3 = io_Stationary_matrix_4_3; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_4_4 = io_Stationary_matrix_4_4; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_4_5 = io_Stationary_matrix_4_5; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_4_6 = io_Stationary_matrix_4_6; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_4_7 = io_Stationary_matrix_4_7; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_5_0 = io_Stationary_matrix_5_0; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_5_1 = io_Stationary_matrix_5_1; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_5_2 = io_Stationary_matrix_5_2; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_5_3 = io_Stationary_matrix_5_3; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_5_4 = io_Stationary_matrix_5_4; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_5_5 = io_Stationary_matrix_5_5; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_5_6 = io_Stationary_matrix_5_6; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_5_7 = io_Stationary_matrix_5_7; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_6_0 = io_Stationary_matrix_6_0; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_6_1 = io_Stationary_matrix_6_1; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_6_2 = io_Stationary_matrix_6_2; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_6_3 = io_Stationary_matrix_6_3; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_6_4 = io_Stationary_matrix_6_4; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_6_5 = io_Stationary_matrix_6_5; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_6_6 = io_Stationary_matrix_6_6; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_6_7 = io_Stationary_matrix_6_7; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_7_0 = io_Stationary_matrix_7_0; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_7_1 = io_Stationary_matrix_7_1; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_7_2 = io_Stationary_matrix_7_2; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_7_3 = io_Stationary_matrix_7_3; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_7_4 = io_Stationary_matrix_7_4; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_7_5 = io_Stationary_matrix_7_5; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_7_6 = io_Stationary_matrix_7_6; // @[FlexDPU.scala 88:27]
  assign ivntop_io_Stationary_matrix_7_7 = io_Stationary_matrix_7_7; // @[FlexDPU.scala 88:27]
  assign MuxesWrapper_io_valid = PathFinder_io_PF_Valid; // @[FlexDPU.scala 77:{21,21}]
  assign MuxesWrapper_io_src_0 = {{16'd0}, PF_0_Source_0}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_io_src_1 = {{16'd0}, PF_0_Source_1}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_io_src_2 = {{16'd0}, PF_0_Source_2}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_io_src_3 = {{16'd0}, PF_0_Source_3}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_io_muxes_0 = {{28'd0}, PF_0_i_mux_bus_0}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_io_muxes_1 = {{28'd0}, PF_0_i_mux_bus_1}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_io_muxes_2 = {{28'd0}, PF_0_i_mux_bus_2}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_io_muxes_3 = {{28'd0}, PF_0_i_mux_bus_3}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_1_io_valid = PathFinder_1_io_PF_Valid; // @[FlexDPU.scala 77:{21,21}]
  assign MuxesWrapper_1_io_src_0 = {{16'd0}, PF_1_Source_0}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_1_io_src_1 = {{16'd0}, PF_1_Source_1}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_1_io_src_2 = {{16'd0}, PF_1_Source_2}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_1_io_src_3 = {{16'd0}, PF_1_Source_3}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_1_io_muxes_0 = {{28'd0}, PF_1_i_mux_bus_0}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_1_io_muxes_1 = {{28'd0}, PF_1_i_mux_bus_1}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_1_io_muxes_2 = {{28'd0}, PF_1_i_mux_bus_2}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_1_io_muxes_3 = {{28'd0}, PF_1_i_mux_bus_3}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_2_io_valid = PathFinder_2_io_PF_Valid; // @[FlexDPU.scala 77:{21,21}]
  assign MuxesWrapper_2_io_src_0 = {{16'd0}, PF_2_Source_0}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_2_io_src_1 = {{16'd0}, PF_2_Source_1}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_2_io_src_2 = {{16'd0}, PF_2_Source_2}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_2_io_src_3 = {{16'd0}, PF_2_Source_3}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_2_io_muxes_0 = {{28'd0}, PF_2_i_mux_bus_0}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_2_io_muxes_1 = {{28'd0}, PF_2_i_mux_bus_1}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_2_io_muxes_2 = {{28'd0}, PF_2_i_mux_bus_2}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_2_io_muxes_3 = {{28'd0}, PF_2_i_mux_bus_3}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_3_io_valid = PathFinder_3_io_PF_Valid; // @[FlexDPU.scala 77:{21,21}]
  assign MuxesWrapper_3_io_src_0 = {{16'd0}, PF_3_Source_0}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_3_io_src_1 = {{16'd0}, PF_3_Source_1}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_3_io_src_2 = {{16'd0}, PF_3_Source_2}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_3_io_src_3 = {{16'd0}, PF_3_Source_3}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_3_io_muxes_0 = {{28'd0}, PF_3_i_mux_bus_0}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_3_io_muxes_1 = {{28'd0}, PF_3_i_mux_bus_1}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_3_io_muxes_2 = {{28'd0}, PF_3_i_mux_bus_2}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_3_io_muxes_3 = {{28'd0}, PF_3_i_mux_bus_3}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_4_io_valid = PathFinder_4_io_PF_Valid; // @[FlexDPU.scala 77:{21,21}]
  assign MuxesWrapper_4_io_src_0 = {{16'd0}, PF_4_Source_0}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_4_io_src_1 = {{16'd0}, PF_4_Source_1}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_4_io_src_2 = {{16'd0}, PF_4_Source_2}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_4_io_src_3 = {{16'd0}, PF_4_Source_3}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_4_io_muxes_0 = {{28'd0}, PF_4_i_mux_bus_0}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_4_io_muxes_1 = {{28'd0}, PF_4_i_mux_bus_1}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_4_io_muxes_2 = {{28'd0}, PF_4_i_mux_bus_2}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_4_io_muxes_3 = {{28'd0}, PF_4_i_mux_bus_3}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_5_io_valid = PathFinder_5_io_PF_Valid; // @[FlexDPU.scala 77:{21,21}]
  assign MuxesWrapper_5_io_src_0 = {{16'd0}, PF_5_Source_0}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_5_io_src_1 = {{16'd0}, PF_5_Source_1}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_5_io_src_2 = {{16'd0}, PF_5_Source_2}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_5_io_src_3 = {{16'd0}, PF_5_Source_3}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_5_io_muxes_0 = {{28'd0}, PF_5_i_mux_bus_0}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_5_io_muxes_1 = {{28'd0}, PF_5_i_mux_bus_1}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_5_io_muxes_2 = {{28'd0}, PF_5_i_mux_bus_2}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_5_io_muxes_3 = {{28'd0}, PF_5_i_mux_bus_3}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_6_io_valid = PathFinder_6_io_PF_Valid; // @[FlexDPU.scala 77:{21,21}]
  assign MuxesWrapper_6_io_src_0 = {{16'd0}, PF_6_Source_0}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_6_io_src_1 = {{16'd0}, PF_6_Source_1}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_6_io_src_2 = {{16'd0}, PF_6_Source_2}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_6_io_src_3 = {{16'd0}, PF_6_Source_3}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_6_io_muxes_0 = {{28'd0}, PF_6_i_mux_bus_0}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_6_io_muxes_1 = {{28'd0}, PF_6_i_mux_bus_1}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_6_io_muxes_2 = {{28'd0}, PF_6_i_mux_bus_2}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_6_io_muxes_3 = {{28'd0}, PF_6_i_mux_bus_3}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_7_io_valid = PathFinder_7_io_PF_Valid; // @[FlexDPU.scala 77:{21,21}]
  assign MuxesWrapper_7_io_src_0 = {{16'd0}, PF_7_Source_0}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_7_io_src_1 = {{16'd0}, PF_7_Source_1}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_7_io_src_2 = {{16'd0}, PF_7_Source_2}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_7_io_src_3 = {{16'd0}, PF_7_Source_3}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_7_io_muxes_0 = {{28'd0}, PF_7_i_mux_bus_0}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_7_io_muxes_1 = {{28'd0}, PF_7_i_mux_bus_1}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_7_io_muxes_2 = {{28'd0}, PF_7_i_mux_bus_2}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_7_io_muxes_3 = {{28'd0}, PF_7_i_mux_bus_3}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_8_io_valid = PathFinder_8_io_PF_Valid; // @[FlexDPU.scala 77:{21,21}]
  assign MuxesWrapper_8_io_src_0 = {{16'd0}, PF_8_Source_0}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_8_io_src_1 = {{16'd0}, PF_8_Source_1}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_8_io_src_2 = {{16'd0}, PF_8_Source_2}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_8_io_src_3 = {{16'd0}, PF_8_Source_3}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_8_io_muxes_0 = {{28'd0}, PF_8_i_mux_bus_0}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_8_io_muxes_1 = {{28'd0}, PF_8_i_mux_bus_1}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_8_io_muxes_2 = {{28'd0}, PF_8_i_mux_bus_2}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_8_io_muxes_3 = {{28'd0}, PF_8_i_mux_bus_3}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_9_io_valid = PathFinder_9_io_PF_Valid; // @[FlexDPU.scala 77:{21,21}]
  assign MuxesWrapper_9_io_src_0 = {{16'd0}, PF_9_Source_0}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_9_io_src_1 = {{16'd0}, PF_9_Source_1}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_9_io_src_2 = {{16'd0}, PF_9_Source_2}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_9_io_src_3 = {{16'd0}, PF_9_Source_3}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_9_io_muxes_0 = {{28'd0}, PF_9_i_mux_bus_0}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_9_io_muxes_1 = {{28'd0}, PF_9_i_mux_bus_1}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_9_io_muxes_2 = {{28'd0}, PF_9_i_mux_bus_2}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_9_io_muxes_3 = {{28'd0}, PF_9_i_mux_bus_3}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_10_io_valid = PathFinder_10_io_PF_Valid; // @[FlexDPU.scala 77:{21,21}]
  assign MuxesWrapper_10_io_src_0 = {{16'd0}, PF_10_Source_0}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_10_io_src_1 = {{16'd0}, PF_10_Source_1}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_10_io_src_2 = {{16'd0}, PF_10_Source_2}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_10_io_src_3 = {{16'd0}, PF_10_Source_3}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_10_io_muxes_0 = {{28'd0}, PF_10_i_mux_bus_0}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_10_io_muxes_1 = {{28'd0}, PF_10_i_mux_bus_1}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_10_io_muxes_2 = {{28'd0}, PF_10_i_mux_bus_2}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_10_io_muxes_3 = {{28'd0}, PF_10_i_mux_bus_3}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_11_io_valid = PathFinder_11_io_PF_Valid; // @[FlexDPU.scala 77:{21,21}]
  assign MuxesWrapper_11_io_src_0 = {{16'd0}, PF_11_Source_0}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_11_io_src_1 = {{16'd0}, PF_11_Source_1}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_11_io_src_2 = {{16'd0}, PF_11_Source_2}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_11_io_src_3 = {{16'd0}, PF_11_Source_3}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_11_io_muxes_0 = {{28'd0}, PF_11_i_mux_bus_0}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_11_io_muxes_1 = {{28'd0}, PF_11_i_mux_bus_1}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_11_io_muxes_2 = {{28'd0}, PF_11_i_mux_bus_2}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_11_io_muxes_3 = {{28'd0}, PF_11_i_mux_bus_3}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_12_io_valid = PathFinder_12_io_PF_Valid; // @[FlexDPU.scala 77:{21,21}]
  assign MuxesWrapper_12_io_src_0 = {{16'd0}, PF_12_Source_0}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_12_io_src_1 = {{16'd0}, PF_12_Source_1}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_12_io_src_2 = {{16'd0}, PF_12_Source_2}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_12_io_src_3 = {{16'd0}, PF_12_Source_3}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_12_io_muxes_0 = {{28'd0}, PF_12_i_mux_bus_0}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_12_io_muxes_1 = {{28'd0}, PF_12_i_mux_bus_1}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_12_io_muxes_2 = {{28'd0}, PF_12_i_mux_bus_2}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_12_io_muxes_3 = {{28'd0}, PF_12_i_mux_bus_3}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_13_io_valid = PathFinder_13_io_PF_Valid; // @[FlexDPU.scala 77:{21,21}]
  assign MuxesWrapper_13_io_src_0 = {{16'd0}, PF_13_Source_0}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_13_io_src_1 = {{16'd0}, PF_13_Source_1}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_13_io_src_2 = {{16'd0}, PF_13_Source_2}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_13_io_src_3 = {{16'd0}, PF_13_Source_3}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_13_io_muxes_0 = {{28'd0}, PF_13_i_mux_bus_0}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_13_io_muxes_1 = {{28'd0}, PF_13_i_mux_bus_1}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_13_io_muxes_2 = {{28'd0}, PF_13_i_mux_bus_2}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_13_io_muxes_3 = {{28'd0}, PF_13_i_mux_bus_3}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_14_io_valid = PathFinder_14_io_PF_Valid; // @[FlexDPU.scala 77:{21,21}]
  assign MuxesWrapper_14_io_src_0 = {{16'd0}, PF_14_Source_0}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_14_io_src_1 = {{16'd0}, PF_14_Source_1}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_14_io_src_2 = {{16'd0}, PF_14_Source_2}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_14_io_src_3 = {{16'd0}, PF_14_Source_3}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_14_io_muxes_0 = {{28'd0}, PF_14_i_mux_bus_0}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_14_io_muxes_1 = {{28'd0}, PF_14_i_mux_bus_1}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_14_io_muxes_2 = {{28'd0}, PF_14_i_mux_bus_2}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_14_io_muxes_3 = {{28'd0}, PF_14_i_mux_bus_3}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_15_io_valid = PathFinder_15_io_PF_Valid; // @[FlexDPU.scala 77:{21,21}]
  assign MuxesWrapper_15_io_src_0 = {{16'd0}, PF_15_Source_0}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_15_io_src_1 = {{16'd0}, PF_15_Source_1}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_15_io_src_2 = {{16'd0}, PF_15_Source_2}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_15_io_src_3 = {{16'd0}, PF_15_Source_3}; // @[FlexDPU.scala 124:33 127:31]
  assign MuxesWrapper_15_io_muxes_0 = {{28'd0}, PF_15_i_mux_bus_0}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_15_io_muxes_1 = {{28'd0}, PF_15_i_mux_bus_1}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_15_io_muxes_2 = {{28'd0}, PF_15_i_mux_bus_2}; // @[FlexDPU.scala 124:33 128:33]
  assign MuxesWrapper_15_io_muxes_3 = {{28'd0}, PF_15_i_mux_bus_3}; // @[FlexDPU.scala 124:33 128:33]
  assign flexdpecom4_clock = clock;
  assign flexdpecom4_reset = reset;
  assign flexdpecom4_io_i_data_valid = 1'h1; // @[FlexDPU.scala 132:27 136:34]
  assign flexdpecom4_io_i_data_bus_0 = nonZeroValues_0[15:0]; // @[FlexDPU.scala 132:27 150:37]
  assign flexdpecom4_io_i_data_bus_1 = nonZeroValues_1[15:0]; // @[FlexDPU.scala 132:27 151:37]
  assign flexdpecom4_io_i_data_bus_2 = nonZeroValues_2[15:0]; // @[FlexDPU.scala 132:27 152:37]
  assign flexdpecom4_io_i_data_bus_3 = nonZeroValues_3[15:0]; // @[FlexDPU.scala 132:27 153:37]
  assign flexdpecom4_io_i_data_bus2_0 = MuxWrapper_0_Osrc_0[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_io_i_data_bus2_1 = MuxWrapper_0_Osrc_1[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_io_i_data_bus2_2 = MuxWrapper_0_Osrc_2[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_io_i_data_bus2_3 = MuxWrapper_0_Osrc_3[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_io_i_vn_0 = ivntop_io_o_vn_0_0; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_io_i_vn_1 = ivntop_io_o_vn_0_1; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_io_i_vn_2 = ivntop_io_o_vn_0_2; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_io_i_vn_3 = ivntop_io_o_vn_0_3; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_io_i_mux_bus_0_0 = _FDPE_0_i_mux_bus_0_0_rev_T_11 | _GEN_1792; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_io_i_mux_bus_0_1 = _FDPE_0_i_mux_bus_0_1_rev_T_11 | _GEN_1798; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_io_i_mux_bus_0_2 = _FDPE_0_i_mux_bus_0_2_rev_T_11 | _GEN_1804; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_io_i_mux_bus_0_3 = _FDPE_0_i_mux_bus_0_3_rev_T_11 | _GEN_1810; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_io_i_mux_bus_1_0 = _FDPE_0_i_mux_bus_1_0_rev_T_11 | _GEN_1816; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_io_i_mux_bus_1_1 = _FDPE_0_i_mux_bus_1_1_rev_T_11 | _GEN_1822; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_io_i_mux_bus_1_2 = _FDPE_0_i_mux_bus_1_2_rev_T_11 | _GEN_1828; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_io_i_mux_bus_2_0 = _FDPE_0_i_mux_bus_2_0_rev_T_11 | _GEN_1834; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_io_i_mux_bus_2_1 = _FDPE_0_i_mux_bus_2_1_rev_T_11 | _GEN_1840; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_io_i_mux_bus_3_0 = _FDPE_0_i_mux_bus_3_0_rev_T_11 | _GEN_1846; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_1_clock = clock;
  assign flexdpecom4_1_reset = reset;
  assign flexdpecom4_1_io_i_data_valid = 1'h1; // @[FlexDPU.scala 132:27 136:34]
  assign flexdpecom4_1_io_i_data_bus_0 = nonZeroValues_4[15:0]; // @[FlexDPU.scala 132:27 150:37]
  assign flexdpecom4_1_io_i_data_bus_1 = nonZeroValues_5[15:0]; // @[FlexDPU.scala 132:27 151:37]
  assign flexdpecom4_1_io_i_data_bus_2 = nonZeroValues_6[15:0]; // @[FlexDPU.scala 132:27 152:37]
  assign flexdpecom4_1_io_i_data_bus_3 = nonZeroValues_7[15:0]; // @[FlexDPU.scala 132:27 153:37]
  assign flexdpecom4_1_io_i_data_bus2_0 = MuxWrapper_1_Osrc_0[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_1_io_i_data_bus2_1 = MuxWrapper_1_Osrc_1[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_1_io_i_data_bus2_2 = MuxWrapper_1_Osrc_2[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_1_io_i_data_bus2_3 = MuxWrapper_1_Osrc_3[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_1_io_i_vn_0 = ivntop_io_o_vn_1_0; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_1_io_i_vn_1 = ivntop_io_o_vn_1_1; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_1_io_i_vn_2 = ivntop_io_o_vn_1_2; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_1_io_i_vn_3 = ivntop_io_o_vn_1_3; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_1_io_i_mux_bus_0_0 = _FDPE_1_i_mux_bus_0_0_rev_T_11 | _GEN_1852; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_1_io_i_mux_bus_0_1 = _FDPE_1_i_mux_bus_0_1_rev_T_11 | _GEN_1858; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_1_io_i_mux_bus_0_2 = _FDPE_1_i_mux_bus_0_2_rev_T_11 | _GEN_1864; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_1_io_i_mux_bus_0_3 = _FDPE_1_i_mux_bus_0_3_rev_T_11 | _GEN_1870; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_1_io_i_mux_bus_1_0 = _FDPE_1_i_mux_bus_1_0_rev_T_11 | _GEN_1876; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_1_io_i_mux_bus_1_1 = _FDPE_1_i_mux_bus_1_1_rev_T_11 | _GEN_1882; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_1_io_i_mux_bus_1_2 = _FDPE_1_i_mux_bus_1_2_rev_T_11 | _GEN_1888; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_1_io_i_mux_bus_2_0 = _FDPE_1_i_mux_bus_2_0_rev_T_11 | _GEN_1894; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_1_io_i_mux_bus_2_1 = _FDPE_1_i_mux_bus_2_1_rev_T_11 | _GEN_1900; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_1_io_i_mux_bus_3_0 = _FDPE_1_i_mux_bus_3_0_rev_T_11 | _GEN_1906; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_2_clock = clock;
  assign flexdpecom4_2_reset = reset;
  assign flexdpecom4_2_io_i_data_valid = 1'h1; // @[FlexDPU.scala 132:27 136:34]
  assign flexdpecom4_2_io_i_data_bus_0 = nonZeroValues_8[15:0]; // @[FlexDPU.scala 132:27 150:37]
  assign flexdpecom4_2_io_i_data_bus_1 = nonZeroValues_9[15:0]; // @[FlexDPU.scala 132:27 151:37]
  assign flexdpecom4_2_io_i_data_bus_2 = nonZeroValues_10[15:0]; // @[FlexDPU.scala 132:27 152:37]
  assign flexdpecom4_2_io_i_data_bus_3 = nonZeroValues_11[15:0]; // @[FlexDPU.scala 132:27 153:37]
  assign flexdpecom4_2_io_i_data_bus2_0 = MuxWrapper_2_Osrc_0[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_2_io_i_data_bus2_1 = MuxWrapper_2_Osrc_1[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_2_io_i_data_bus2_2 = MuxWrapper_2_Osrc_2[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_2_io_i_data_bus2_3 = MuxWrapper_2_Osrc_3[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_2_io_i_vn_0 = ivntop_io_o_vn_2_0; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_2_io_i_vn_1 = ivntop_io_o_vn_2_1; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_2_io_i_vn_2 = ivntop_io_o_vn_2_2; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_2_io_i_vn_3 = ivntop_io_o_vn_2_3; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_2_io_i_mux_bus_0_0 = _FDPE_2_i_mux_bus_0_0_rev_T_11 | _GEN_1912; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_2_io_i_mux_bus_0_1 = _FDPE_2_i_mux_bus_0_1_rev_T_11 | _GEN_1918; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_2_io_i_mux_bus_0_2 = _FDPE_2_i_mux_bus_0_2_rev_T_11 | _GEN_1924; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_2_io_i_mux_bus_0_3 = _FDPE_2_i_mux_bus_0_3_rev_T_11 | _GEN_1930; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_2_io_i_mux_bus_1_0 = _FDPE_2_i_mux_bus_1_0_rev_T_11 | _GEN_1936; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_2_io_i_mux_bus_1_1 = _FDPE_2_i_mux_bus_1_1_rev_T_11 | _GEN_1942; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_2_io_i_mux_bus_1_2 = _FDPE_2_i_mux_bus_1_2_rev_T_11 | _GEN_1948; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_2_io_i_mux_bus_2_0 = _FDPE_2_i_mux_bus_2_0_rev_T_11 | _GEN_1954; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_2_io_i_mux_bus_2_1 = _FDPE_2_i_mux_bus_2_1_rev_T_11 | _GEN_1960; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_2_io_i_mux_bus_3_0 = _FDPE_2_i_mux_bus_3_0_rev_T_11 | _GEN_1966; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_3_clock = clock;
  assign flexdpecom4_3_reset = reset;
  assign flexdpecom4_3_io_i_data_valid = 1'h1; // @[FlexDPU.scala 132:27 136:34]
  assign flexdpecom4_3_io_i_data_bus_0 = nonZeroValues_12[15:0]; // @[FlexDPU.scala 132:27 150:37]
  assign flexdpecom4_3_io_i_data_bus_1 = nonZeroValues_13[15:0]; // @[FlexDPU.scala 132:27 151:37]
  assign flexdpecom4_3_io_i_data_bus_2 = nonZeroValues_14[15:0]; // @[FlexDPU.scala 132:27 152:37]
  assign flexdpecom4_3_io_i_data_bus_3 = nonZeroValues_15[15:0]; // @[FlexDPU.scala 132:27 153:37]
  assign flexdpecom4_3_io_i_data_bus2_0 = MuxWrapper_3_Osrc_0[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_3_io_i_data_bus2_1 = MuxWrapper_3_Osrc_1[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_3_io_i_data_bus2_2 = MuxWrapper_3_Osrc_2[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_3_io_i_data_bus2_3 = MuxWrapper_3_Osrc_3[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_3_io_i_vn_0 = ivntop_io_o_vn_3_0; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_3_io_i_vn_1 = ivntop_io_o_vn_3_1; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_3_io_i_vn_2 = ivntop_io_o_vn_3_2; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_3_io_i_vn_3 = ivntop_io_o_vn_3_3; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_3_io_i_mux_bus_0_0 = _FDPE_3_i_mux_bus_0_0_rev_T_11 | _GEN_1972; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_3_io_i_mux_bus_0_1 = _FDPE_3_i_mux_bus_0_1_rev_T_11 | _GEN_1978; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_3_io_i_mux_bus_0_2 = _FDPE_3_i_mux_bus_0_2_rev_T_11 | _GEN_1984; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_3_io_i_mux_bus_0_3 = _FDPE_3_i_mux_bus_0_3_rev_T_11 | _GEN_1990; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_3_io_i_mux_bus_1_0 = _FDPE_3_i_mux_bus_1_0_rev_T_11 | _GEN_1996; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_3_io_i_mux_bus_1_1 = _FDPE_3_i_mux_bus_1_1_rev_T_11 | _GEN_2002; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_3_io_i_mux_bus_1_2 = _FDPE_3_i_mux_bus_1_2_rev_T_11 | _GEN_2008; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_3_io_i_mux_bus_2_0 = _FDPE_3_i_mux_bus_2_0_rev_T_11 | _GEN_2014; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_3_io_i_mux_bus_2_1 = _FDPE_3_i_mux_bus_2_1_rev_T_11 | _GEN_2020; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_3_io_i_mux_bus_3_0 = _FDPE_3_i_mux_bus_3_0_rev_T_11 | _GEN_2026; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_4_clock = clock;
  assign flexdpecom4_4_reset = reset;
  assign flexdpecom4_4_io_i_data_valid = 1'h1; // @[FlexDPU.scala 132:27 136:34]
  assign flexdpecom4_4_io_i_data_bus_0 = nonZeroValues_16[15:0]; // @[FlexDPU.scala 132:27 150:37]
  assign flexdpecom4_4_io_i_data_bus_1 = nonZeroValues_17[15:0]; // @[FlexDPU.scala 132:27 151:37]
  assign flexdpecom4_4_io_i_data_bus_2 = nonZeroValues_18[15:0]; // @[FlexDPU.scala 132:27 152:37]
  assign flexdpecom4_4_io_i_data_bus_3 = nonZeroValues_19[15:0]; // @[FlexDPU.scala 132:27 153:37]
  assign flexdpecom4_4_io_i_data_bus2_0 = MuxWrapper_4_Osrc_0[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_4_io_i_data_bus2_1 = MuxWrapper_4_Osrc_1[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_4_io_i_data_bus2_2 = MuxWrapper_4_Osrc_2[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_4_io_i_data_bus2_3 = MuxWrapper_4_Osrc_3[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_4_io_i_vn_0 = ivntop_io_o_vn_4_0; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_4_io_i_vn_1 = ivntop_io_o_vn_4_1; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_4_io_i_vn_2 = ivntop_io_o_vn_4_2; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_4_io_i_vn_3 = ivntop_io_o_vn_4_3; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_4_io_i_mux_bus_0_0 = _FDPE_4_i_mux_bus_0_0_rev_T_11 | _GEN_2032; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_4_io_i_mux_bus_0_1 = _FDPE_4_i_mux_bus_0_1_rev_T_11 | _GEN_2038; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_4_io_i_mux_bus_0_2 = _FDPE_4_i_mux_bus_0_2_rev_T_11 | _GEN_2044; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_4_io_i_mux_bus_0_3 = _FDPE_4_i_mux_bus_0_3_rev_T_11 | _GEN_2050; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_4_io_i_mux_bus_1_0 = _FDPE_4_i_mux_bus_1_0_rev_T_11 | _GEN_2056; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_4_io_i_mux_bus_1_1 = _FDPE_4_i_mux_bus_1_1_rev_T_11 | _GEN_2062; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_4_io_i_mux_bus_1_2 = _FDPE_4_i_mux_bus_1_2_rev_T_11 | _GEN_2068; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_4_io_i_mux_bus_2_0 = _FDPE_4_i_mux_bus_2_0_rev_T_11 | _GEN_2074; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_4_io_i_mux_bus_2_1 = _FDPE_4_i_mux_bus_2_1_rev_T_11 | _GEN_2080; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_4_io_i_mux_bus_3_0 = _FDPE_4_i_mux_bus_3_0_rev_T_11 | _GEN_2086; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_5_clock = clock;
  assign flexdpecom4_5_reset = reset;
  assign flexdpecom4_5_io_i_data_valid = 1'h1; // @[FlexDPU.scala 132:27 136:34]
  assign flexdpecom4_5_io_i_data_bus_0 = nonZeroValues_20[15:0]; // @[FlexDPU.scala 132:27 150:37]
  assign flexdpecom4_5_io_i_data_bus_1 = nonZeroValues_21[15:0]; // @[FlexDPU.scala 132:27 151:37]
  assign flexdpecom4_5_io_i_data_bus_2 = nonZeroValues_22[15:0]; // @[FlexDPU.scala 132:27 152:37]
  assign flexdpecom4_5_io_i_data_bus_3 = nonZeroValues_23[15:0]; // @[FlexDPU.scala 132:27 153:37]
  assign flexdpecom4_5_io_i_data_bus2_0 = MuxWrapper_5_Osrc_0[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_5_io_i_data_bus2_1 = MuxWrapper_5_Osrc_1[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_5_io_i_data_bus2_2 = MuxWrapper_5_Osrc_2[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_5_io_i_data_bus2_3 = MuxWrapper_5_Osrc_3[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_5_io_i_vn_0 = ivntop_io_o_vn_5_0; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_5_io_i_vn_1 = ivntop_io_o_vn_5_1; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_5_io_i_vn_2 = ivntop_io_o_vn_5_2; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_5_io_i_vn_3 = ivntop_io_o_vn_5_3; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_5_io_i_mux_bus_0_0 = _FDPE_5_i_mux_bus_0_0_rev_T_11 | _GEN_2092; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_5_io_i_mux_bus_0_1 = _FDPE_5_i_mux_bus_0_1_rev_T_11 | _GEN_2098; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_5_io_i_mux_bus_0_2 = _FDPE_5_i_mux_bus_0_2_rev_T_11 | _GEN_2104; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_5_io_i_mux_bus_0_3 = _FDPE_5_i_mux_bus_0_3_rev_T_11 | _GEN_2110; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_5_io_i_mux_bus_1_0 = _FDPE_5_i_mux_bus_1_0_rev_T_11 | _GEN_2116; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_5_io_i_mux_bus_1_1 = _FDPE_5_i_mux_bus_1_1_rev_T_11 | _GEN_2122; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_5_io_i_mux_bus_1_2 = _FDPE_5_i_mux_bus_1_2_rev_T_11 | _GEN_2128; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_5_io_i_mux_bus_2_0 = _FDPE_5_i_mux_bus_2_0_rev_T_11 | _GEN_2134; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_5_io_i_mux_bus_2_1 = _FDPE_5_i_mux_bus_2_1_rev_T_11 | _GEN_2140; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_5_io_i_mux_bus_3_0 = _FDPE_5_i_mux_bus_3_0_rev_T_11 | _GEN_2146; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_6_clock = clock;
  assign flexdpecom4_6_reset = reset;
  assign flexdpecom4_6_io_i_data_valid = 1'h1; // @[FlexDPU.scala 132:27 136:34]
  assign flexdpecom4_6_io_i_data_bus_0 = nonZeroValues_24[15:0]; // @[FlexDPU.scala 132:27 150:37]
  assign flexdpecom4_6_io_i_data_bus_1 = nonZeroValues_25[15:0]; // @[FlexDPU.scala 132:27 151:37]
  assign flexdpecom4_6_io_i_data_bus_2 = nonZeroValues_26[15:0]; // @[FlexDPU.scala 132:27 152:37]
  assign flexdpecom4_6_io_i_data_bus_3 = nonZeroValues_27[15:0]; // @[FlexDPU.scala 132:27 153:37]
  assign flexdpecom4_6_io_i_data_bus2_0 = MuxWrapper_6_Osrc_0[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_6_io_i_data_bus2_1 = MuxWrapper_6_Osrc_1[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_6_io_i_data_bus2_2 = MuxWrapper_6_Osrc_2[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_6_io_i_data_bus2_3 = MuxWrapper_6_Osrc_3[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_6_io_i_vn_0 = ivntop_io_o_vn_6_0; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_6_io_i_vn_1 = ivntop_io_o_vn_6_1; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_6_io_i_vn_2 = ivntop_io_o_vn_6_2; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_6_io_i_vn_3 = ivntop_io_o_vn_6_3; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_6_io_i_mux_bus_0_0 = _FDPE_6_i_mux_bus_0_0_rev_T_11 | _GEN_2152; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_6_io_i_mux_bus_0_1 = _FDPE_6_i_mux_bus_0_1_rev_T_11 | _GEN_2158; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_6_io_i_mux_bus_0_2 = _FDPE_6_i_mux_bus_0_2_rev_T_11 | _GEN_2164; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_6_io_i_mux_bus_0_3 = _FDPE_6_i_mux_bus_0_3_rev_T_11 | _GEN_2170; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_6_io_i_mux_bus_1_0 = _FDPE_6_i_mux_bus_1_0_rev_T_11 | _GEN_2176; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_6_io_i_mux_bus_1_1 = _FDPE_6_i_mux_bus_1_1_rev_T_11 | _GEN_2182; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_6_io_i_mux_bus_1_2 = _FDPE_6_i_mux_bus_1_2_rev_T_11 | _GEN_2188; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_6_io_i_mux_bus_2_0 = _FDPE_6_i_mux_bus_2_0_rev_T_11 | _GEN_2194; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_6_io_i_mux_bus_2_1 = _FDPE_6_i_mux_bus_2_1_rev_T_11 | _GEN_2200; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_6_io_i_mux_bus_3_0 = _FDPE_6_i_mux_bus_3_0_rev_T_11 | _GEN_2206; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_7_clock = clock;
  assign flexdpecom4_7_reset = reset;
  assign flexdpecom4_7_io_i_data_valid = 1'h1; // @[FlexDPU.scala 132:27 136:34]
  assign flexdpecom4_7_io_i_data_bus_0 = nonZeroValues_28[15:0]; // @[FlexDPU.scala 132:27 150:37]
  assign flexdpecom4_7_io_i_data_bus_1 = nonZeroValues_29[15:0]; // @[FlexDPU.scala 132:27 151:37]
  assign flexdpecom4_7_io_i_data_bus_2 = nonZeroValues_30[15:0]; // @[FlexDPU.scala 132:27 152:37]
  assign flexdpecom4_7_io_i_data_bus_3 = nonZeroValues_31[15:0]; // @[FlexDPU.scala 132:27 153:37]
  assign flexdpecom4_7_io_i_data_bus2_0 = MuxWrapper_7_Osrc_0[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_7_io_i_data_bus2_1 = MuxWrapper_7_Osrc_1[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_7_io_i_data_bus2_2 = MuxWrapper_7_Osrc_2[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_7_io_i_data_bus2_3 = MuxWrapper_7_Osrc_3[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_7_io_i_vn_0 = ivntop_io_o_vn_7_0; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_7_io_i_vn_1 = ivntop_io_o_vn_7_1; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_7_io_i_vn_2 = ivntop_io_o_vn_7_2; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_7_io_i_vn_3 = ivntop_io_o_vn_7_3; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_7_io_i_mux_bus_0_0 = _FDPE_7_i_mux_bus_0_0_rev_T_11 | _GEN_2212; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_7_io_i_mux_bus_0_1 = _FDPE_7_i_mux_bus_0_1_rev_T_11 | _GEN_2218; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_7_io_i_mux_bus_0_2 = _FDPE_7_i_mux_bus_0_2_rev_T_11 | _GEN_2224; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_7_io_i_mux_bus_0_3 = _FDPE_7_i_mux_bus_0_3_rev_T_11 | _GEN_2230; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_7_io_i_mux_bus_1_0 = _FDPE_7_i_mux_bus_1_0_rev_T_11 | _GEN_2236; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_7_io_i_mux_bus_1_1 = _FDPE_7_i_mux_bus_1_1_rev_T_11 | _GEN_2242; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_7_io_i_mux_bus_1_2 = _FDPE_7_i_mux_bus_1_2_rev_T_11 | _GEN_2248; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_7_io_i_mux_bus_2_0 = _FDPE_7_i_mux_bus_2_0_rev_T_11 | _GEN_2254; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_7_io_i_mux_bus_2_1 = _FDPE_7_i_mux_bus_2_1_rev_T_11 | _GEN_2260; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_7_io_i_mux_bus_3_0 = _FDPE_7_i_mux_bus_3_0_rev_T_11 | _GEN_2266; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_8_clock = clock;
  assign flexdpecom4_8_reset = reset;
  assign flexdpecom4_8_io_i_data_valid = 1'h1; // @[FlexDPU.scala 132:27 136:34]
  assign flexdpecom4_8_io_i_data_bus_0 = nonZeroValues_32[15:0]; // @[FlexDPU.scala 132:27 150:37]
  assign flexdpecom4_8_io_i_data_bus_1 = nonZeroValues_33[15:0]; // @[FlexDPU.scala 132:27 151:37]
  assign flexdpecom4_8_io_i_data_bus_2 = nonZeroValues_34[15:0]; // @[FlexDPU.scala 132:27 152:37]
  assign flexdpecom4_8_io_i_data_bus_3 = nonZeroValues_35[15:0]; // @[FlexDPU.scala 132:27 153:37]
  assign flexdpecom4_8_io_i_data_bus2_0 = MuxWrapper_8_Osrc_0[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_8_io_i_data_bus2_1 = MuxWrapper_8_Osrc_1[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_8_io_i_data_bus2_2 = MuxWrapper_8_Osrc_2[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_8_io_i_data_bus2_3 = MuxWrapper_8_Osrc_3[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_8_io_i_vn_0 = ivntop_io_o_vn_8_0; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_8_io_i_vn_1 = ivntop_io_o_vn_8_1; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_8_io_i_vn_2 = ivntop_io_o_vn_8_2; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_8_io_i_vn_3 = ivntop_io_o_vn_8_3; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_8_io_i_mux_bus_0_0 = _FDPE_8_i_mux_bus_0_0_rev_T_11 | _GEN_2272; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_8_io_i_mux_bus_0_1 = _FDPE_8_i_mux_bus_0_1_rev_T_11 | _GEN_2278; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_8_io_i_mux_bus_0_2 = _FDPE_8_i_mux_bus_0_2_rev_T_11 | _GEN_2284; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_8_io_i_mux_bus_0_3 = _FDPE_8_i_mux_bus_0_3_rev_T_11 | _GEN_2290; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_8_io_i_mux_bus_1_0 = _FDPE_8_i_mux_bus_1_0_rev_T_11 | _GEN_2296; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_8_io_i_mux_bus_1_1 = _FDPE_8_i_mux_bus_1_1_rev_T_11 | _GEN_2302; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_8_io_i_mux_bus_1_2 = _FDPE_8_i_mux_bus_1_2_rev_T_11 | _GEN_2308; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_8_io_i_mux_bus_2_0 = _FDPE_8_i_mux_bus_2_0_rev_T_11 | _GEN_2314; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_8_io_i_mux_bus_2_1 = _FDPE_8_i_mux_bus_2_1_rev_T_11 | _GEN_2320; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_8_io_i_mux_bus_3_0 = _FDPE_8_i_mux_bus_3_0_rev_T_11 | _GEN_2326; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_9_clock = clock;
  assign flexdpecom4_9_reset = reset;
  assign flexdpecom4_9_io_i_data_valid = 1'h1; // @[FlexDPU.scala 132:27 136:34]
  assign flexdpecom4_9_io_i_data_bus_0 = nonZeroValues_36[15:0]; // @[FlexDPU.scala 132:27 150:37]
  assign flexdpecom4_9_io_i_data_bus_1 = nonZeroValues_37[15:0]; // @[FlexDPU.scala 132:27 151:37]
  assign flexdpecom4_9_io_i_data_bus_2 = nonZeroValues_38[15:0]; // @[FlexDPU.scala 132:27 152:37]
  assign flexdpecom4_9_io_i_data_bus_3 = nonZeroValues_39[15:0]; // @[FlexDPU.scala 132:27 153:37]
  assign flexdpecom4_9_io_i_data_bus2_0 = MuxWrapper_9_Osrc_0[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_9_io_i_data_bus2_1 = MuxWrapper_9_Osrc_1[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_9_io_i_data_bus2_2 = MuxWrapper_9_Osrc_2[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_9_io_i_data_bus2_3 = MuxWrapper_9_Osrc_3[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_9_io_i_vn_0 = ivntop_io_o_vn_9_0; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_9_io_i_vn_1 = ivntop_io_o_vn_9_1; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_9_io_i_vn_2 = ivntop_io_o_vn_9_2; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_9_io_i_vn_3 = ivntop_io_o_vn_9_3; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_9_io_i_mux_bus_0_0 = _FDPE_9_i_mux_bus_0_0_rev_T_11 | _GEN_2332; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_9_io_i_mux_bus_0_1 = _FDPE_9_i_mux_bus_0_1_rev_T_11 | _GEN_2338; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_9_io_i_mux_bus_0_2 = _FDPE_9_i_mux_bus_0_2_rev_T_11 | _GEN_2344; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_9_io_i_mux_bus_0_3 = _FDPE_9_i_mux_bus_0_3_rev_T_11 | _GEN_2350; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_9_io_i_mux_bus_1_0 = _FDPE_9_i_mux_bus_1_0_rev_T_11 | _GEN_2356; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_9_io_i_mux_bus_1_1 = _FDPE_9_i_mux_bus_1_1_rev_T_11 | _GEN_2362; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_9_io_i_mux_bus_1_2 = _FDPE_9_i_mux_bus_1_2_rev_T_11 | _GEN_2368; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_9_io_i_mux_bus_2_0 = _FDPE_9_i_mux_bus_2_0_rev_T_11 | _GEN_2374; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_9_io_i_mux_bus_2_1 = _FDPE_9_i_mux_bus_2_1_rev_T_11 | _GEN_2380; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_9_io_i_mux_bus_3_0 = _FDPE_9_i_mux_bus_3_0_rev_T_11 | _GEN_2386; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_10_clock = clock;
  assign flexdpecom4_10_reset = reset;
  assign flexdpecom4_10_io_i_data_valid = 1'h1; // @[FlexDPU.scala 132:27 136:34]
  assign flexdpecom4_10_io_i_data_bus_0 = nonZeroValues_40[15:0]; // @[FlexDPU.scala 132:27 150:37]
  assign flexdpecom4_10_io_i_data_bus_1 = nonZeroValues_41[15:0]; // @[FlexDPU.scala 132:27 151:37]
  assign flexdpecom4_10_io_i_data_bus_2 = nonZeroValues_42[15:0]; // @[FlexDPU.scala 132:27 152:37]
  assign flexdpecom4_10_io_i_data_bus_3 = nonZeroValues_43[15:0]; // @[FlexDPU.scala 132:27 153:37]
  assign flexdpecom4_10_io_i_data_bus2_0 = MuxWrapper_10_Osrc_0[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_10_io_i_data_bus2_1 = MuxWrapper_10_Osrc_1[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_10_io_i_data_bus2_2 = MuxWrapper_10_Osrc_2[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_10_io_i_data_bus2_3 = MuxWrapper_10_Osrc_3[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_10_io_i_vn_0 = ivntop_io_o_vn_10_0; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_10_io_i_vn_1 = ivntop_io_o_vn_10_1; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_10_io_i_vn_2 = ivntop_io_o_vn_10_2; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_10_io_i_vn_3 = ivntop_io_o_vn_10_3; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_10_io_i_mux_bus_0_0 = _FDPE_10_i_mux_bus_0_0_rev_T_11 | _GEN_2392; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_10_io_i_mux_bus_0_1 = _FDPE_10_i_mux_bus_0_1_rev_T_11 | _GEN_2398; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_10_io_i_mux_bus_0_2 = _FDPE_10_i_mux_bus_0_2_rev_T_11 | _GEN_2404; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_10_io_i_mux_bus_0_3 = _FDPE_10_i_mux_bus_0_3_rev_T_11 | _GEN_2410; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_10_io_i_mux_bus_1_0 = _FDPE_10_i_mux_bus_1_0_rev_T_11 | _GEN_2416; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_10_io_i_mux_bus_1_1 = _FDPE_10_i_mux_bus_1_1_rev_T_11 | _GEN_2422; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_10_io_i_mux_bus_1_2 = _FDPE_10_i_mux_bus_1_2_rev_T_11 | _GEN_2428; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_10_io_i_mux_bus_2_0 = _FDPE_10_i_mux_bus_2_0_rev_T_11 | _GEN_2434; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_10_io_i_mux_bus_2_1 = _FDPE_10_i_mux_bus_2_1_rev_T_11 | _GEN_2440; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_10_io_i_mux_bus_3_0 = _FDPE_10_i_mux_bus_3_0_rev_T_11 | _GEN_2446; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_11_clock = clock;
  assign flexdpecom4_11_reset = reset;
  assign flexdpecom4_11_io_i_data_valid = 1'h1; // @[FlexDPU.scala 132:27 136:34]
  assign flexdpecom4_11_io_i_data_bus_0 = nonZeroValues_44[15:0]; // @[FlexDPU.scala 132:27 150:37]
  assign flexdpecom4_11_io_i_data_bus_1 = nonZeroValues_45[15:0]; // @[FlexDPU.scala 132:27 151:37]
  assign flexdpecom4_11_io_i_data_bus_2 = nonZeroValues_46[15:0]; // @[FlexDPU.scala 132:27 152:37]
  assign flexdpecom4_11_io_i_data_bus_3 = nonZeroValues_47[15:0]; // @[FlexDPU.scala 132:27 153:37]
  assign flexdpecom4_11_io_i_data_bus2_0 = MuxWrapper_11_Osrc_0[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_11_io_i_data_bus2_1 = MuxWrapper_11_Osrc_1[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_11_io_i_data_bus2_2 = MuxWrapper_11_Osrc_2[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_11_io_i_data_bus2_3 = MuxWrapper_11_Osrc_3[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_11_io_i_vn_0 = ivntop_io_o_vn_11_0; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_11_io_i_vn_1 = ivntop_io_o_vn_11_1; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_11_io_i_vn_2 = ivntop_io_o_vn_11_2; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_11_io_i_vn_3 = ivntop_io_o_vn_11_3; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_11_io_i_mux_bus_0_0 = _FDPE_11_i_mux_bus_0_0_rev_T_11 | _GEN_2452; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_11_io_i_mux_bus_0_1 = _FDPE_11_i_mux_bus_0_1_rev_T_11 | _GEN_2458; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_11_io_i_mux_bus_0_2 = _FDPE_11_i_mux_bus_0_2_rev_T_11 | _GEN_2464; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_11_io_i_mux_bus_0_3 = _FDPE_11_i_mux_bus_0_3_rev_T_11 | _GEN_2470; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_11_io_i_mux_bus_1_0 = _FDPE_11_i_mux_bus_1_0_rev_T_11 | _GEN_2476; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_11_io_i_mux_bus_1_1 = _FDPE_11_i_mux_bus_1_1_rev_T_11 | _GEN_2482; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_11_io_i_mux_bus_1_2 = _FDPE_11_i_mux_bus_1_2_rev_T_11 | _GEN_2488; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_11_io_i_mux_bus_2_0 = _FDPE_11_i_mux_bus_2_0_rev_T_11 | _GEN_2494; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_11_io_i_mux_bus_2_1 = _FDPE_11_i_mux_bus_2_1_rev_T_11 | _GEN_2500; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_11_io_i_mux_bus_3_0 = _FDPE_11_i_mux_bus_3_0_rev_T_11 | _GEN_2506; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_12_clock = clock;
  assign flexdpecom4_12_reset = reset;
  assign flexdpecom4_12_io_i_data_valid = 1'h1; // @[FlexDPU.scala 132:27 136:34]
  assign flexdpecom4_12_io_i_data_bus_0 = nonZeroValues_48[15:0]; // @[FlexDPU.scala 132:27 150:37]
  assign flexdpecom4_12_io_i_data_bus_1 = nonZeroValues_49[15:0]; // @[FlexDPU.scala 132:27 151:37]
  assign flexdpecom4_12_io_i_data_bus_2 = nonZeroValues_50[15:0]; // @[FlexDPU.scala 132:27 152:37]
  assign flexdpecom4_12_io_i_data_bus_3 = nonZeroValues_51[15:0]; // @[FlexDPU.scala 132:27 153:37]
  assign flexdpecom4_12_io_i_data_bus2_0 = MuxWrapper_12_Osrc_0[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_12_io_i_data_bus2_1 = MuxWrapper_12_Osrc_1[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_12_io_i_data_bus2_2 = MuxWrapper_12_Osrc_2[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_12_io_i_data_bus2_3 = MuxWrapper_12_Osrc_3[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_12_io_i_vn_0 = ivntop_io_o_vn_12_0; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_12_io_i_vn_1 = ivntop_io_o_vn_12_1; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_12_io_i_vn_2 = ivntop_io_o_vn_12_2; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_12_io_i_vn_3 = ivntop_io_o_vn_12_3; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_12_io_i_mux_bus_0_0 = _FDPE_12_i_mux_bus_0_0_rev_T_11 | _GEN_2512; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_12_io_i_mux_bus_0_1 = _FDPE_12_i_mux_bus_0_1_rev_T_11 | _GEN_2518; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_12_io_i_mux_bus_0_2 = _FDPE_12_i_mux_bus_0_2_rev_T_11 | _GEN_2524; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_12_io_i_mux_bus_0_3 = _FDPE_12_i_mux_bus_0_3_rev_T_11 | _GEN_2530; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_12_io_i_mux_bus_1_0 = _FDPE_12_i_mux_bus_1_0_rev_T_11 | _GEN_2536; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_12_io_i_mux_bus_1_1 = _FDPE_12_i_mux_bus_1_1_rev_T_11 | _GEN_2542; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_12_io_i_mux_bus_1_2 = _FDPE_12_i_mux_bus_1_2_rev_T_11 | _GEN_2548; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_12_io_i_mux_bus_2_0 = _FDPE_12_i_mux_bus_2_0_rev_T_11 | _GEN_2554; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_12_io_i_mux_bus_2_1 = _FDPE_12_i_mux_bus_2_1_rev_T_11 | _GEN_2560; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_12_io_i_mux_bus_3_0 = _FDPE_12_i_mux_bus_3_0_rev_T_11 | _GEN_2566; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_13_clock = clock;
  assign flexdpecom4_13_reset = reset;
  assign flexdpecom4_13_io_i_data_valid = 1'h1; // @[FlexDPU.scala 132:27 136:34]
  assign flexdpecom4_13_io_i_data_bus_0 = nonZeroValues_52[15:0]; // @[FlexDPU.scala 132:27 150:37]
  assign flexdpecom4_13_io_i_data_bus_1 = nonZeroValues_53[15:0]; // @[FlexDPU.scala 132:27 151:37]
  assign flexdpecom4_13_io_i_data_bus_2 = nonZeroValues_54[15:0]; // @[FlexDPU.scala 132:27 152:37]
  assign flexdpecom4_13_io_i_data_bus_3 = nonZeroValues_55[15:0]; // @[FlexDPU.scala 132:27 153:37]
  assign flexdpecom4_13_io_i_data_bus2_0 = MuxWrapper_13_Osrc_0[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_13_io_i_data_bus2_1 = MuxWrapper_13_Osrc_1[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_13_io_i_data_bus2_2 = MuxWrapper_13_Osrc_2[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_13_io_i_data_bus2_3 = MuxWrapper_13_Osrc_3[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_13_io_i_vn_0 = ivntop_io_o_vn_13_0; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_13_io_i_vn_1 = ivntop_io_o_vn_13_1; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_13_io_i_vn_2 = ivntop_io_o_vn_13_2; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_13_io_i_vn_3 = ivntop_io_o_vn_13_3; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_13_io_i_mux_bus_0_0 = _FDPE_13_i_mux_bus_0_0_rev_T_11 | _GEN_2572; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_13_io_i_mux_bus_0_1 = _FDPE_13_i_mux_bus_0_1_rev_T_11 | _GEN_2578; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_13_io_i_mux_bus_0_2 = _FDPE_13_i_mux_bus_0_2_rev_T_11 | _GEN_2584; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_13_io_i_mux_bus_0_3 = _FDPE_13_i_mux_bus_0_3_rev_T_11 | _GEN_2590; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_13_io_i_mux_bus_1_0 = _FDPE_13_i_mux_bus_1_0_rev_T_11 | _GEN_2596; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_13_io_i_mux_bus_1_1 = _FDPE_13_i_mux_bus_1_1_rev_T_11 | _GEN_2602; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_13_io_i_mux_bus_1_2 = _FDPE_13_i_mux_bus_1_2_rev_T_11 | _GEN_2608; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_13_io_i_mux_bus_2_0 = _FDPE_13_i_mux_bus_2_0_rev_T_11 | _GEN_2614; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_13_io_i_mux_bus_2_1 = _FDPE_13_i_mux_bus_2_1_rev_T_11 | _GEN_2620; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_13_io_i_mux_bus_3_0 = _FDPE_13_i_mux_bus_3_0_rev_T_11 | _GEN_2626; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_14_clock = clock;
  assign flexdpecom4_14_reset = reset;
  assign flexdpecom4_14_io_i_data_valid = 1'h1; // @[FlexDPU.scala 132:27 136:34]
  assign flexdpecom4_14_io_i_data_bus_0 = nonZeroValues_56[15:0]; // @[FlexDPU.scala 132:27 150:37]
  assign flexdpecom4_14_io_i_data_bus_1 = nonZeroValues_57[15:0]; // @[FlexDPU.scala 132:27 151:37]
  assign flexdpecom4_14_io_i_data_bus_2 = nonZeroValues_58[15:0]; // @[FlexDPU.scala 132:27 152:37]
  assign flexdpecom4_14_io_i_data_bus_3 = nonZeroValues_59[15:0]; // @[FlexDPU.scala 132:27 153:37]
  assign flexdpecom4_14_io_i_data_bus2_0 = MuxWrapper_14_Osrc_0[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_14_io_i_data_bus2_1 = MuxWrapper_14_Osrc_1[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_14_io_i_data_bus2_2 = MuxWrapper_14_Osrc_2[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_14_io_i_data_bus2_3 = MuxWrapper_14_Osrc_3[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_14_io_i_vn_0 = ivntop_io_o_vn_14_0; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_14_io_i_vn_1 = ivntop_io_o_vn_14_1; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_14_io_i_vn_2 = ivntop_io_o_vn_14_2; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_14_io_i_vn_3 = ivntop_io_o_vn_14_3; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_14_io_i_mux_bus_0_0 = _FDPE_14_i_mux_bus_0_0_rev_T_11 | _GEN_2632; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_14_io_i_mux_bus_0_1 = _FDPE_14_i_mux_bus_0_1_rev_T_11 | _GEN_2638; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_14_io_i_mux_bus_0_2 = _FDPE_14_i_mux_bus_0_2_rev_T_11 | _GEN_2644; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_14_io_i_mux_bus_0_3 = _FDPE_14_i_mux_bus_0_3_rev_T_11 | _GEN_2650; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_14_io_i_mux_bus_1_0 = _FDPE_14_i_mux_bus_1_0_rev_T_11 | _GEN_2656; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_14_io_i_mux_bus_1_1 = _FDPE_14_i_mux_bus_1_1_rev_T_11 | _GEN_2662; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_14_io_i_mux_bus_1_2 = _FDPE_14_i_mux_bus_1_2_rev_T_11 | _GEN_2668; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_14_io_i_mux_bus_2_0 = _FDPE_14_i_mux_bus_2_0_rev_T_11 | _GEN_2674; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_14_io_i_mux_bus_2_1 = _FDPE_14_i_mux_bus_2_1_rev_T_11 | _GEN_2680; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_14_io_i_mux_bus_3_0 = _FDPE_14_i_mux_bus_3_0_rev_T_11 | _GEN_2686; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_15_clock = clock;
  assign flexdpecom4_15_reset = reset;
  assign flexdpecom4_15_io_i_data_valid = 1'h1; // @[FlexDPU.scala 132:27 136:34]
  assign flexdpecom4_15_io_i_data_bus_0 = nonZeroValues_60[15:0]; // @[FlexDPU.scala 132:27 150:37]
  assign flexdpecom4_15_io_i_data_bus_1 = nonZeroValues_61[15:0]; // @[FlexDPU.scala 132:27 151:37]
  assign flexdpecom4_15_io_i_data_bus_2 = nonZeroValues_62[15:0]; // @[FlexDPU.scala 132:27 152:37]
  assign flexdpecom4_15_io_i_data_bus_3 = nonZeroValues_63[15:0]; // @[FlexDPU.scala 132:27 153:37]
  assign flexdpecom4_15_io_i_data_bus2_0 = MuxWrapper_15_Osrc_0[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_15_io_i_data_bus2_1 = MuxWrapper_15_Osrc_1[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_15_io_i_data_bus2_2 = MuxWrapper_15_Osrc_2[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_15_io_i_data_bus2_3 = MuxWrapper_15_Osrc_3[15:0]; // @[FlexDPU.scala 132:27 144:33]
  assign flexdpecom4_15_io_i_vn_0 = ivntop_io_o_vn_15_0; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_15_io_i_vn_1 = ivntop_io_o_vn_15_1; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_15_io_i_vn_2 = ivntop_io_o_vn_15_2; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_15_io_i_vn_3 = ivntop_io_o_vn_15_3; // @[FlexDPU.scala 132:27 139:37]
  assign flexdpecom4_15_io_i_mux_bus_0_0 = _FDPE_15_i_mux_bus_0_0_rev_T_11 | _GEN_2692; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_15_io_i_mux_bus_0_1 = _FDPE_15_i_mux_bus_0_1_rev_T_11 | _GEN_2698; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_15_io_i_mux_bus_0_2 = _FDPE_15_i_mux_bus_0_2_rev_T_11 | _GEN_2704; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_15_io_i_mux_bus_0_3 = _FDPE_15_i_mux_bus_0_3_rev_T_11 | _GEN_2710; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_15_io_i_mux_bus_1_0 = _FDPE_15_i_mux_bus_1_0_rev_T_11 | _GEN_2716; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_15_io_i_mux_bus_1_1 = _FDPE_15_i_mux_bus_1_1_rev_T_11 | _GEN_2722; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_15_io_i_mux_bus_1_2 = _FDPE_15_i_mux_bus_1_2_rev_T_11 | _GEN_2728; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_15_io_i_mux_bus_2_0 = _FDPE_15_i_mux_bus_2_0_rev_T_11 | _GEN_2734; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_15_io_i_mux_bus_2_1 = _FDPE_15_i_mux_bus_2_1_rev_T_11 | _GEN_2740; // @[FlexDPU.scala 68:17]
  assign flexdpecom4_15_io_i_mux_bus_3_0 = _FDPE_15_i_mux_bus_3_0_rev_T_11 | _GEN_2746; // @[FlexDPU.scala 68:17]
  always @(posedge clock) begin
    if (5'h0 < remainingDistribution) begin // @[FlexDPU.scala 25:29]
      used_FlexDPE_0 <= _used_FlexDPE_0_T_2;
    end else begin
      used_FlexDPE_0 <= equalDistribution;
    end
    if (5'h1 < remainingDistribution) begin // @[FlexDPU.scala 25:29]
      used_FlexDPE_1 <= _used_FlexDPE_0_T_2;
    end else begin
      used_FlexDPE_1 <= equalDistribution;
    end
    if (5'h2 < remainingDistribution) begin // @[FlexDPU.scala 25:29]
      used_FlexDPE_2 <= _used_FlexDPE_0_T_2;
    end else begin
      used_FlexDPE_2 <= equalDistribution;
    end
    if (5'h3 < remainingDistribution) begin // @[FlexDPU.scala 25:29]
      used_FlexDPE_3 <= _used_FlexDPE_0_T_2;
    end else begin
      used_FlexDPE_3 <= equalDistribution;
    end
    if (5'h4 < remainingDistribution) begin // @[FlexDPU.scala 25:29]
      used_FlexDPE_4 <= _used_FlexDPE_0_T_2;
    end else begin
      used_FlexDPE_4 <= equalDistribution;
    end
    if (5'h5 < remainingDistribution) begin // @[FlexDPU.scala 25:29]
      used_FlexDPE_5 <= _used_FlexDPE_0_T_2;
    end else begin
      used_FlexDPE_5 <= equalDistribution;
    end
    if (5'h6 < remainingDistribution) begin // @[FlexDPU.scala 25:29]
      used_FlexDPE_6 <= _used_FlexDPE_0_T_2;
    end else begin
      used_FlexDPE_6 <= equalDistribution;
    end
    if (5'h7 < remainingDistribution) begin // @[FlexDPU.scala 25:29]
      used_FlexDPE_7 <= _used_FlexDPE_0_T_2;
    end else begin
      used_FlexDPE_7 <= equalDistribution;
    end
    if (5'h8 < remainingDistribution) begin // @[FlexDPU.scala 25:29]
      used_FlexDPE_8 <= _used_FlexDPE_0_T_2;
    end else begin
      used_FlexDPE_8 <= equalDistribution;
    end
    if (5'h9 < remainingDistribution) begin // @[FlexDPU.scala 25:29]
      used_FlexDPE_9 <= _used_FlexDPE_0_T_2;
    end else begin
      used_FlexDPE_9 <= equalDistribution;
    end
    if (5'ha < remainingDistribution) begin // @[FlexDPU.scala 25:29]
      used_FlexDPE_10 <= _used_FlexDPE_0_T_2;
    end else begin
      used_FlexDPE_10 <= equalDistribution;
    end
    if (5'hb < remainingDistribution) begin // @[FlexDPU.scala 25:29]
      used_FlexDPE_11 <= _used_FlexDPE_0_T_2;
    end else begin
      used_FlexDPE_11 <= equalDistribution;
    end
    if (5'hc < remainingDistribution) begin // @[FlexDPU.scala 25:29]
      used_FlexDPE_12 <= _used_FlexDPE_0_T_2;
    end else begin
      used_FlexDPE_12 <= equalDistribution;
    end
    if (5'hd < remainingDistribution) begin // @[FlexDPU.scala 25:29]
      used_FlexDPE_13 <= _used_FlexDPE_0_T_2;
    end else begin
      used_FlexDPE_13 <= equalDistribution;
    end
    if (5'he < remainingDistribution) begin // @[FlexDPU.scala 25:29]
      used_FlexDPE_14 <= _used_FlexDPE_0_T_2;
    end else begin
      used_FlexDPE_14 <= equalDistribution;
    end
    if (5'hf < remainingDistribution) begin // @[FlexDPU.scala 25:29]
      used_FlexDPE_15 <= _used_FlexDPE_0_T_2;
    end else begin
      used_FlexDPE_15 <= equalDistribution;
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_0 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'h0 == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_0 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_1 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'h1 == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_1 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_2 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'h2 == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_2 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_3 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'h3 == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_3 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_4 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'h4 == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_4 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_5 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'h5 == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_5 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_6 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'h6 == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_6 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_7 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'h7 == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_7 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_8 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'h8 == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_8 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_9 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'h9 == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_9 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_10 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'ha == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_10 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_11 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'hb == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_11 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_12 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'hc == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_12 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_13 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'hd == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_13 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_14 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'he == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_14 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_15 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'hf == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_15 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_16 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'h10 == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_16 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_17 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'h11 == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_17 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_18 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'h12 == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_18 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_19 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'h13 == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_19 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_20 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'h14 == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_20 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_21 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'h15 == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_21 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_22 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'h16 == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_22 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_23 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'h17 == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_23 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_24 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'h18 == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_24 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_25 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'h19 == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_25 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_26 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'h1a == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_26 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_27 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'h1b == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_27 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_28 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'h1c == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_28 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_29 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'h1d == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_29 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_30 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'h1e == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_30 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_31 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'h1f == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_31 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_32 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'h20 == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_32 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_33 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'h21 == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_33 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_34 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'h22 == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_34 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_35 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'h23 == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_35 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_36 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'h24 == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_36 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_37 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'h25 == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_37 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_38 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'h26 == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_38 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_39 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'h27 == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_39 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_40 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'h28 == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_40 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_41 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'h29 == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_41 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_42 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'h2a == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_42 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_43 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'h2b == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_43 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_44 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'h2c == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_44 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_45 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'h2d == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_45 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_46 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'h2e == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_46 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_47 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'h2f == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_47 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_48 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'h30 == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_48 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_49 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'h31 == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_49 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_50 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'h32 == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_50 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_51 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'h33 == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_51 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_52 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'h34 == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_52 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_53 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'h35 == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_53 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_54 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'h36 == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_54 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_55 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'h37 == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_55 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_56 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'h38 == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_56 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_57 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'h39 == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_57 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_58 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'h3a == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_58 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_59 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'h3b == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_59 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_60 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'h3c == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_60 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_61 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'h3d == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_61 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_62 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'h3e == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_62 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 31:32]
      nonZeroValues_63 <= 32'h0; // @[FlexDPU.scala 31:32]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      if (6'h3f == index[5:0]) begin // @[FlexDPU.scala 39:30]
        nonZeroValues_63 <= _nonZeroValues_T_3; // @[FlexDPU.scala 39:30]
      end
    end
    if (reset) begin // @[FlexDPU.scala 32:24]
      index <= 32'h0; // @[FlexDPU.scala 32:24]
    end else if (_GEN_63 != 16'h0) begin // @[FlexDPU.scala 38:54]
      index <= _index_T_1; // @[FlexDPU.scala 40:15]
    end
    if (reset) begin // @[FlexDPU.scala 33:24]
      iloop <= 32'h0; // @[FlexDPU.scala 33:24]
    end else if (iloop < 32'h7 & _Statvalid_T_1) begin // @[FlexDPU.scala 43:77]
      iloop <= _iloop_T_1; // @[FlexDPU.scala 44:15]
    end
    if (reset) begin // @[FlexDPU.scala 34:24]
      jloop <= 32'h0; // @[FlexDPU.scala 34:24]
    end else if (iloop <= 32'h7 & jloop < 32'h7) begin // @[FlexDPU.scala 47:76]
      jloop <= _jloop_T_1; // @[FlexDPU.scala 48:15]
    end else if (!(_Statvalid_T_2)) begin // @[FlexDPU.scala 49:83]
      jloop <= 32'h0; // @[FlexDPU.scala 52:15]
    end
    if (reset) begin // @[FlexDPU.scala 35:28]
      Statvalid <= 1'h0; // @[FlexDPU.scala 35:28]
    end else begin
      Statvalid <= iloop == 32'h7 & jloop == 32'h7; // @[FlexDPU.scala 37:15]
    end
    if (reset) begin // @[FlexDPU.scala 61:33]
      PF1_Stream_Col_0 <= 32'h0; // @[FlexDPU.scala 61:33]
    end else if (Statvalid & check) begin // @[FlexDPU.scala 112:29]
      PF1_Stream_Col_0 <= {{16'd0}, _GEN_274}; // @[FlexDPU.scala 189:31]
    end
    if (reset) begin // @[FlexDPU.scala 61:33]
      PF1_Stream_Col_1 <= 32'h0; // @[FlexDPU.scala 61:33]
    end else if (Statvalid & check) begin // @[FlexDPU.scala 112:29]
      PF1_Stream_Col_1 <= {{16'd0}, _GEN_282}; // @[FlexDPU.scala 189:31]
    end
    if (reset) begin // @[FlexDPU.scala 61:33]
      PF1_Stream_Col_2 <= 32'h0; // @[FlexDPU.scala 61:33]
    end else if (Statvalid & check) begin // @[FlexDPU.scala 112:29]
      PF1_Stream_Col_2 <= {{16'd0}, _GEN_290}; // @[FlexDPU.scala 189:31]
    end
    if (reset) begin // @[FlexDPU.scala 61:33]
      PF1_Stream_Col_3 <= 32'h0; // @[FlexDPU.scala 61:33]
    end else if (Statvalid & check) begin // @[FlexDPU.scala 112:29]
      PF1_Stream_Col_3 <= {{16'd0}, _GEN_298}; // @[FlexDPU.scala 189:31]
    end
    if (reset) begin // @[FlexDPU.scala 61:33]
      PF1_Stream_Col_4 <= 32'h0; // @[FlexDPU.scala 61:33]
    end else if (Statvalid & check) begin // @[FlexDPU.scala 112:29]
      PF1_Stream_Col_4 <= {{16'd0}, _GEN_306}; // @[FlexDPU.scala 189:31]
    end
    if (reset) begin // @[FlexDPU.scala 61:33]
      PF1_Stream_Col_5 <= 32'h0; // @[FlexDPU.scala 61:33]
    end else if (Statvalid & check) begin // @[FlexDPU.scala 112:29]
      PF1_Stream_Col_5 <= {{16'd0}, _GEN_314}; // @[FlexDPU.scala 189:31]
    end
    if (reset) begin // @[FlexDPU.scala 61:33]
      PF1_Stream_Col_6 <= 32'h0; // @[FlexDPU.scala 61:33]
    end else if (Statvalid & check) begin // @[FlexDPU.scala 112:29]
      PF1_Stream_Col_6 <= {{16'd0}, _GEN_322}; // @[FlexDPU.scala 189:31]
    end
    if (reset) begin // @[FlexDPU.scala 61:33]
      PF1_Stream_Col_7 <= 32'h0; // @[FlexDPU.scala 61:33]
    end else if (Statvalid & check) begin // @[FlexDPU.scala 112:29]
      PF1_Stream_Col_7 <= {{16'd0}, _GEN_330}; // @[FlexDPU.scala 189:31]
    end
    if (reset) begin // @[FlexDPU.scala 62:30]
      ModuleIndex <= 32'h0; // @[FlexDPU.scala 62:30]
    end else if (Statvalid & check) begin // @[FlexDPU.scala 112:29]
      if (!(ModuleIndex == 32'h7 & PF_0_PF_Valid)) begin // @[FlexDPU.scala 182:71]
        if (PF_0_PF_Valid) begin // @[FlexDPU.scala 177:29]
          ModuleIndex <= _ModuleIndex_T_1; // @[FlexDPU.scala 179:25]
        end
      end
    end
    if (reset) begin // @[FlexDPU.scala 99:24]
      delay <= 32'h0; // @[FlexDPU.scala 99:24]
    end else if (!(ivntop_io_ProcessValid)) begin // @[FlexDPU.scala 104:29]
      if (delay < 32'hbb8) begin // @[FlexDPU.scala 106:32]
        delay <= _delay_T_1; // @[FlexDPU.scala 107:11]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  used_FlexDPE_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  used_FlexDPE_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  used_FlexDPE_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  used_FlexDPE_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  used_FlexDPE_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  used_FlexDPE_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  used_FlexDPE_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  used_FlexDPE_7 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  used_FlexDPE_8 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  used_FlexDPE_9 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  used_FlexDPE_10 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  used_FlexDPE_11 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  used_FlexDPE_12 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  used_FlexDPE_13 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  used_FlexDPE_14 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  used_FlexDPE_15 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  nonZeroValues_0 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  nonZeroValues_1 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  nonZeroValues_2 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  nonZeroValues_3 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  nonZeroValues_4 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  nonZeroValues_5 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  nonZeroValues_6 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  nonZeroValues_7 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  nonZeroValues_8 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  nonZeroValues_9 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  nonZeroValues_10 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  nonZeroValues_11 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  nonZeroValues_12 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  nonZeroValues_13 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  nonZeroValues_14 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  nonZeroValues_15 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  nonZeroValues_16 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  nonZeroValues_17 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  nonZeroValues_18 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  nonZeroValues_19 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  nonZeroValues_20 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  nonZeroValues_21 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  nonZeroValues_22 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  nonZeroValues_23 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  nonZeroValues_24 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  nonZeroValues_25 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  nonZeroValues_26 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  nonZeroValues_27 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  nonZeroValues_28 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  nonZeroValues_29 = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  nonZeroValues_30 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  nonZeroValues_31 = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  nonZeroValues_32 = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  nonZeroValues_33 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  nonZeroValues_34 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  nonZeroValues_35 = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  nonZeroValues_36 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  nonZeroValues_37 = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  nonZeroValues_38 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  nonZeroValues_39 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  nonZeroValues_40 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  nonZeroValues_41 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  nonZeroValues_42 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  nonZeroValues_43 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  nonZeroValues_44 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  nonZeroValues_45 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  nonZeroValues_46 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  nonZeroValues_47 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  nonZeroValues_48 = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  nonZeroValues_49 = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  nonZeroValues_50 = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  nonZeroValues_51 = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  nonZeroValues_52 = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  nonZeroValues_53 = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  nonZeroValues_54 = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  nonZeroValues_55 = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  nonZeroValues_56 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  nonZeroValues_57 = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  nonZeroValues_58 = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  nonZeroValues_59 = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  nonZeroValues_60 = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  nonZeroValues_61 = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  nonZeroValues_62 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  nonZeroValues_63 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  index = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  iloop = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  jloop = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  Statvalid = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  PF1_Stream_Col_0 = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  PF1_Stream_Col_1 = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  PF1_Stream_Col_2 = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  PF1_Stream_Col_3 = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  PF1_Stream_Col_4 = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  PF1_Stream_Col_5 = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  PF1_Stream_Col_6 = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  PF1_Stream_Col_7 = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  ModuleIndex = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  delay = _RAND_93[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Top(
  input         clock,
  input         reset,
  input  [31:0] io_Stationary_matrix_0_0,
  input  [31:0] io_Stationary_matrix_0_1,
  input  [31:0] io_Stationary_matrix_0_2,
  input  [31:0] io_Stationary_matrix_0_3,
  input  [31:0] io_Stationary_matrix_0_4,
  input  [31:0] io_Stationary_matrix_0_5,
  input  [31:0] io_Stationary_matrix_0_6,
  input  [31:0] io_Stationary_matrix_0_7,
  input  [31:0] io_Stationary_matrix_1_0,
  input  [31:0] io_Stationary_matrix_1_1,
  input  [31:0] io_Stationary_matrix_1_2,
  input  [31:0] io_Stationary_matrix_1_3,
  input  [31:0] io_Stationary_matrix_1_4,
  input  [31:0] io_Stationary_matrix_1_5,
  input  [31:0] io_Stationary_matrix_1_6,
  input  [31:0] io_Stationary_matrix_1_7,
  input  [31:0] io_Stationary_matrix_2_0,
  input  [31:0] io_Stationary_matrix_2_1,
  input  [31:0] io_Stationary_matrix_2_2,
  input  [31:0] io_Stationary_matrix_2_3,
  input  [31:0] io_Stationary_matrix_2_4,
  input  [31:0] io_Stationary_matrix_2_5,
  input  [31:0] io_Stationary_matrix_2_6,
  input  [31:0] io_Stationary_matrix_2_7,
  input  [31:0] io_Stationary_matrix_3_0,
  input  [31:0] io_Stationary_matrix_3_1,
  input  [31:0] io_Stationary_matrix_3_2,
  input  [31:0] io_Stationary_matrix_3_3,
  input  [31:0] io_Stationary_matrix_3_4,
  input  [31:0] io_Stationary_matrix_3_5,
  input  [31:0] io_Stationary_matrix_3_6,
  input  [31:0] io_Stationary_matrix_3_7,
  input  [31:0] io_Stationary_matrix_4_0,
  input  [31:0] io_Stationary_matrix_4_1,
  input  [31:0] io_Stationary_matrix_4_2,
  input  [31:0] io_Stationary_matrix_4_3,
  input  [31:0] io_Stationary_matrix_4_4,
  input  [31:0] io_Stationary_matrix_4_5,
  input  [31:0] io_Stationary_matrix_4_6,
  input  [31:0] io_Stationary_matrix_4_7,
  input  [31:0] io_Stationary_matrix_5_0,
  input  [31:0] io_Stationary_matrix_5_1,
  input  [31:0] io_Stationary_matrix_5_2,
  input  [31:0] io_Stationary_matrix_5_3,
  input  [31:0] io_Stationary_matrix_5_4,
  input  [31:0] io_Stationary_matrix_5_5,
  input  [31:0] io_Stationary_matrix_5_6,
  input  [31:0] io_Stationary_matrix_5_7,
  input  [31:0] io_Stationary_matrix_6_0,
  input  [31:0] io_Stationary_matrix_6_1,
  input  [31:0] io_Stationary_matrix_6_2,
  input  [31:0] io_Stationary_matrix_6_3,
  input  [31:0] io_Stationary_matrix_6_4,
  input  [31:0] io_Stationary_matrix_6_5,
  input  [31:0] io_Stationary_matrix_6_6,
  input  [31:0] io_Stationary_matrix_6_7,
  input  [31:0] io_Stationary_matrix_7_0,
  input  [31:0] io_Stationary_matrix_7_1,
  input  [31:0] io_Stationary_matrix_7_2,
  input  [31:0] io_Stationary_matrix_7_3,
  input  [31:0] io_Stationary_matrix_7_4,
  input  [31:0] io_Stationary_matrix_7_5,
  input  [31:0] io_Stationary_matrix_7_6,
  input  [31:0] io_Stationary_matrix_7_7,
  input  [31:0] io_Streaming_matrix_0_0,
  input  [31:0] io_Streaming_matrix_0_1,
  input  [31:0] io_Streaming_matrix_0_2,
  input  [31:0] io_Streaming_matrix_0_3,
  input  [31:0] io_Streaming_matrix_0_4,
  input  [31:0] io_Streaming_matrix_0_5,
  input  [31:0] io_Streaming_matrix_0_6,
  input  [31:0] io_Streaming_matrix_0_7,
  input  [31:0] io_Streaming_matrix_1_0,
  input  [31:0] io_Streaming_matrix_1_1,
  input  [31:0] io_Streaming_matrix_1_2,
  input  [31:0] io_Streaming_matrix_1_3,
  input  [31:0] io_Streaming_matrix_1_4,
  input  [31:0] io_Streaming_matrix_1_5,
  input  [31:0] io_Streaming_matrix_1_6,
  input  [31:0] io_Streaming_matrix_1_7,
  input  [31:0] io_Streaming_matrix_2_0,
  input  [31:0] io_Streaming_matrix_2_1,
  input  [31:0] io_Streaming_matrix_2_2,
  input  [31:0] io_Streaming_matrix_2_3,
  input  [31:0] io_Streaming_matrix_2_4,
  input  [31:0] io_Streaming_matrix_2_5,
  input  [31:0] io_Streaming_matrix_2_6,
  input  [31:0] io_Streaming_matrix_2_7,
  input  [31:0] io_Streaming_matrix_3_0,
  input  [31:0] io_Streaming_matrix_3_1,
  input  [31:0] io_Streaming_matrix_3_2,
  input  [31:0] io_Streaming_matrix_3_3,
  input  [31:0] io_Streaming_matrix_3_4,
  input  [31:0] io_Streaming_matrix_3_5,
  input  [31:0] io_Streaming_matrix_3_6,
  input  [31:0] io_Streaming_matrix_3_7,
  input  [31:0] io_Streaming_matrix_4_0,
  input  [31:0] io_Streaming_matrix_4_1,
  input  [31:0] io_Streaming_matrix_4_2,
  input  [31:0] io_Streaming_matrix_4_3,
  input  [31:0] io_Streaming_matrix_4_4,
  input  [31:0] io_Streaming_matrix_4_5,
  input  [31:0] io_Streaming_matrix_4_6,
  input  [31:0] io_Streaming_matrix_4_7,
  input  [31:0] io_Streaming_matrix_5_0,
  input  [31:0] io_Streaming_matrix_5_1,
  input  [31:0] io_Streaming_matrix_5_2,
  input  [31:0] io_Streaming_matrix_5_3,
  input  [31:0] io_Streaming_matrix_5_4,
  input  [31:0] io_Streaming_matrix_5_5,
  input  [31:0] io_Streaming_matrix_5_6,
  input  [31:0] io_Streaming_matrix_5_7,
  input  [31:0] io_Streaming_matrix_6_0,
  input  [31:0] io_Streaming_matrix_6_1,
  input  [31:0] io_Streaming_matrix_6_2,
  input  [31:0] io_Streaming_matrix_6_3,
  input  [31:0] io_Streaming_matrix_6_4,
  input  [31:0] io_Streaming_matrix_6_5,
  input  [31:0] io_Streaming_matrix_6_6,
  input  [31:0] io_Streaming_matrix_6_7,
  input  [31:0] io_Streaming_matrix_7_0,
  input  [31:0] io_Streaming_matrix_7_1,
  input  [31:0] io_Streaming_matrix_7_2,
  input  [31:0] io_Streaming_matrix_7_3,
  input  [31:0] io_Streaming_matrix_7_4,
  input  [31:0] io_Streaming_matrix_7_5,
  input  [31:0] io_Streaming_matrix_7_6,
  input  [31:0] io_Streaming_matrix_7_7,
  output [31:0] io_Third_Matrix_0_0,
  output [31:0] io_Third_Matrix_0_1,
  output [31:0] io_Third_Matrix_0_2,
  output [31:0] io_Third_Matrix_0_3,
  output [31:0] io_Third_Matrix_0_4,
  output [31:0] io_Third_Matrix_0_5,
  output [31:0] io_Third_Matrix_0_6,
  output [31:0] io_Third_Matrix_0_7,
  output [31:0] io_Third_Matrix_1_0,
  output [31:0] io_Third_Matrix_1_1,
  output [31:0] io_Third_Matrix_1_2,
  output [31:0] io_Third_Matrix_1_3,
  output [31:0] io_Third_Matrix_1_4,
  output [31:0] io_Third_Matrix_1_5,
  output [31:0] io_Third_Matrix_1_6,
  output [31:0] io_Third_Matrix_1_7,
  output [31:0] io_Third_Matrix_2_0,
  output [31:0] io_Third_Matrix_2_1,
  output [31:0] io_Third_Matrix_2_2,
  output [31:0] io_Third_Matrix_2_3,
  output [31:0] io_Third_Matrix_2_4,
  output [31:0] io_Third_Matrix_2_5,
  output [31:0] io_Third_Matrix_2_6,
  output [31:0] io_Third_Matrix_2_7,
  output [31:0] io_Third_Matrix_3_0,
  output [31:0] io_Third_Matrix_3_1,
  output [31:0] io_Third_Matrix_3_2,
  output [31:0] io_Third_Matrix_3_3,
  output [31:0] io_Third_Matrix_3_4,
  output [31:0] io_Third_Matrix_3_5,
  output [31:0] io_Third_Matrix_3_6,
  output [31:0] io_Third_Matrix_3_7,
  output [31:0] io_Third_Matrix_4_0,
  output [31:0] io_Third_Matrix_4_1,
  output [31:0] io_Third_Matrix_4_2,
  output [31:0] io_Third_Matrix_4_3,
  output [31:0] io_Third_Matrix_4_4,
  output [31:0] io_Third_Matrix_4_5,
  output [31:0] io_Third_Matrix_4_6,
  output [31:0] io_Third_Matrix_4_7,
  output [31:0] io_Third_Matrix_5_0,
  output [31:0] io_Third_Matrix_5_1,
  output [31:0] io_Third_Matrix_5_2,
  output [31:0] io_Third_Matrix_5_3,
  output [31:0] io_Third_Matrix_5_4,
  output [31:0] io_Third_Matrix_5_5,
  output [31:0] io_Third_Matrix_5_6,
  output [31:0] io_Third_Matrix_5_7,
  output [31:0] io_Third_Matrix_6_0,
  output [31:0] io_Third_Matrix_6_1,
  output [31:0] io_Third_Matrix_6_2,
  output [31:0] io_Third_Matrix_6_3,
  output [31:0] io_Third_Matrix_6_4,
  output [31:0] io_Third_Matrix_6_5,
  output [31:0] io_Third_Matrix_6_6,
  output [31:0] io_Third_Matrix_6_7,
  output [31:0] io_Third_Matrix_7_0,
  output [31:0] io_Third_Matrix_7_1,
  output [31:0] io_Third_Matrix_7_2,
  output [31:0] io_Third_Matrix_7_3,
  output [31:0] io_Third_Matrix_7_4,
  output [31:0] io_Third_Matrix_7_5,
  output [31:0] io_Third_Matrix_7_6,
  output [31:0] io_Third_Matrix_7_7
);
  wire  PreProcessor_clock; // @[TOP.scala 14:30]
  wire  PreProcessor_reset; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_0_0; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_0_1; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_0_2; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_0_3; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_0_4; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_0_5; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_0_6; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_0_7; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_1_0; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_1_1; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_1_2; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_1_3; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_1_4; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_1_5; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_1_6; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_1_7; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_2_0; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_2_1; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_2_2; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_2_3; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_2_4; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_2_5; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_2_6; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_2_7; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_3_0; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_3_1; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_3_2; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_3_3; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_3_4; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_3_5; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_3_6; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_3_7; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_4_0; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_4_1; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_4_2; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_4_3; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_4_4; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_4_5; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_4_6; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_4_7; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_5_0; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_5_1; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_5_2; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_5_3; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_5_4; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_5_5; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_5_6; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_5_7; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_6_0; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_6_1; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_6_2; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_6_3; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_6_4; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_6_5; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_6_6; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_6_7; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_7_0; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_7_1; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_7_2; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_7_3; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_7_4; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_7_5; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_7_6; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat1_7_7; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_0_0; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_0_1; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_0_2; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_0_3; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_0_4; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_0_5; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_0_6; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_0_7; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_1_0; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_1_1; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_1_2; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_1_3; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_1_4; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_1_5; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_1_6; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_1_7; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_2_0; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_2_1; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_2_2; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_2_3; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_2_4; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_2_5; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_2_6; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_2_7; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_3_0; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_3_1; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_3_2; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_3_3; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_3_4; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_3_5; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_3_6; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_3_7; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_4_0; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_4_1; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_4_2; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_4_3; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_4_4; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_4_5; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_4_6; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_4_7; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_5_0; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_5_1; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_5_2; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_5_3; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_5_4; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_5_5; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_5_6; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_5_7; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_6_0; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_6_1; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_6_2; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_6_3; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_6_4; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_6_5; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_6_6; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_6_7; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_7_0; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_7_1; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_7_2; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_7_3; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_7_4; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_7_5; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_7_6; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_mat2_7_7; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_0_0; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_0_1; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_0_2; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_0_3; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_0_4; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_0_5; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_0_6; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_0_7; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_1_0; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_1_1; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_1_2; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_1_3; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_1_4; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_1_5; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_1_6; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_1_7; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_2_0; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_2_1; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_2_2; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_2_3; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_2_4; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_2_5; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_2_6; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_2_7; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_3_0; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_3_1; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_3_2; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_3_3; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_3_4; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_3_5; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_3_6; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_3_7; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_4_0; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_4_1; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_4_2; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_4_3; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_4_4; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_4_5; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_4_6; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_4_7; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_5_0; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_5_1; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_5_2; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_5_3; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_5_4; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_5_5; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_5_6; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_5_7; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_6_0; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_6_1; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_6_2; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_6_3; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_6_4; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_6_5; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_6_6; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_6_7; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_7_0; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_7_1; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_7_2; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_7_3; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_7_4; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_7_5; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_7_6; // @[TOP.scala 14:30]
  wire [15:0] PreProcessor_io_compressedBitmap_7_7; // @[TOP.scala 14:30]
  wire  FDPU_clock; // @[TOP.scala 25:26]
  wire  FDPU_reset; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_0_0; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_0_1; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_0_2; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_0_3; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_0_4; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_0_5; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_0_6; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_0_7; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_1_0; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_1_1; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_1_2; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_1_3; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_1_4; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_1_5; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_1_6; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_1_7; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_2_0; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_2_1; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_2_2; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_2_3; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_2_4; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_2_5; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_2_6; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_2_7; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_3_0; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_3_1; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_3_2; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_3_3; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_3_4; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_3_5; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_3_6; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_3_7; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_4_0; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_4_1; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_4_2; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_4_3; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_4_4; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_4_5; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_4_6; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_4_7; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_5_0; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_5_1; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_5_2; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_5_3; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_5_4; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_5_5; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_5_6; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_5_7; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_6_0; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_6_1; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_6_2; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_6_3; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_6_4; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_6_5; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_6_6; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_6_7; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_7_0; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_7_1; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_7_2; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_7_3; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_7_4; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_7_5; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_7_6; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Stationary_matrix_7_7; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_0_0; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_0_1; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_0_2; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_0_3; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_0_4; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_0_5; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_0_6; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_0_7; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_1_0; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_1_1; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_1_2; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_1_3; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_1_4; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_1_5; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_1_6; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_1_7; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_2_0; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_2_1; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_2_2; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_2_3; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_2_4; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_2_5; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_2_6; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_2_7; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_3_0; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_3_1; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_3_2; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_3_3; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_3_4; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_3_5; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_3_6; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_3_7; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_4_0; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_4_1; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_4_2; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_4_3; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_4_4; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_4_5; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_4_6; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_4_7; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_5_0; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_5_1; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_5_2; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_5_3; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_5_4; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_5_5; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_5_6; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_5_7; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_6_0; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_6_1; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_6_2; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_6_3; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_6_4; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_6_5; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_6_6; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_6_7; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_7_0; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_7_1; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_7_2; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_7_3; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_7_4; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_7_5; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_7_6; // @[TOP.scala 25:26]
  wire [15:0] FDPU_io_Streaming_matrix_7_7; // @[TOP.scala 25:26]
  Regor PreProcessor ( // @[TOP.scala 14:30]
    .clock(PreProcessor_clock),
    .reset(PreProcessor_reset),
    .io_mat1_0_0(PreProcessor_io_mat1_0_0),
    .io_mat1_0_1(PreProcessor_io_mat1_0_1),
    .io_mat1_0_2(PreProcessor_io_mat1_0_2),
    .io_mat1_0_3(PreProcessor_io_mat1_0_3),
    .io_mat1_0_4(PreProcessor_io_mat1_0_4),
    .io_mat1_0_5(PreProcessor_io_mat1_0_5),
    .io_mat1_0_6(PreProcessor_io_mat1_0_6),
    .io_mat1_0_7(PreProcessor_io_mat1_0_7),
    .io_mat1_1_0(PreProcessor_io_mat1_1_0),
    .io_mat1_1_1(PreProcessor_io_mat1_1_1),
    .io_mat1_1_2(PreProcessor_io_mat1_1_2),
    .io_mat1_1_3(PreProcessor_io_mat1_1_3),
    .io_mat1_1_4(PreProcessor_io_mat1_1_4),
    .io_mat1_1_5(PreProcessor_io_mat1_1_5),
    .io_mat1_1_6(PreProcessor_io_mat1_1_6),
    .io_mat1_1_7(PreProcessor_io_mat1_1_7),
    .io_mat1_2_0(PreProcessor_io_mat1_2_0),
    .io_mat1_2_1(PreProcessor_io_mat1_2_1),
    .io_mat1_2_2(PreProcessor_io_mat1_2_2),
    .io_mat1_2_3(PreProcessor_io_mat1_2_3),
    .io_mat1_2_4(PreProcessor_io_mat1_2_4),
    .io_mat1_2_5(PreProcessor_io_mat1_2_5),
    .io_mat1_2_6(PreProcessor_io_mat1_2_6),
    .io_mat1_2_7(PreProcessor_io_mat1_2_7),
    .io_mat1_3_0(PreProcessor_io_mat1_3_0),
    .io_mat1_3_1(PreProcessor_io_mat1_3_1),
    .io_mat1_3_2(PreProcessor_io_mat1_3_2),
    .io_mat1_3_3(PreProcessor_io_mat1_3_3),
    .io_mat1_3_4(PreProcessor_io_mat1_3_4),
    .io_mat1_3_5(PreProcessor_io_mat1_3_5),
    .io_mat1_3_6(PreProcessor_io_mat1_3_6),
    .io_mat1_3_7(PreProcessor_io_mat1_3_7),
    .io_mat1_4_0(PreProcessor_io_mat1_4_0),
    .io_mat1_4_1(PreProcessor_io_mat1_4_1),
    .io_mat1_4_2(PreProcessor_io_mat1_4_2),
    .io_mat1_4_3(PreProcessor_io_mat1_4_3),
    .io_mat1_4_4(PreProcessor_io_mat1_4_4),
    .io_mat1_4_5(PreProcessor_io_mat1_4_5),
    .io_mat1_4_6(PreProcessor_io_mat1_4_6),
    .io_mat1_4_7(PreProcessor_io_mat1_4_7),
    .io_mat1_5_0(PreProcessor_io_mat1_5_0),
    .io_mat1_5_1(PreProcessor_io_mat1_5_1),
    .io_mat1_5_2(PreProcessor_io_mat1_5_2),
    .io_mat1_5_3(PreProcessor_io_mat1_5_3),
    .io_mat1_5_4(PreProcessor_io_mat1_5_4),
    .io_mat1_5_5(PreProcessor_io_mat1_5_5),
    .io_mat1_5_6(PreProcessor_io_mat1_5_6),
    .io_mat1_5_7(PreProcessor_io_mat1_5_7),
    .io_mat1_6_0(PreProcessor_io_mat1_6_0),
    .io_mat1_6_1(PreProcessor_io_mat1_6_1),
    .io_mat1_6_2(PreProcessor_io_mat1_6_2),
    .io_mat1_6_3(PreProcessor_io_mat1_6_3),
    .io_mat1_6_4(PreProcessor_io_mat1_6_4),
    .io_mat1_6_5(PreProcessor_io_mat1_6_5),
    .io_mat1_6_6(PreProcessor_io_mat1_6_6),
    .io_mat1_6_7(PreProcessor_io_mat1_6_7),
    .io_mat1_7_0(PreProcessor_io_mat1_7_0),
    .io_mat1_7_1(PreProcessor_io_mat1_7_1),
    .io_mat1_7_2(PreProcessor_io_mat1_7_2),
    .io_mat1_7_3(PreProcessor_io_mat1_7_3),
    .io_mat1_7_4(PreProcessor_io_mat1_7_4),
    .io_mat1_7_5(PreProcessor_io_mat1_7_5),
    .io_mat1_7_6(PreProcessor_io_mat1_7_6),
    .io_mat1_7_7(PreProcessor_io_mat1_7_7),
    .io_mat2_0_0(PreProcessor_io_mat2_0_0),
    .io_mat2_0_1(PreProcessor_io_mat2_0_1),
    .io_mat2_0_2(PreProcessor_io_mat2_0_2),
    .io_mat2_0_3(PreProcessor_io_mat2_0_3),
    .io_mat2_0_4(PreProcessor_io_mat2_0_4),
    .io_mat2_0_5(PreProcessor_io_mat2_0_5),
    .io_mat2_0_6(PreProcessor_io_mat2_0_6),
    .io_mat2_0_7(PreProcessor_io_mat2_0_7),
    .io_mat2_1_0(PreProcessor_io_mat2_1_0),
    .io_mat2_1_1(PreProcessor_io_mat2_1_1),
    .io_mat2_1_2(PreProcessor_io_mat2_1_2),
    .io_mat2_1_3(PreProcessor_io_mat2_1_3),
    .io_mat2_1_4(PreProcessor_io_mat2_1_4),
    .io_mat2_1_5(PreProcessor_io_mat2_1_5),
    .io_mat2_1_6(PreProcessor_io_mat2_1_6),
    .io_mat2_1_7(PreProcessor_io_mat2_1_7),
    .io_mat2_2_0(PreProcessor_io_mat2_2_0),
    .io_mat2_2_1(PreProcessor_io_mat2_2_1),
    .io_mat2_2_2(PreProcessor_io_mat2_2_2),
    .io_mat2_2_3(PreProcessor_io_mat2_2_3),
    .io_mat2_2_4(PreProcessor_io_mat2_2_4),
    .io_mat2_2_5(PreProcessor_io_mat2_2_5),
    .io_mat2_2_6(PreProcessor_io_mat2_2_6),
    .io_mat2_2_7(PreProcessor_io_mat2_2_7),
    .io_mat2_3_0(PreProcessor_io_mat2_3_0),
    .io_mat2_3_1(PreProcessor_io_mat2_3_1),
    .io_mat2_3_2(PreProcessor_io_mat2_3_2),
    .io_mat2_3_3(PreProcessor_io_mat2_3_3),
    .io_mat2_3_4(PreProcessor_io_mat2_3_4),
    .io_mat2_3_5(PreProcessor_io_mat2_3_5),
    .io_mat2_3_6(PreProcessor_io_mat2_3_6),
    .io_mat2_3_7(PreProcessor_io_mat2_3_7),
    .io_mat2_4_0(PreProcessor_io_mat2_4_0),
    .io_mat2_4_1(PreProcessor_io_mat2_4_1),
    .io_mat2_4_2(PreProcessor_io_mat2_4_2),
    .io_mat2_4_3(PreProcessor_io_mat2_4_3),
    .io_mat2_4_4(PreProcessor_io_mat2_4_4),
    .io_mat2_4_5(PreProcessor_io_mat2_4_5),
    .io_mat2_4_6(PreProcessor_io_mat2_4_6),
    .io_mat2_4_7(PreProcessor_io_mat2_4_7),
    .io_mat2_5_0(PreProcessor_io_mat2_5_0),
    .io_mat2_5_1(PreProcessor_io_mat2_5_1),
    .io_mat2_5_2(PreProcessor_io_mat2_5_2),
    .io_mat2_5_3(PreProcessor_io_mat2_5_3),
    .io_mat2_5_4(PreProcessor_io_mat2_5_4),
    .io_mat2_5_5(PreProcessor_io_mat2_5_5),
    .io_mat2_5_6(PreProcessor_io_mat2_5_6),
    .io_mat2_5_7(PreProcessor_io_mat2_5_7),
    .io_mat2_6_0(PreProcessor_io_mat2_6_0),
    .io_mat2_6_1(PreProcessor_io_mat2_6_1),
    .io_mat2_6_2(PreProcessor_io_mat2_6_2),
    .io_mat2_6_3(PreProcessor_io_mat2_6_3),
    .io_mat2_6_4(PreProcessor_io_mat2_6_4),
    .io_mat2_6_5(PreProcessor_io_mat2_6_5),
    .io_mat2_6_6(PreProcessor_io_mat2_6_6),
    .io_mat2_6_7(PreProcessor_io_mat2_6_7),
    .io_mat2_7_0(PreProcessor_io_mat2_7_0),
    .io_mat2_7_1(PreProcessor_io_mat2_7_1),
    .io_mat2_7_2(PreProcessor_io_mat2_7_2),
    .io_mat2_7_3(PreProcessor_io_mat2_7_3),
    .io_mat2_7_4(PreProcessor_io_mat2_7_4),
    .io_mat2_7_5(PreProcessor_io_mat2_7_5),
    .io_mat2_7_6(PreProcessor_io_mat2_7_6),
    .io_mat2_7_7(PreProcessor_io_mat2_7_7),
    .io_compressedBitmap_0_0(PreProcessor_io_compressedBitmap_0_0),
    .io_compressedBitmap_0_1(PreProcessor_io_compressedBitmap_0_1),
    .io_compressedBitmap_0_2(PreProcessor_io_compressedBitmap_0_2),
    .io_compressedBitmap_0_3(PreProcessor_io_compressedBitmap_0_3),
    .io_compressedBitmap_0_4(PreProcessor_io_compressedBitmap_0_4),
    .io_compressedBitmap_0_5(PreProcessor_io_compressedBitmap_0_5),
    .io_compressedBitmap_0_6(PreProcessor_io_compressedBitmap_0_6),
    .io_compressedBitmap_0_7(PreProcessor_io_compressedBitmap_0_7),
    .io_compressedBitmap_1_0(PreProcessor_io_compressedBitmap_1_0),
    .io_compressedBitmap_1_1(PreProcessor_io_compressedBitmap_1_1),
    .io_compressedBitmap_1_2(PreProcessor_io_compressedBitmap_1_2),
    .io_compressedBitmap_1_3(PreProcessor_io_compressedBitmap_1_3),
    .io_compressedBitmap_1_4(PreProcessor_io_compressedBitmap_1_4),
    .io_compressedBitmap_1_5(PreProcessor_io_compressedBitmap_1_5),
    .io_compressedBitmap_1_6(PreProcessor_io_compressedBitmap_1_6),
    .io_compressedBitmap_1_7(PreProcessor_io_compressedBitmap_1_7),
    .io_compressedBitmap_2_0(PreProcessor_io_compressedBitmap_2_0),
    .io_compressedBitmap_2_1(PreProcessor_io_compressedBitmap_2_1),
    .io_compressedBitmap_2_2(PreProcessor_io_compressedBitmap_2_2),
    .io_compressedBitmap_2_3(PreProcessor_io_compressedBitmap_2_3),
    .io_compressedBitmap_2_4(PreProcessor_io_compressedBitmap_2_4),
    .io_compressedBitmap_2_5(PreProcessor_io_compressedBitmap_2_5),
    .io_compressedBitmap_2_6(PreProcessor_io_compressedBitmap_2_6),
    .io_compressedBitmap_2_7(PreProcessor_io_compressedBitmap_2_7),
    .io_compressedBitmap_3_0(PreProcessor_io_compressedBitmap_3_0),
    .io_compressedBitmap_3_1(PreProcessor_io_compressedBitmap_3_1),
    .io_compressedBitmap_3_2(PreProcessor_io_compressedBitmap_3_2),
    .io_compressedBitmap_3_3(PreProcessor_io_compressedBitmap_3_3),
    .io_compressedBitmap_3_4(PreProcessor_io_compressedBitmap_3_4),
    .io_compressedBitmap_3_5(PreProcessor_io_compressedBitmap_3_5),
    .io_compressedBitmap_3_6(PreProcessor_io_compressedBitmap_3_6),
    .io_compressedBitmap_3_7(PreProcessor_io_compressedBitmap_3_7),
    .io_compressedBitmap_4_0(PreProcessor_io_compressedBitmap_4_0),
    .io_compressedBitmap_4_1(PreProcessor_io_compressedBitmap_4_1),
    .io_compressedBitmap_4_2(PreProcessor_io_compressedBitmap_4_2),
    .io_compressedBitmap_4_3(PreProcessor_io_compressedBitmap_4_3),
    .io_compressedBitmap_4_4(PreProcessor_io_compressedBitmap_4_4),
    .io_compressedBitmap_4_5(PreProcessor_io_compressedBitmap_4_5),
    .io_compressedBitmap_4_6(PreProcessor_io_compressedBitmap_4_6),
    .io_compressedBitmap_4_7(PreProcessor_io_compressedBitmap_4_7),
    .io_compressedBitmap_5_0(PreProcessor_io_compressedBitmap_5_0),
    .io_compressedBitmap_5_1(PreProcessor_io_compressedBitmap_5_1),
    .io_compressedBitmap_5_2(PreProcessor_io_compressedBitmap_5_2),
    .io_compressedBitmap_5_3(PreProcessor_io_compressedBitmap_5_3),
    .io_compressedBitmap_5_4(PreProcessor_io_compressedBitmap_5_4),
    .io_compressedBitmap_5_5(PreProcessor_io_compressedBitmap_5_5),
    .io_compressedBitmap_5_6(PreProcessor_io_compressedBitmap_5_6),
    .io_compressedBitmap_5_7(PreProcessor_io_compressedBitmap_5_7),
    .io_compressedBitmap_6_0(PreProcessor_io_compressedBitmap_6_0),
    .io_compressedBitmap_6_1(PreProcessor_io_compressedBitmap_6_1),
    .io_compressedBitmap_6_2(PreProcessor_io_compressedBitmap_6_2),
    .io_compressedBitmap_6_3(PreProcessor_io_compressedBitmap_6_3),
    .io_compressedBitmap_6_4(PreProcessor_io_compressedBitmap_6_4),
    .io_compressedBitmap_6_5(PreProcessor_io_compressedBitmap_6_5),
    .io_compressedBitmap_6_6(PreProcessor_io_compressedBitmap_6_6),
    .io_compressedBitmap_6_7(PreProcessor_io_compressedBitmap_6_7),
    .io_compressedBitmap_7_0(PreProcessor_io_compressedBitmap_7_0),
    .io_compressedBitmap_7_1(PreProcessor_io_compressedBitmap_7_1),
    .io_compressedBitmap_7_2(PreProcessor_io_compressedBitmap_7_2),
    .io_compressedBitmap_7_3(PreProcessor_io_compressedBitmap_7_3),
    .io_compressedBitmap_7_4(PreProcessor_io_compressedBitmap_7_4),
    .io_compressedBitmap_7_5(PreProcessor_io_compressedBitmap_7_5),
    .io_compressedBitmap_7_6(PreProcessor_io_compressedBitmap_7_6),
    .io_compressedBitmap_7_7(PreProcessor_io_compressedBitmap_7_7)
  );
  FlexDPU FDPU ( // @[TOP.scala 25:26]
    .clock(FDPU_clock),
    .reset(FDPU_reset),
    .io_Stationary_matrix_0_0(FDPU_io_Stationary_matrix_0_0),
    .io_Stationary_matrix_0_1(FDPU_io_Stationary_matrix_0_1),
    .io_Stationary_matrix_0_2(FDPU_io_Stationary_matrix_0_2),
    .io_Stationary_matrix_0_3(FDPU_io_Stationary_matrix_0_3),
    .io_Stationary_matrix_0_4(FDPU_io_Stationary_matrix_0_4),
    .io_Stationary_matrix_0_5(FDPU_io_Stationary_matrix_0_5),
    .io_Stationary_matrix_0_6(FDPU_io_Stationary_matrix_0_6),
    .io_Stationary_matrix_0_7(FDPU_io_Stationary_matrix_0_7),
    .io_Stationary_matrix_1_0(FDPU_io_Stationary_matrix_1_0),
    .io_Stationary_matrix_1_1(FDPU_io_Stationary_matrix_1_1),
    .io_Stationary_matrix_1_2(FDPU_io_Stationary_matrix_1_2),
    .io_Stationary_matrix_1_3(FDPU_io_Stationary_matrix_1_3),
    .io_Stationary_matrix_1_4(FDPU_io_Stationary_matrix_1_4),
    .io_Stationary_matrix_1_5(FDPU_io_Stationary_matrix_1_5),
    .io_Stationary_matrix_1_6(FDPU_io_Stationary_matrix_1_6),
    .io_Stationary_matrix_1_7(FDPU_io_Stationary_matrix_1_7),
    .io_Stationary_matrix_2_0(FDPU_io_Stationary_matrix_2_0),
    .io_Stationary_matrix_2_1(FDPU_io_Stationary_matrix_2_1),
    .io_Stationary_matrix_2_2(FDPU_io_Stationary_matrix_2_2),
    .io_Stationary_matrix_2_3(FDPU_io_Stationary_matrix_2_3),
    .io_Stationary_matrix_2_4(FDPU_io_Stationary_matrix_2_4),
    .io_Stationary_matrix_2_5(FDPU_io_Stationary_matrix_2_5),
    .io_Stationary_matrix_2_6(FDPU_io_Stationary_matrix_2_6),
    .io_Stationary_matrix_2_7(FDPU_io_Stationary_matrix_2_7),
    .io_Stationary_matrix_3_0(FDPU_io_Stationary_matrix_3_0),
    .io_Stationary_matrix_3_1(FDPU_io_Stationary_matrix_3_1),
    .io_Stationary_matrix_3_2(FDPU_io_Stationary_matrix_3_2),
    .io_Stationary_matrix_3_3(FDPU_io_Stationary_matrix_3_3),
    .io_Stationary_matrix_3_4(FDPU_io_Stationary_matrix_3_4),
    .io_Stationary_matrix_3_5(FDPU_io_Stationary_matrix_3_5),
    .io_Stationary_matrix_3_6(FDPU_io_Stationary_matrix_3_6),
    .io_Stationary_matrix_3_7(FDPU_io_Stationary_matrix_3_7),
    .io_Stationary_matrix_4_0(FDPU_io_Stationary_matrix_4_0),
    .io_Stationary_matrix_4_1(FDPU_io_Stationary_matrix_4_1),
    .io_Stationary_matrix_4_2(FDPU_io_Stationary_matrix_4_2),
    .io_Stationary_matrix_4_3(FDPU_io_Stationary_matrix_4_3),
    .io_Stationary_matrix_4_4(FDPU_io_Stationary_matrix_4_4),
    .io_Stationary_matrix_4_5(FDPU_io_Stationary_matrix_4_5),
    .io_Stationary_matrix_4_6(FDPU_io_Stationary_matrix_4_6),
    .io_Stationary_matrix_4_7(FDPU_io_Stationary_matrix_4_7),
    .io_Stationary_matrix_5_0(FDPU_io_Stationary_matrix_5_0),
    .io_Stationary_matrix_5_1(FDPU_io_Stationary_matrix_5_1),
    .io_Stationary_matrix_5_2(FDPU_io_Stationary_matrix_5_2),
    .io_Stationary_matrix_5_3(FDPU_io_Stationary_matrix_5_3),
    .io_Stationary_matrix_5_4(FDPU_io_Stationary_matrix_5_4),
    .io_Stationary_matrix_5_5(FDPU_io_Stationary_matrix_5_5),
    .io_Stationary_matrix_5_6(FDPU_io_Stationary_matrix_5_6),
    .io_Stationary_matrix_5_7(FDPU_io_Stationary_matrix_5_7),
    .io_Stationary_matrix_6_0(FDPU_io_Stationary_matrix_6_0),
    .io_Stationary_matrix_6_1(FDPU_io_Stationary_matrix_6_1),
    .io_Stationary_matrix_6_2(FDPU_io_Stationary_matrix_6_2),
    .io_Stationary_matrix_6_3(FDPU_io_Stationary_matrix_6_3),
    .io_Stationary_matrix_6_4(FDPU_io_Stationary_matrix_6_4),
    .io_Stationary_matrix_6_5(FDPU_io_Stationary_matrix_6_5),
    .io_Stationary_matrix_6_6(FDPU_io_Stationary_matrix_6_6),
    .io_Stationary_matrix_6_7(FDPU_io_Stationary_matrix_6_7),
    .io_Stationary_matrix_7_0(FDPU_io_Stationary_matrix_7_0),
    .io_Stationary_matrix_7_1(FDPU_io_Stationary_matrix_7_1),
    .io_Stationary_matrix_7_2(FDPU_io_Stationary_matrix_7_2),
    .io_Stationary_matrix_7_3(FDPU_io_Stationary_matrix_7_3),
    .io_Stationary_matrix_7_4(FDPU_io_Stationary_matrix_7_4),
    .io_Stationary_matrix_7_5(FDPU_io_Stationary_matrix_7_5),
    .io_Stationary_matrix_7_6(FDPU_io_Stationary_matrix_7_6),
    .io_Stationary_matrix_7_7(FDPU_io_Stationary_matrix_7_7),
    .io_Streaming_matrix_0_0(FDPU_io_Streaming_matrix_0_0),
    .io_Streaming_matrix_0_1(FDPU_io_Streaming_matrix_0_1),
    .io_Streaming_matrix_0_2(FDPU_io_Streaming_matrix_0_2),
    .io_Streaming_matrix_0_3(FDPU_io_Streaming_matrix_0_3),
    .io_Streaming_matrix_0_4(FDPU_io_Streaming_matrix_0_4),
    .io_Streaming_matrix_0_5(FDPU_io_Streaming_matrix_0_5),
    .io_Streaming_matrix_0_6(FDPU_io_Streaming_matrix_0_6),
    .io_Streaming_matrix_0_7(FDPU_io_Streaming_matrix_0_7),
    .io_Streaming_matrix_1_0(FDPU_io_Streaming_matrix_1_0),
    .io_Streaming_matrix_1_1(FDPU_io_Streaming_matrix_1_1),
    .io_Streaming_matrix_1_2(FDPU_io_Streaming_matrix_1_2),
    .io_Streaming_matrix_1_3(FDPU_io_Streaming_matrix_1_3),
    .io_Streaming_matrix_1_4(FDPU_io_Streaming_matrix_1_4),
    .io_Streaming_matrix_1_5(FDPU_io_Streaming_matrix_1_5),
    .io_Streaming_matrix_1_6(FDPU_io_Streaming_matrix_1_6),
    .io_Streaming_matrix_1_7(FDPU_io_Streaming_matrix_1_7),
    .io_Streaming_matrix_2_0(FDPU_io_Streaming_matrix_2_0),
    .io_Streaming_matrix_2_1(FDPU_io_Streaming_matrix_2_1),
    .io_Streaming_matrix_2_2(FDPU_io_Streaming_matrix_2_2),
    .io_Streaming_matrix_2_3(FDPU_io_Streaming_matrix_2_3),
    .io_Streaming_matrix_2_4(FDPU_io_Streaming_matrix_2_4),
    .io_Streaming_matrix_2_5(FDPU_io_Streaming_matrix_2_5),
    .io_Streaming_matrix_2_6(FDPU_io_Streaming_matrix_2_6),
    .io_Streaming_matrix_2_7(FDPU_io_Streaming_matrix_2_7),
    .io_Streaming_matrix_3_0(FDPU_io_Streaming_matrix_3_0),
    .io_Streaming_matrix_3_1(FDPU_io_Streaming_matrix_3_1),
    .io_Streaming_matrix_3_2(FDPU_io_Streaming_matrix_3_2),
    .io_Streaming_matrix_3_3(FDPU_io_Streaming_matrix_3_3),
    .io_Streaming_matrix_3_4(FDPU_io_Streaming_matrix_3_4),
    .io_Streaming_matrix_3_5(FDPU_io_Streaming_matrix_3_5),
    .io_Streaming_matrix_3_6(FDPU_io_Streaming_matrix_3_6),
    .io_Streaming_matrix_3_7(FDPU_io_Streaming_matrix_3_7),
    .io_Streaming_matrix_4_0(FDPU_io_Streaming_matrix_4_0),
    .io_Streaming_matrix_4_1(FDPU_io_Streaming_matrix_4_1),
    .io_Streaming_matrix_4_2(FDPU_io_Streaming_matrix_4_2),
    .io_Streaming_matrix_4_3(FDPU_io_Streaming_matrix_4_3),
    .io_Streaming_matrix_4_4(FDPU_io_Streaming_matrix_4_4),
    .io_Streaming_matrix_4_5(FDPU_io_Streaming_matrix_4_5),
    .io_Streaming_matrix_4_6(FDPU_io_Streaming_matrix_4_6),
    .io_Streaming_matrix_4_7(FDPU_io_Streaming_matrix_4_7),
    .io_Streaming_matrix_5_0(FDPU_io_Streaming_matrix_5_0),
    .io_Streaming_matrix_5_1(FDPU_io_Streaming_matrix_5_1),
    .io_Streaming_matrix_5_2(FDPU_io_Streaming_matrix_5_2),
    .io_Streaming_matrix_5_3(FDPU_io_Streaming_matrix_5_3),
    .io_Streaming_matrix_5_4(FDPU_io_Streaming_matrix_5_4),
    .io_Streaming_matrix_5_5(FDPU_io_Streaming_matrix_5_5),
    .io_Streaming_matrix_5_6(FDPU_io_Streaming_matrix_5_6),
    .io_Streaming_matrix_5_7(FDPU_io_Streaming_matrix_5_7),
    .io_Streaming_matrix_6_0(FDPU_io_Streaming_matrix_6_0),
    .io_Streaming_matrix_6_1(FDPU_io_Streaming_matrix_6_1),
    .io_Streaming_matrix_6_2(FDPU_io_Streaming_matrix_6_2),
    .io_Streaming_matrix_6_3(FDPU_io_Streaming_matrix_6_3),
    .io_Streaming_matrix_6_4(FDPU_io_Streaming_matrix_6_4),
    .io_Streaming_matrix_6_5(FDPU_io_Streaming_matrix_6_5),
    .io_Streaming_matrix_6_6(FDPU_io_Streaming_matrix_6_6),
    .io_Streaming_matrix_6_7(FDPU_io_Streaming_matrix_6_7),
    .io_Streaming_matrix_7_0(FDPU_io_Streaming_matrix_7_0),
    .io_Streaming_matrix_7_1(FDPU_io_Streaming_matrix_7_1),
    .io_Streaming_matrix_7_2(FDPU_io_Streaming_matrix_7_2),
    .io_Streaming_matrix_7_3(FDPU_io_Streaming_matrix_7_3),
    .io_Streaming_matrix_7_4(FDPU_io_Streaming_matrix_7_4),
    .io_Streaming_matrix_7_5(FDPU_io_Streaming_matrix_7_5),
    .io_Streaming_matrix_7_6(FDPU_io_Streaming_matrix_7_6),
    .io_Streaming_matrix_7_7(FDPU_io_Streaming_matrix_7_7)
  );
  assign io_Third_Matrix_0_0 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_0_1 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_0_2 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_0_3 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_0_4 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_0_5 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_0_6 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_0_7 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_1_0 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_1_1 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_1_2 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_1_3 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_1_4 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_1_5 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_1_6 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_1_7 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_2_0 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_2_1 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_2_2 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_2_3 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_2_4 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_2_5 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_2_6 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_2_7 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_3_0 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_3_1 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_3_2 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_3_3 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_3_4 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_3_5 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_3_6 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_3_7 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_4_0 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_4_1 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_4_2 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_4_3 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_4_4 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_4_5 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_4_6 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_4_7 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_5_0 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_5_1 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_5_2 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_5_3 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_5_4 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_5_5 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_5_6 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_5_7 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_6_0 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_6_1 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_6_2 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_6_3 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_6_4 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_6_5 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_6_6 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_6_7 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_7_0 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_7_1 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_7_2 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_7_3 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_7_4 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_7_5 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_7_6 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign io_Third_Matrix_7_7 = 32'h0; // @[TOP.scala 24:25 31:25 33:25]
  assign PreProcessor_clock = clock;
  assign PreProcessor_reset = reset;
  assign PreProcessor_io_mat1_0_0 = io_Stationary_matrix_0_0[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_0_1 = io_Stationary_matrix_0_1[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_0_2 = io_Stationary_matrix_0_2[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_0_3 = io_Stationary_matrix_0_3[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_0_4 = io_Stationary_matrix_0_4[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_0_5 = io_Stationary_matrix_0_5[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_0_6 = io_Stationary_matrix_0_6[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_0_7 = io_Stationary_matrix_0_7[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_1_0 = io_Stationary_matrix_1_0[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_1_1 = io_Stationary_matrix_1_1[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_1_2 = io_Stationary_matrix_1_2[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_1_3 = io_Stationary_matrix_1_3[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_1_4 = io_Stationary_matrix_1_4[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_1_5 = io_Stationary_matrix_1_5[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_1_6 = io_Stationary_matrix_1_6[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_1_7 = io_Stationary_matrix_1_7[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_2_0 = io_Stationary_matrix_2_0[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_2_1 = io_Stationary_matrix_2_1[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_2_2 = io_Stationary_matrix_2_2[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_2_3 = io_Stationary_matrix_2_3[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_2_4 = io_Stationary_matrix_2_4[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_2_5 = io_Stationary_matrix_2_5[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_2_6 = io_Stationary_matrix_2_6[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_2_7 = io_Stationary_matrix_2_7[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_3_0 = io_Stationary_matrix_3_0[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_3_1 = io_Stationary_matrix_3_1[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_3_2 = io_Stationary_matrix_3_2[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_3_3 = io_Stationary_matrix_3_3[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_3_4 = io_Stationary_matrix_3_4[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_3_5 = io_Stationary_matrix_3_5[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_3_6 = io_Stationary_matrix_3_6[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_3_7 = io_Stationary_matrix_3_7[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_4_0 = io_Stationary_matrix_4_0[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_4_1 = io_Stationary_matrix_4_1[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_4_2 = io_Stationary_matrix_4_2[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_4_3 = io_Stationary_matrix_4_3[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_4_4 = io_Stationary_matrix_4_4[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_4_5 = io_Stationary_matrix_4_5[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_4_6 = io_Stationary_matrix_4_6[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_4_7 = io_Stationary_matrix_4_7[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_5_0 = io_Stationary_matrix_5_0[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_5_1 = io_Stationary_matrix_5_1[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_5_2 = io_Stationary_matrix_5_2[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_5_3 = io_Stationary_matrix_5_3[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_5_4 = io_Stationary_matrix_5_4[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_5_5 = io_Stationary_matrix_5_5[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_5_6 = io_Stationary_matrix_5_6[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_5_7 = io_Stationary_matrix_5_7[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_6_0 = io_Stationary_matrix_6_0[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_6_1 = io_Stationary_matrix_6_1[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_6_2 = io_Stationary_matrix_6_2[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_6_3 = io_Stationary_matrix_6_3[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_6_4 = io_Stationary_matrix_6_4[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_6_5 = io_Stationary_matrix_6_5[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_6_6 = io_Stationary_matrix_6_6[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_6_7 = io_Stationary_matrix_6_7[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_7_0 = io_Stationary_matrix_7_0[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_7_1 = io_Stationary_matrix_7_1[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_7_2 = io_Stationary_matrix_7_2[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_7_3 = io_Stationary_matrix_7_3[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_7_4 = io_Stationary_matrix_7_4[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_7_5 = io_Stationary_matrix_7_5[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_7_6 = io_Stationary_matrix_7_6[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat1_7_7 = io_Stationary_matrix_7_7[15:0]; // @[TOP.scala 15:26]
  assign PreProcessor_io_mat2_0_0 = io_Streaming_matrix_0_0[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_0_1 = io_Streaming_matrix_0_1[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_0_2 = io_Streaming_matrix_0_2[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_0_3 = io_Streaming_matrix_0_3[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_0_4 = io_Streaming_matrix_0_4[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_0_5 = io_Streaming_matrix_0_5[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_0_6 = io_Streaming_matrix_0_6[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_0_7 = io_Streaming_matrix_0_7[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_1_0 = io_Streaming_matrix_1_0[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_1_1 = io_Streaming_matrix_1_1[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_1_2 = io_Streaming_matrix_1_2[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_1_3 = io_Streaming_matrix_1_3[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_1_4 = io_Streaming_matrix_1_4[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_1_5 = io_Streaming_matrix_1_5[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_1_6 = io_Streaming_matrix_1_6[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_1_7 = io_Streaming_matrix_1_7[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_2_0 = io_Streaming_matrix_2_0[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_2_1 = io_Streaming_matrix_2_1[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_2_2 = io_Streaming_matrix_2_2[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_2_3 = io_Streaming_matrix_2_3[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_2_4 = io_Streaming_matrix_2_4[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_2_5 = io_Streaming_matrix_2_5[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_2_6 = io_Streaming_matrix_2_6[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_2_7 = io_Streaming_matrix_2_7[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_3_0 = io_Streaming_matrix_3_0[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_3_1 = io_Streaming_matrix_3_1[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_3_2 = io_Streaming_matrix_3_2[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_3_3 = io_Streaming_matrix_3_3[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_3_4 = io_Streaming_matrix_3_4[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_3_5 = io_Streaming_matrix_3_5[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_3_6 = io_Streaming_matrix_3_6[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_3_7 = io_Streaming_matrix_3_7[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_4_0 = io_Streaming_matrix_4_0[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_4_1 = io_Streaming_matrix_4_1[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_4_2 = io_Streaming_matrix_4_2[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_4_3 = io_Streaming_matrix_4_3[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_4_4 = io_Streaming_matrix_4_4[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_4_5 = io_Streaming_matrix_4_5[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_4_6 = io_Streaming_matrix_4_6[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_4_7 = io_Streaming_matrix_4_7[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_5_0 = io_Streaming_matrix_5_0[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_5_1 = io_Streaming_matrix_5_1[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_5_2 = io_Streaming_matrix_5_2[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_5_3 = io_Streaming_matrix_5_3[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_5_4 = io_Streaming_matrix_5_4[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_5_5 = io_Streaming_matrix_5_5[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_5_6 = io_Streaming_matrix_5_6[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_5_7 = io_Streaming_matrix_5_7[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_6_0 = io_Streaming_matrix_6_0[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_6_1 = io_Streaming_matrix_6_1[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_6_2 = io_Streaming_matrix_6_2[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_6_3 = io_Streaming_matrix_6_3[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_6_4 = io_Streaming_matrix_6_4[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_6_5 = io_Streaming_matrix_6_5[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_6_6 = io_Streaming_matrix_6_6[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_6_7 = io_Streaming_matrix_6_7[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_7_0 = io_Streaming_matrix_7_0[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_7_1 = io_Streaming_matrix_7_1[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_7_2 = io_Streaming_matrix_7_2[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_7_3 = io_Streaming_matrix_7_3[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_7_4 = io_Streaming_matrix_7_4[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_7_5 = io_Streaming_matrix_7_5[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_7_6 = io_Streaming_matrix_7_6[15:0]; // @[TOP.scala 16:26]
  assign PreProcessor_io_mat2_7_7 = io_Streaming_matrix_7_7[15:0]; // @[TOP.scala 16:26]
  assign FDPU_clock = clock;
  assign FDPU_reset = reset;
  assign FDPU_io_Stationary_matrix_0_0 = PreProcessor_io_compressedBitmap_0_0; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_0_1 = PreProcessor_io_compressedBitmap_0_1; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_0_2 = PreProcessor_io_compressedBitmap_0_2; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_0_3 = PreProcessor_io_compressedBitmap_0_3; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_0_4 = PreProcessor_io_compressedBitmap_0_4; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_0_5 = PreProcessor_io_compressedBitmap_0_5; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_0_6 = PreProcessor_io_compressedBitmap_0_6; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_0_7 = PreProcessor_io_compressedBitmap_0_7; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_1_0 = PreProcessor_io_compressedBitmap_1_0; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_1_1 = PreProcessor_io_compressedBitmap_1_1; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_1_2 = PreProcessor_io_compressedBitmap_1_2; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_1_3 = PreProcessor_io_compressedBitmap_1_3; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_1_4 = PreProcessor_io_compressedBitmap_1_4; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_1_5 = PreProcessor_io_compressedBitmap_1_5; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_1_6 = PreProcessor_io_compressedBitmap_1_6; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_1_7 = PreProcessor_io_compressedBitmap_1_7; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_2_0 = PreProcessor_io_compressedBitmap_2_0; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_2_1 = PreProcessor_io_compressedBitmap_2_1; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_2_2 = PreProcessor_io_compressedBitmap_2_2; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_2_3 = PreProcessor_io_compressedBitmap_2_3; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_2_4 = PreProcessor_io_compressedBitmap_2_4; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_2_5 = PreProcessor_io_compressedBitmap_2_5; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_2_6 = PreProcessor_io_compressedBitmap_2_6; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_2_7 = PreProcessor_io_compressedBitmap_2_7; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_3_0 = PreProcessor_io_compressedBitmap_3_0; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_3_1 = PreProcessor_io_compressedBitmap_3_1; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_3_2 = PreProcessor_io_compressedBitmap_3_2; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_3_3 = PreProcessor_io_compressedBitmap_3_3; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_3_4 = PreProcessor_io_compressedBitmap_3_4; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_3_5 = PreProcessor_io_compressedBitmap_3_5; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_3_6 = PreProcessor_io_compressedBitmap_3_6; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_3_7 = PreProcessor_io_compressedBitmap_3_7; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_4_0 = PreProcessor_io_compressedBitmap_4_0; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_4_1 = PreProcessor_io_compressedBitmap_4_1; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_4_2 = PreProcessor_io_compressedBitmap_4_2; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_4_3 = PreProcessor_io_compressedBitmap_4_3; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_4_4 = PreProcessor_io_compressedBitmap_4_4; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_4_5 = PreProcessor_io_compressedBitmap_4_5; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_4_6 = PreProcessor_io_compressedBitmap_4_6; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_4_7 = PreProcessor_io_compressedBitmap_4_7; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_5_0 = PreProcessor_io_compressedBitmap_5_0; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_5_1 = PreProcessor_io_compressedBitmap_5_1; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_5_2 = PreProcessor_io_compressedBitmap_5_2; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_5_3 = PreProcessor_io_compressedBitmap_5_3; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_5_4 = PreProcessor_io_compressedBitmap_5_4; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_5_5 = PreProcessor_io_compressedBitmap_5_5; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_5_6 = PreProcessor_io_compressedBitmap_5_6; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_5_7 = PreProcessor_io_compressedBitmap_5_7; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_6_0 = PreProcessor_io_compressedBitmap_6_0; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_6_1 = PreProcessor_io_compressedBitmap_6_1; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_6_2 = PreProcessor_io_compressedBitmap_6_2; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_6_3 = PreProcessor_io_compressedBitmap_6_3; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_6_4 = PreProcessor_io_compressedBitmap_6_4; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_6_5 = PreProcessor_io_compressedBitmap_6_5; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_6_6 = PreProcessor_io_compressedBitmap_6_6; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_6_7 = PreProcessor_io_compressedBitmap_6_7; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_7_0 = PreProcessor_io_compressedBitmap_7_0; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_7_1 = PreProcessor_io_compressedBitmap_7_1; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_7_2 = PreProcessor_io_compressedBitmap_7_2; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_7_3 = PreProcessor_io_compressedBitmap_7_3; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_7_4 = PreProcessor_io_compressedBitmap_7_4; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_7_5 = PreProcessor_io_compressedBitmap_7_5; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_7_6 = PreProcessor_io_compressedBitmap_7_6; // @[TOP.scala 28:35]
  assign FDPU_io_Stationary_matrix_7_7 = PreProcessor_io_compressedBitmap_7_7; // @[TOP.scala 28:35]
  assign FDPU_io_Streaming_matrix_0_0 = io_Streaming_matrix_0_0[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_0_1 = io_Streaming_matrix_0_1[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_0_2 = io_Streaming_matrix_0_2[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_0_3 = io_Streaming_matrix_0_3[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_0_4 = io_Streaming_matrix_0_4[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_0_5 = io_Streaming_matrix_0_5[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_0_6 = io_Streaming_matrix_0_6[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_0_7 = io_Streaming_matrix_0_7[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_1_0 = io_Streaming_matrix_1_0[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_1_1 = io_Streaming_matrix_1_1[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_1_2 = io_Streaming_matrix_1_2[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_1_3 = io_Streaming_matrix_1_3[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_1_4 = io_Streaming_matrix_1_4[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_1_5 = io_Streaming_matrix_1_5[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_1_6 = io_Streaming_matrix_1_6[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_1_7 = io_Streaming_matrix_1_7[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_2_0 = io_Streaming_matrix_2_0[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_2_1 = io_Streaming_matrix_2_1[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_2_2 = io_Streaming_matrix_2_2[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_2_3 = io_Streaming_matrix_2_3[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_2_4 = io_Streaming_matrix_2_4[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_2_5 = io_Streaming_matrix_2_5[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_2_6 = io_Streaming_matrix_2_6[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_2_7 = io_Streaming_matrix_2_7[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_3_0 = io_Streaming_matrix_3_0[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_3_1 = io_Streaming_matrix_3_1[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_3_2 = io_Streaming_matrix_3_2[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_3_3 = io_Streaming_matrix_3_3[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_3_4 = io_Streaming_matrix_3_4[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_3_5 = io_Streaming_matrix_3_5[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_3_6 = io_Streaming_matrix_3_6[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_3_7 = io_Streaming_matrix_3_7[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_4_0 = io_Streaming_matrix_4_0[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_4_1 = io_Streaming_matrix_4_1[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_4_2 = io_Streaming_matrix_4_2[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_4_3 = io_Streaming_matrix_4_3[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_4_4 = io_Streaming_matrix_4_4[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_4_5 = io_Streaming_matrix_4_5[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_4_6 = io_Streaming_matrix_4_6[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_4_7 = io_Streaming_matrix_4_7[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_5_0 = io_Streaming_matrix_5_0[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_5_1 = io_Streaming_matrix_5_1[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_5_2 = io_Streaming_matrix_5_2[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_5_3 = io_Streaming_matrix_5_3[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_5_4 = io_Streaming_matrix_5_4[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_5_5 = io_Streaming_matrix_5_5[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_5_6 = io_Streaming_matrix_5_6[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_5_7 = io_Streaming_matrix_5_7[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_6_0 = io_Streaming_matrix_6_0[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_6_1 = io_Streaming_matrix_6_1[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_6_2 = io_Streaming_matrix_6_2[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_6_3 = io_Streaming_matrix_6_3[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_6_4 = io_Streaming_matrix_6_4[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_6_5 = io_Streaming_matrix_6_5[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_6_6 = io_Streaming_matrix_6_6[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_6_7 = io_Streaming_matrix_6_7[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_7_0 = io_Streaming_matrix_7_0[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_7_1 = io_Streaming_matrix_7_1[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_7_2 = io_Streaming_matrix_7_2[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_7_3 = io_Streaming_matrix_7_3[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_7_4 = io_Streaming_matrix_7_4[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_7_5 = io_Streaming_matrix_7_5[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_7_6 = io_Streaming_matrix_7_6[15:0]; // @[TOP.scala 29:34]
  assign FDPU_io_Streaming_matrix_7_7 = io_Streaming_matrix_7_7[15:0]; // @[TOP.scala 29:34]
endmodule
