module InputSwitch(
  output [31:0] io_y,
  output [31:0] io_z,
  input  [31:0] io_in
);
  assign io_y = io_in; // @[Switches.scala 13:8]
  assign io_z = io_in; // @[Switches.scala 14:8]
endmodule
module BenesMux(
  output [31:0] io_o,
  input  [31:0] io_a,
  input  [31:0] io_b,
  input         io_sel
);
  assign io_o = io_sel ? io_b : io_a; // @[Switches.scala 65:14]
endmodule
module OutputSwitch(
  output [31:0] io_y,
  input  [31:0] io_in0,
  input  [31:0] io_in1,
  input         io_sel
);
  wire [31:0] mux0_io_o; // @[Switches.scala 26:20]
  wire [31:0] mux0_io_a; // @[Switches.scala 26:20]
  wire [31:0] mux0_io_b; // @[Switches.scala 26:20]
  wire  mux0_io_sel; // @[Switches.scala 26:20]
  BenesMux mux0 ( // @[Switches.scala 26:20]
    .io_o(mux0_io_o),
    .io_a(mux0_io_a),
    .io_b(mux0_io_b),
    .io_sel(mux0_io_sel)
  );
  assign io_y = mux0_io_o; // @[Switches.scala 30:8]
  assign mux0_io_a = io_in0; // @[Switches.scala 27:13]
  assign mux0_io_b = io_in1; // @[Switches.scala 28:13]
  assign mux0_io_sel = io_sel; // @[Switches.scala 29:15]
endmodule
module Switch(
  output [31:0] io_y,
  output [31:0] io_z,
  input  [31:0] io_in0,
  input  [31:0] io_in1,
  input         io_sel0,
  input         io_sel1
);
  wire [31:0] mux0_io_o; // @[Switches.scala 44:20]
  wire [31:0] mux0_io_a; // @[Switches.scala 44:20]
  wire [31:0] mux0_io_b; // @[Switches.scala 44:20]
  wire  mux0_io_sel; // @[Switches.scala 44:20]
  wire [31:0] mux1_io_o; // @[Switches.scala 45:20]
  wire [31:0] mux1_io_a; // @[Switches.scala 45:20]
  wire [31:0] mux1_io_b; // @[Switches.scala 45:20]
  wire  mux1_io_sel; // @[Switches.scala 45:20]
  BenesMux mux0 ( // @[Switches.scala 44:20]
    .io_o(mux0_io_o),
    .io_a(mux0_io_a),
    .io_b(mux0_io_b),
    .io_sel(mux0_io_sel)
  );
  BenesMux mux1 ( // @[Switches.scala 45:20]
    .io_o(mux1_io_o),
    .io_a(mux1_io_a),
    .io_b(mux1_io_b),
    .io_sel(mux1_io_sel)
  );
  assign io_y = mux0_io_o; // @[Switches.scala 52:8]
  assign io_z = mux1_io_o; // @[Switches.scala 53:8]
  assign mux0_io_a = io_in0; // @[Switches.scala 46:13]
  assign mux0_io_b = io_in1; // @[Switches.scala 47:13]
  assign mux0_io_sel = io_sel0; // @[Switches.scala 48:15]
  assign mux1_io_a = io_in0; // @[Switches.scala 49:13]
  assign mux1_io_b = io_in1; // @[Switches.scala 50:13]
  assign mux1_io_sel = io_sel1; // @[Switches.scala 51:15]
endmodule
module Benes(
  input         clock,
  input         reset,
  input  [31:0] io_i_data_bus_0,
  input  [31:0] io_i_data_bus_1,
  input  [31:0] io_i_data_bus_2,
  input  [31:0] io_i_data_bus_3,
  input  [31:0] io_i_data_bus_4,
  input  [31:0] io_i_data_bus_5,
  input  [31:0] io_i_data_bus_6,
  input  [31:0] io_i_data_bus_7,
  input  [31:0] io_i_data_bus_8,
  input  [31:0] io_i_data_bus_9,
  input  [31:0] io_i_data_bus_10,
  input  [31:0] io_i_data_bus_11,
  input  [31:0] io_i_data_bus_12,
  input  [31:0] io_i_data_bus_13,
  input  [31:0] io_i_data_bus_14,
  input  [31:0] io_i_data_bus_15,
  input  [31:0] io_i_data_bus_16,
  input  [31:0] io_i_data_bus_17,
  input  [31:0] io_i_data_bus_18,
  input  [31:0] io_i_data_bus_19,
  input  [31:0] io_i_data_bus_20,
  input  [31:0] io_i_data_bus_21,
  input  [31:0] io_i_data_bus_22,
  input  [31:0] io_i_data_bus_23,
  input  [31:0] io_i_data_bus_24,
  input  [31:0] io_i_data_bus_25,
  input  [31:0] io_i_data_bus_26,
  input  [31:0] io_i_data_bus_27,
  input  [31:0] io_i_data_bus_28,
  input  [31:0] io_i_data_bus_29,
  input  [31:0] io_i_data_bus_30,
  input  [31:0] io_i_data_bus_31,
  input         io_i_mux_bus_0,
  input         io_i_mux_bus_1,
  input         io_i_mux_bus_2,
  input         io_i_mux_bus_3,
  input         io_i_mux_bus_4,
  input         io_i_mux_bus_5,
  input         io_i_mux_bus_6,
  input         io_i_mux_bus_7,
  input         io_i_mux_bus_8,
  input         io_i_mux_bus_9,
  input         io_i_mux_bus_10,
  input         io_i_mux_bus_11,
  input         io_i_mux_bus_12,
  input         io_i_mux_bus_13,
  input         io_i_mux_bus_14,
  input         io_i_mux_bus_15,
  input         io_i_mux_bus_16,
  input         io_i_mux_bus_17,
  input         io_i_mux_bus_18,
  input         io_i_mux_bus_19,
  input         io_i_mux_bus_20,
  input         io_i_mux_bus_21,
  input         io_i_mux_bus_22,
  input         io_i_mux_bus_23,
  input         io_i_mux_bus_24,
  input         io_i_mux_bus_25,
  input         io_i_mux_bus_26,
  input         io_i_mux_bus_27,
  input         io_i_mux_bus_28,
  input         io_i_mux_bus_29,
  input         io_i_mux_bus_30,
  input         io_i_mux_bus_31,
  input         io_i_mux_bus_32,
  input         io_i_mux_bus_33,
  input         io_i_mux_bus_34,
  input         io_i_mux_bus_35,
  input         io_i_mux_bus_36,
  input         io_i_mux_bus_37,
  input         io_i_mux_bus_38,
  input         io_i_mux_bus_39,
  input         io_i_mux_bus_40,
  input         io_i_mux_bus_41,
  input         io_i_mux_bus_42,
  input         io_i_mux_bus_43,
  input         io_i_mux_bus_44,
  input         io_i_mux_bus_45,
  input         io_i_mux_bus_46,
  input         io_i_mux_bus_47,
  input         io_i_mux_bus_48,
  input         io_i_mux_bus_49,
  input         io_i_mux_bus_50,
  input         io_i_mux_bus_51,
  input         io_i_mux_bus_52,
  input         io_i_mux_bus_53,
  input         io_i_mux_bus_54,
  input         io_i_mux_bus_55,
  input         io_i_mux_bus_56,
  input         io_i_mux_bus_57,
  input         io_i_mux_bus_58,
  input         io_i_mux_bus_59,
  input         io_i_mux_bus_60,
  input         io_i_mux_bus_61,
  input         io_i_mux_bus_62,
  input         io_i_mux_bus_63,
  input         io_i_mux_bus_64,
  input         io_i_mux_bus_65,
  input         io_i_mux_bus_66,
  input         io_i_mux_bus_67,
  input         io_i_mux_bus_68,
  input         io_i_mux_bus_69,
  input         io_i_mux_bus_70,
  input         io_i_mux_bus_71,
  input         io_i_mux_bus_72,
  input         io_i_mux_bus_73,
  input         io_i_mux_bus_74,
  input         io_i_mux_bus_75,
  input         io_i_mux_bus_76,
  input         io_i_mux_bus_77,
  input         io_i_mux_bus_78,
  input         io_i_mux_bus_79,
  input         io_i_mux_bus_80,
  input         io_i_mux_bus_81,
  input         io_i_mux_bus_82,
  input         io_i_mux_bus_83,
  input         io_i_mux_bus_84,
  input         io_i_mux_bus_85,
  input         io_i_mux_bus_86,
  input         io_i_mux_bus_87,
  input         io_i_mux_bus_88,
  input         io_i_mux_bus_89,
  input         io_i_mux_bus_90,
  input         io_i_mux_bus_91,
  input         io_i_mux_bus_92,
  input         io_i_mux_bus_93,
  input         io_i_mux_bus_94,
  input         io_i_mux_bus_95,
  input         io_i_mux_bus_96,
  input         io_i_mux_bus_97,
  input         io_i_mux_bus_98,
  input         io_i_mux_bus_99,
  input         io_i_mux_bus_100,
  input         io_i_mux_bus_101,
  input         io_i_mux_bus_102,
  input         io_i_mux_bus_103,
  input         io_i_mux_bus_104,
  input         io_i_mux_bus_105,
  input         io_i_mux_bus_106,
  input         io_i_mux_bus_107,
  input         io_i_mux_bus_108,
  input         io_i_mux_bus_109,
  input         io_i_mux_bus_110,
  input         io_i_mux_bus_111,
  input         io_i_mux_bus_112,
  input         io_i_mux_bus_113,
  input         io_i_mux_bus_114,
  input         io_i_mux_bus_115,
  input         io_i_mux_bus_116,
  input         io_i_mux_bus_117,
  input         io_i_mux_bus_118,
  input         io_i_mux_bus_119,
  input         io_i_mux_bus_120,
  input         io_i_mux_bus_121,
  input         io_i_mux_bus_122,
  input         io_i_mux_bus_123,
  input         io_i_mux_bus_124,
  input         io_i_mux_bus_125,
  input         io_i_mux_bus_126,
  input         io_i_mux_bus_127,
  input         io_i_mux_bus_128,
  input         io_i_mux_bus_129,
  input         io_i_mux_bus_130,
  input         io_i_mux_bus_131,
  input         io_i_mux_bus_132,
  input         io_i_mux_bus_133,
  input         io_i_mux_bus_134,
  input         io_i_mux_bus_135,
  input         io_i_mux_bus_136,
  input         io_i_mux_bus_137,
  input         io_i_mux_bus_138,
  input         io_i_mux_bus_139,
  input         io_i_mux_bus_140,
  input         io_i_mux_bus_141,
  input         io_i_mux_bus_142,
  input         io_i_mux_bus_143,
  input         io_i_mux_bus_144,
  input         io_i_mux_bus_145,
  input         io_i_mux_bus_146,
  input         io_i_mux_bus_147,
  input         io_i_mux_bus_148,
  input         io_i_mux_bus_149,
  input         io_i_mux_bus_150,
  input         io_i_mux_bus_151,
  input         io_i_mux_bus_152,
  input         io_i_mux_bus_153,
  input         io_i_mux_bus_154,
  input         io_i_mux_bus_155,
  input         io_i_mux_bus_156,
  input         io_i_mux_bus_157,
  input         io_i_mux_bus_158,
  input         io_i_mux_bus_159,
  input         io_i_mux_bus_160,
  input         io_i_mux_bus_161,
  input         io_i_mux_bus_162,
  input         io_i_mux_bus_163,
  input         io_i_mux_bus_164,
  input         io_i_mux_bus_165,
  input         io_i_mux_bus_166,
  input         io_i_mux_bus_167,
  input         io_i_mux_bus_168,
  input         io_i_mux_bus_169,
  input         io_i_mux_bus_170,
  input         io_i_mux_bus_171,
  input         io_i_mux_bus_172,
  input         io_i_mux_bus_173,
  input         io_i_mux_bus_174,
  input         io_i_mux_bus_175,
  input         io_i_mux_bus_176,
  input         io_i_mux_bus_177,
  input         io_i_mux_bus_178,
  input         io_i_mux_bus_179,
  input         io_i_mux_bus_180,
  input         io_i_mux_bus_181,
  input         io_i_mux_bus_182,
  input         io_i_mux_bus_183,
  input         io_i_mux_bus_184,
  input         io_i_mux_bus_185,
  input         io_i_mux_bus_186,
  input         io_i_mux_bus_187,
  input         io_i_mux_bus_188,
  input         io_i_mux_bus_189,
  input         io_i_mux_bus_190,
  input         io_i_mux_bus_191,
  input         io_i_mux_bus_192,
  input         io_i_mux_bus_193,
  input         io_i_mux_bus_194,
  input         io_i_mux_bus_195,
  input         io_i_mux_bus_196,
  input         io_i_mux_bus_197,
  input         io_i_mux_bus_198,
  input         io_i_mux_bus_199,
  input         io_i_mux_bus_200,
  input         io_i_mux_bus_201,
  input         io_i_mux_bus_202,
  input         io_i_mux_bus_203,
  input         io_i_mux_bus_204,
  input         io_i_mux_bus_205,
  input         io_i_mux_bus_206,
  input         io_i_mux_bus_207,
  input         io_i_mux_bus_208,
  input         io_i_mux_bus_209,
  input         io_i_mux_bus_210,
  input         io_i_mux_bus_211,
  input         io_i_mux_bus_212,
  input         io_i_mux_bus_213,
  input         io_i_mux_bus_214,
  input         io_i_mux_bus_215,
  input         io_i_mux_bus_216,
  input         io_i_mux_bus_217,
  input         io_i_mux_bus_218,
  input         io_i_mux_bus_219,
  input         io_i_mux_bus_220,
  input         io_i_mux_bus_221,
  input         io_i_mux_bus_222,
  input         io_i_mux_bus_223,
  input         io_i_mux_bus_224,
  input         io_i_mux_bus_225,
  input         io_i_mux_bus_226,
  input         io_i_mux_bus_227,
  input         io_i_mux_bus_228,
  input         io_i_mux_bus_229,
  input         io_i_mux_bus_230,
  input         io_i_mux_bus_231,
  input         io_i_mux_bus_232,
  input         io_i_mux_bus_233,
  input         io_i_mux_bus_234,
  input         io_i_mux_bus_235,
  input         io_i_mux_bus_236,
  input         io_i_mux_bus_237,
  input         io_i_mux_bus_238,
  input         io_i_mux_bus_239,
  input         io_i_mux_bus_240,
  input         io_i_mux_bus_241,
  input         io_i_mux_bus_242,
  input         io_i_mux_bus_243,
  input         io_i_mux_bus_244,
  input         io_i_mux_bus_245,
  input         io_i_mux_bus_246,
  input         io_i_mux_bus_247,
  input         io_i_mux_bus_248,
  input         io_i_mux_bus_249,
  input         io_i_mux_bus_250,
  input         io_i_mux_bus_251,
  input         io_i_mux_bus_252,
  input         io_i_mux_bus_253,
  input         io_i_mux_bus_254,
  input         io_i_mux_bus_255,
  input         io_i_mux_bus_256,
  input         io_i_mux_bus_257,
  input         io_i_mux_bus_258,
  input         io_i_mux_bus_259,
  input         io_i_mux_bus_260,
  input         io_i_mux_bus_261,
  input         io_i_mux_bus_262,
  input         io_i_mux_bus_263,
  input         io_i_mux_bus_264,
  input         io_i_mux_bus_265,
  input         io_i_mux_bus_266,
  input         io_i_mux_bus_267,
  input         io_i_mux_bus_268,
  input         io_i_mux_bus_269,
  input         io_i_mux_bus_270,
  input         io_i_mux_bus_271,
  input         io_i_mux_bus_272,
  input         io_i_mux_bus_273,
  input         io_i_mux_bus_274,
  input         io_i_mux_bus_275,
  input         io_i_mux_bus_276,
  input         io_i_mux_bus_277,
  input         io_i_mux_bus_278,
  input         io_i_mux_bus_279,
  input         io_i_mux_bus_280,
  input         io_i_mux_bus_281,
  input         io_i_mux_bus_282,
  input         io_i_mux_bus_283,
  input         io_i_mux_bus_284,
  input         io_i_mux_bus_285,
  input         io_i_mux_bus_286,
  input         io_i_mux_bus_287,
  input         io_i_mux_bus_288,
  input         io_i_mux_bus_289,
  input         io_i_mux_bus_290,
  input         io_i_mux_bus_291,
  input         io_i_mux_bus_292,
  input         io_i_mux_bus_293,
  input         io_i_mux_bus_294,
  input         io_i_mux_bus_295,
  input         io_i_mux_bus_296,
  input         io_i_mux_bus_297,
  input         io_i_mux_bus_298,
  input         io_i_mux_bus_299,
  input         io_i_mux_bus_300,
  input         io_i_mux_bus_301,
  input         io_i_mux_bus_302,
  input         io_i_mux_bus_303,
  input         io_i_mux_bus_304,
  input         io_i_mux_bus_305,
  input         io_i_mux_bus_306,
  input         io_i_mux_bus_307,
  input         io_i_mux_bus_308,
  input         io_i_mux_bus_309,
  input         io_i_mux_bus_310,
  input         io_i_mux_bus_311,
  input         io_i_mux_bus_312,
  input         io_i_mux_bus_313,
  input         io_i_mux_bus_314,
  input         io_i_mux_bus_315,
  input         io_i_mux_bus_316,
  input         io_i_mux_bus_317,
  input         io_i_mux_bus_318,
  input         io_i_mux_bus_319,
  input         io_i_mux_bus_320,
  input         io_i_mux_bus_321,
  input         io_i_mux_bus_322,
  input         io_i_mux_bus_323,
  input         io_i_mux_bus_324,
  input         io_i_mux_bus_325,
  input         io_i_mux_bus_326,
  input         io_i_mux_bus_327,
  input         io_i_mux_bus_328,
  input         io_i_mux_bus_329,
  input         io_i_mux_bus_330,
  input         io_i_mux_bus_331,
  input         io_i_mux_bus_332,
  input         io_i_mux_bus_333,
  input         io_i_mux_bus_334,
  input         io_i_mux_bus_335,
  input         io_i_mux_bus_336,
  input         io_i_mux_bus_337,
  input         io_i_mux_bus_338,
  input         io_i_mux_bus_339,
  input         io_i_mux_bus_340,
  input         io_i_mux_bus_341,
  input         io_i_mux_bus_342,
  input         io_i_mux_bus_343,
  input         io_i_mux_bus_344,
  input         io_i_mux_bus_345,
  input         io_i_mux_bus_346,
  input         io_i_mux_bus_347,
  input         io_i_mux_bus_348,
  input         io_i_mux_bus_349,
  input         io_i_mux_bus_350,
  input         io_i_mux_bus_351,
  input         io_i_mux_bus_352,
  input         io_i_mux_bus_353,
  input         io_i_mux_bus_354,
  input         io_i_mux_bus_355,
  input         io_i_mux_bus_356,
  input         io_i_mux_bus_357,
  input         io_i_mux_bus_358,
  input         io_i_mux_bus_359,
  input         io_i_mux_bus_360,
  input         io_i_mux_bus_361,
  input         io_i_mux_bus_362,
  input         io_i_mux_bus_363,
  input         io_i_mux_bus_364,
  input         io_i_mux_bus_365,
  input         io_i_mux_bus_366,
  input         io_i_mux_bus_367,
  input         io_i_mux_bus_368,
  input         io_i_mux_bus_369,
  input         io_i_mux_bus_370,
  input         io_i_mux_bus_371,
  input         io_i_mux_bus_372,
  input         io_i_mux_bus_373,
  input         io_i_mux_bus_374,
  input         io_i_mux_bus_375,
  input         io_i_mux_bus_376,
  input         io_i_mux_bus_377,
  input         io_i_mux_bus_378,
  input         io_i_mux_bus_379,
  input         io_i_mux_bus_380,
  input         io_i_mux_bus_381,
  input         io_i_mux_bus_382,
  input         io_i_mux_bus_383,
  input         io_i_mux_bus_384,
  input         io_i_mux_bus_385,
  input         io_i_mux_bus_386,
  input         io_i_mux_bus_387,
  input         io_i_mux_bus_388,
  input         io_i_mux_bus_389,
  input         io_i_mux_bus_390,
  input         io_i_mux_bus_391,
  input         io_i_mux_bus_392,
  input         io_i_mux_bus_393,
  input         io_i_mux_bus_394,
  input         io_i_mux_bus_395,
  input         io_i_mux_bus_396,
  input         io_i_mux_bus_397,
  input         io_i_mux_bus_398,
  input         io_i_mux_bus_399,
  input         io_i_mux_bus_400,
  input         io_i_mux_bus_401,
  input         io_i_mux_bus_402,
  input         io_i_mux_bus_403,
  input         io_i_mux_bus_404,
  input         io_i_mux_bus_405,
  input         io_i_mux_bus_406,
  input         io_i_mux_bus_407,
  input         io_i_mux_bus_408,
  input         io_i_mux_bus_409,
  input         io_i_mux_bus_410,
  input         io_i_mux_bus_411,
  input         io_i_mux_bus_412,
  input         io_i_mux_bus_413,
  input         io_i_mux_bus_414,
  input         io_i_mux_bus_415,
  input         io_i_mux_bus_416,
  input         io_i_mux_bus_417,
  input         io_i_mux_bus_418,
  input         io_i_mux_bus_419,
  input         io_i_mux_bus_420,
  input         io_i_mux_bus_421,
  input         io_i_mux_bus_422,
  input         io_i_mux_bus_423,
  input         io_i_mux_bus_424,
  input         io_i_mux_bus_425,
  input         io_i_mux_bus_426,
  input         io_i_mux_bus_427,
  input         io_i_mux_bus_428,
  input         io_i_mux_bus_429,
  input         io_i_mux_bus_430,
  input         io_i_mux_bus_431,
  input         io_i_mux_bus_432,
  input         io_i_mux_bus_433,
  input         io_i_mux_bus_434,
  input         io_i_mux_bus_435,
  input         io_i_mux_bus_436,
  input         io_i_mux_bus_437,
  input         io_i_mux_bus_438,
  input         io_i_mux_bus_439,
  input         io_i_mux_bus_440,
  input         io_i_mux_bus_441,
  input         io_i_mux_bus_442,
  input         io_i_mux_bus_443,
  input         io_i_mux_bus_444,
  input         io_i_mux_bus_445,
  input         io_i_mux_bus_446,
  input         io_i_mux_bus_447,
  input         io_i_mux_bus_448,
  input         io_i_mux_bus_449,
  input         io_i_mux_bus_450,
  input         io_i_mux_bus_451,
  input         io_i_mux_bus_452,
  input         io_i_mux_bus_453,
  input         io_i_mux_bus_454,
  input         io_i_mux_bus_455,
  input         io_i_mux_bus_456,
  input         io_i_mux_bus_457,
  input         io_i_mux_bus_458,
  input         io_i_mux_bus_459,
  input         io_i_mux_bus_460,
  input         io_i_mux_bus_461,
  input         io_i_mux_bus_462,
  input         io_i_mux_bus_463,
  input         io_i_mux_bus_464,
  input         io_i_mux_bus_465,
  input         io_i_mux_bus_466,
  input         io_i_mux_bus_467,
  input         io_i_mux_bus_468,
  input         io_i_mux_bus_469,
  input         io_i_mux_bus_470,
  input         io_i_mux_bus_471,
  input         io_i_mux_bus_472,
  input         io_i_mux_bus_473,
  input         io_i_mux_bus_474,
  input         io_i_mux_bus_475,
  input         io_i_mux_bus_476,
  input         io_i_mux_bus_477,
  input         io_i_mux_bus_478,
  input         io_i_mux_bus_479,
  input         io_i_mux_bus_480,
  input         io_i_mux_bus_481,
  input         io_i_mux_bus_482,
  input         io_i_mux_bus_483,
  input         io_i_mux_bus_484,
  input         io_i_mux_bus_485,
  input         io_i_mux_bus_486,
  input         io_i_mux_bus_487,
  input         io_i_mux_bus_488,
  input         io_i_mux_bus_489,
  input         io_i_mux_bus_490,
  input         io_i_mux_bus_491,
  input         io_i_mux_bus_492,
  input         io_i_mux_bus_493,
  input         io_i_mux_bus_494,
  input         io_i_mux_bus_495,
  input         io_i_mux_bus_496,
  input         io_i_mux_bus_497,
  input         io_i_mux_bus_498,
  input         io_i_mux_bus_499,
  input         io_i_mux_bus_500,
  input         io_i_mux_bus_501,
  input         io_i_mux_bus_502,
  input         io_i_mux_bus_503,
  input         io_i_mux_bus_504,
  input         io_i_mux_bus_505,
  input         io_i_mux_bus_506,
  input         io_i_mux_bus_507,
  input         io_i_mux_bus_508,
  input         io_i_mux_bus_509,
  input         io_i_mux_bus_510,
  input         io_i_mux_bus_511,
  input         io_i_mux_bus_512,
  input         io_i_mux_bus_513,
  input         io_i_mux_bus_514,
  input         io_i_mux_bus_515,
  input         io_i_mux_bus_516,
  input         io_i_mux_bus_517,
  input         io_i_mux_bus_518,
  input         io_i_mux_bus_519,
  input         io_i_mux_bus_520,
  input         io_i_mux_bus_521,
  input         io_i_mux_bus_522,
  input         io_i_mux_bus_523,
  input         io_i_mux_bus_524,
  input         io_i_mux_bus_525,
  input         io_i_mux_bus_526,
  input         io_i_mux_bus_527,
  input         io_i_mux_bus_528,
  input         io_i_mux_bus_529,
  input         io_i_mux_bus_530,
  input         io_i_mux_bus_531,
  input         io_i_mux_bus_532,
  input         io_i_mux_bus_533,
  input         io_i_mux_bus_534,
  input         io_i_mux_bus_535,
  input         io_i_mux_bus_536,
  input         io_i_mux_bus_537,
  input         io_i_mux_bus_538,
  input         io_i_mux_bus_539,
  input         io_i_mux_bus_540,
  input         io_i_mux_bus_541,
  input         io_i_mux_bus_542,
  input         io_i_mux_bus_543,
  input         io_i_mux_bus_544,
  input         io_i_mux_bus_545,
  input         io_i_mux_bus_546,
  input         io_i_mux_bus_547,
  input         io_i_mux_bus_548,
  input         io_i_mux_bus_549,
  input         io_i_mux_bus_550,
  input         io_i_mux_bus_551,
  input         io_i_mux_bus_552,
  input         io_i_mux_bus_553,
  input         io_i_mux_bus_554,
  input         io_i_mux_bus_555,
  input         io_i_mux_bus_556,
  input         io_i_mux_bus_557,
  input         io_i_mux_bus_558,
  input         io_i_mux_bus_559,
  input         io_i_mux_bus_560,
  input         io_i_mux_bus_561,
  input         io_i_mux_bus_562,
  input         io_i_mux_bus_563,
  input         io_i_mux_bus_564,
  input         io_i_mux_bus_565,
  input         io_i_mux_bus_566,
  input         io_i_mux_bus_567,
  input         io_i_mux_bus_568,
  input         io_i_mux_bus_569,
  input         io_i_mux_bus_570,
  input         io_i_mux_bus_571,
  input         io_i_mux_bus_572,
  input         io_i_mux_bus_573,
  input         io_i_mux_bus_574,
  input         io_i_mux_bus_575,
  input         io_i_mux_bus_576,
  input         io_i_mux_bus_577,
  input         io_i_mux_bus_578,
  input         io_i_mux_bus_579,
  input         io_i_mux_bus_580,
  input         io_i_mux_bus_581,
  input         io_i_mux_bus_582,
  input         io_i_mux_bus_583,
  input         io_i_mux_bus_584,
  input         io_i_mux_bus_585,
  input         io_i_mux_bus_586,
  input         io_i_mux_bus_587,
  input         io_i_mux_bus_588,
  input         io_i_mux_bus_589,
  input         io_i_mux_bus_590,
  input         io_i_mux_bus_591,
  input         io_i_mux_bus_592,
  input         io_i_mux_bus_593,
  input         io_i_mux_bus_594,
  input         io_i_mux_bus_595,
  input         io_i_mux_bus_596,
  input         io_i_mux_bus_597,
  input         io_i_mux_bus_598,
  input         io_i_mux_bus_599,
  input         io_i_mux_bus_600,
  input         io_i_mux_bus_601,
  input         io_i_mux_bus_602,
  input         io_i_mux_bus_603,
  input         io_i_mux_bus_604,
  input         io_i_mux_bus_605,
  input         io_i_mux_bus_606,
  input         io_i_mux_bus_607,
  output [31:0] io_o_dist_bus_0,
  output [31:0] io_o_dist_bus_1,
  output [31:0] io_o_dist_bus_2,
  output [31:0] io_o_dist_bus_3,
  output [31:0] io_o_dist_bus_4,
  output [31:0] io_o_dist_bus_5,
  output [31:0] io_o_dist_bus_6,
  output [31:0] io_o_dist_bus_7,
  output [31:0] io_o_dist_bus_8,
  output [31:0] io_o_dist_bus_9,
  output [31:0] io_o_dist_bus_10,
  output [31:0] io_o_dist_bus_11,
  output [31:0] io_o_dist_bus_12,
  output [31:0] io_o_dist_bus_13,
  output [31:0] io_o_dist_bus_14,
  output [31:0] io_o_dist_bus_15,
  output [31:0] io_o_dist_bus_16,
  output [31:0] io_o_dist_bus_17,
  output [31:0] io_o_dist_bus_18,
  output [31:0] io_o_dist_bus_19,
  output [31:0] io_o_dist_bus_20,
  output [31:0] io_o_dist_bus_21,
  output [31:0] io_o_dist_bus_22,
  output [31:0] io_o_dist_bus_23,
  output [31:0] io_o_dist_bus_24,
  output [31:0] io_o_dist_bus_25,
  output [31:0] io_o_dist_bus_26,
  output [31:0] io_o_dist_bus_27,
  output [31:0] io_o_dist_bus_28,
  output [31:0] io_o_dist_bus_29,
  output [31:0] io_o_dist_bus_30,
  output [31:0] io_o_dist_bus_31
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] in_switch_io_y; // @[Benes.scala 89:27]
  wire [31:0] in_switch_io_z; // @[Benes.scala 89:27]
  wire [31:0] in_switch_io_in; // @[Benes.scala 89:27]
  wire [31:0] in_switch_1_io_y; // @[Benes.scala 89:27]
  wire [31:0] in_switch_1_io_z; // @[Benes.scala 89:27]
  wire [31:0] in_switch_1_io_in; // @[Benes.scala 89:27]
  wire [31:0] in_switch_2_io_y; // @[Benes.scala 89:27]
  wire [31:0] in_switch_2_io_z; // @[Benes.scala 89:27]
  wire [31:0] in_switch_2_io_in; // @[Benes.scala 89:27]
  wire [31:0] in_switch_3_io_y; // @[Benes.scala 89:27]
  wire [31:0] in_switch_3_io_z; // @[Benes.scala 89:27]
  wire [31:0] in_switch_3_io_in; // @[Benes.scala 89:27]
  wire [31:0] in_switch_4_io_y; // @[Benes.scala 89:27]
  wire [31:0] in_switch_4_io_z; // @[Benes.scala 89:27]
  wire [31:0] in_switch_4_io_in; // @[Benes.scala 89:27]
  wire [31:0] in_switch_5_io_y; // @[Benes.scala 89:27]
  wire [31:0] in_switch_5_io_z; // @[Benes.scala 89:27]
  wire [31:0] in_switch_5_io_in; // @[Benes.scala 89:27]
  wire [31:0] in_switch_6_io_y; // @[Benes.scala 89:27]
  wire [31:0] in_switch_6_io_z; // @[Benes.scala 89:27]
  wire [31:0] in_switch_6_io_in; // @[Benes.scala 89:27]
  wire [31:0] in_switch_7_io_y; // @[Benes.scala 89:27]
  wire [31:0] in_switch_7_io_z; // @[Benes.scala 89:27]
  wire [31:0] in_switch_7_io_in; // @[Benes.scala 89:27]
  wire [31:0] in_switch_8_io_y; // @[Benes.scala 89:27]
  wire [31:0] in_switch_8_io_z; // @[Benes.scala 89:27]
  wire [31:0] in_switch_8_io_in; // @[Benes.scala 89:27]
  wire [31:0] in_switch_9_io_y; // @[Benes.scala 89:27]
  wire [31:0] in_switch_9_io_z; // @[Benes.scala 89:27]
  wire [31:0] in_switch_9_io_in; // @[Benes.scala 89:27]
  wire [31:0] in_switch_10_io_y; // @[Benes.scala 89:27]
  wire [31:0] in_switch_10_io_z; // @[Benes.scala 89:27]
  wire [31:0] in_switch_10_io_in; // @[Benes.scala 89:27]
  wire [31:0] in_switch_11_io_y; // @[Benes.scala 89:27]
  wire [31:0] in_switch_11_io_z; // @[Benes.scala 89:27]
  wire [31:0] in_switch_11_io_in; // @[Benes.scala 89:27]
  wire [31:0] in_switch_12_io_y; // @[Benes.scala 89:27]
  wire [31:0] in_switch_12_io_z; // @[Benes.scala 89:27]
  wire [31:0] in_switch_12_io_in; // @[Benes.scala 89:27]
  wire [31:0] in_switch_13_io_y; // @[Benes.scala 89:27]
  wire [31:0] in_switch_13_io_z; // @[Benes.scala 89:27]
  wire [31:0] in_switch_13_io_in; // @[Benes.scala 89:27]
  wire [31:0] in_switch_14_io_y; // @[Benes.scala 89:27]
  wire [31:0] in_switch_14_io_z; // @[Benes.scala 89:27]
  wire [31:0] in_switch_14_io_in; // @[Benes.scala 89:27]
  wire [31:0] in_switch_15_io_y; // @[Benes.scala 89:27]
  wire [31:0] in_switch_15_io_z; // @[Benes.scala 89:27]
  wire [31:0] in_switch_15_io_in; // @[Benes.scala 89:27]
  wire [31:0] in_switch_16_io_y; // @[Benes.scala 89:27]
  wire [31:0] in_switch_16_io_z; // @[Benes.scala 89:27]
  wire [31:0] in_switch_16_io_in; // @[Benes.scala 89:27]
  wire [31:0] in_switch_17_io_y; // @[Benes.scala 89:27]
  wire [31:0] in_switch_17_io_z; // @[Benes.scala 89:27]
  wire [31:0] in_switch_17_io_in; // @[Benes.scala 89:27]
  wire [31:0] in_switch_18_io_y; // @[Benes.scala 89:27]
  wire [31:0] in_switch_18_io_z; // @[Benes.scala 89:27]
  wire [31:0] in_switch_18_io_in; // @[Benes.scala 89:27]
  wire [31:0] in_switch_19_io_y; // @[Benes.scala 89:27]
  wire [31:0] in_switch_19_io_z; // @[Benes.scala 89:27]
  wire [31:0] in_switch_19_io_in; // @[Benes.scala 89:27]
  wire [31:0] in_switch_20_io_y; // @[Benes.scala 89:27]
  wire [31:0] in_switch_20_io_z; // @[Benes.scala 89:27]
  wire [31:0] in_switch_20_io_in; // @[Benes.scala 89:27]
  wire [31:0] in_switch_21_io_y; // @[Benes.scala 89:27]
  wire [31:0] in_switch_21_io_z; // @[Benes.scala 89:27]
  wire [31:0] in_switch_21_io_in; // @[Benes.scala 89:27]
  wire [31:0] in_switch_22_io_y; // @[Benes.scala 89:27]
  wire [31:0] in_switch_22_io_z; // @[Benes.scala 89:27]
  wire [31:0] in_switch_22_io_in; // @[Benes.scala 89:27]
  wire [31:0] in_switch_23_io_y; // @[Benes.scala 89:27]
  wire [31:0] in_switch_23_io_z; // @[Benes.scala 89:27]
  wire [31:0] in_switch_23_io_in; // @[Benes.scala 89:27]
  wire [31:0] in_switch_24_io_y; // @[Benes.scala 89:27]
  wire [31:0] in_switch_24_io_z; // @[Benes.scala 89:27]
  wire [31:0] in_switch_24_io_in; // @[Benes.scala 89:27]
  wire [31:0] in_switch_25_io_y; // @[Benes.scala 89:27]
  wire [31:0] in_switch_25_io_z; // @[Benes.scala 89:27]
  wire [31:0] in_switch_25_io_in; // @[Benes.scala 89:27]
  wire [31:0] in_switch_26_io_y; // @[Benes.scala 89:27]
  wire [31:0] in_switch_26_io_z; // @[Benes.scala 89:27]
  wire [31:0] in_switch_26_io_in; // @[Benes.scala 89:27]
  wire [31:0] in_switch_27_io_y; // @[Benes.scala 89:27]
  wire [31:0] in_switch_27_io_z; // @[Benes.scala 89:27]
  wire [31:0] in_switch_27_io_in; // @[Benes.scala 89:27]
  wire [31:0] in_switch_28_io_y; // @[Benes.scala 89:27]
  wire [31:0] in_switch_28_io_z; // @[Benes.scala 89:27]
  wire [31:0] in_switch_28_io_in; // @[Benes.scala 89:27]
  wire [31:0] in_switch_29_io_y; // @[Benes.scala 89:27]
  wire [31:0] in_switch_29_io_z; // @[Benes.scala 89:27]
  wire [31:0] in_switch_29_io_in; // @[Benes.scala 89:27]
  wire [31:0] in_switch_30_io_y; // @[Benes.scala 89:27]
  wire [31:0] in_switch_30_io_z; // @[Benes.scala 89:27]
  wire [31:0] in_switch_30_io_in; // @[Benes.scala 89:27]
  wire [31:0] in_switch_31_io_y; // @[Benes.scala 89:27]
  wire [31:0] in_switch_31_io_z; // @[Benes.scala 89:27]
  wire [31:0] in_switch_31_io_in; // @[Benes.scala 89:27]
  wire [31:0] out_switch_io_y; // @[Benes.scala 98:28]
  wire [31:0] out_switch_io_in0; // @[Benes.scala 98:28]
  wire [31:0] out_switch_io_in1; // @[Benes.scala 98:28]
  wire  out_switch_io_sel; // @[Benes.scala 98:28]
  wire [31:0] out_switch_1_io_y; // @[Benes.scala 98:28]
  wire [31:0] out_switch_1_io_in0; // @[Benes.scala 98:28]
  wire [31:0] out_switch_1_io_in1; // @[Benes.scala 98:28]
  wire  out_switch_1_io_sel; // @[Benes.scala 98:28]
  wire [31:0] out_switch_2_io_y; // @[Benes.scala 98:28]
  wire [31:0] out_switch_2_io_in0; // @[Benes.scala 98:28]
  wire [31:0] out_switch_2_io_in1; // @[Benes.scala 98:28]
  wire  out_switch_2_io_sel; // @[Benes.scala 98:28]
  wire [31:0] out_switch_3_io_y; // @[Benes.scala 98:28]
  wire [31:0] out_switch_3_io_in0; // @[Benes.scala 98:28]
  wire [31:0] out_switch_3_io_in1; // @[Benes.scala 98:28]
  wire  out_switch_3_io_sel; // @[Benes.scala 98:28]
  wire [31:0] out_switch_4_io_y; // @[Benes.scala 98:28]
  wire [31:0] out_switch_4_io_in0; // @[Benes.scala 98:28]
  wire [31:0] out_switch_4_io_in1; // @[Benes.scala 98:28]
  wire  out_switch_4_io_sel; // @[Benes.scala 98:28]
  wire [31:0] out_switch_5_io_y; // @[Benes.scala 98:28]
  wire [31:0] out_switch_5_io_in0; // @[Benes.scala 98:28]
  wire [31:0] out_switch_5_io_in1; // @[Benes.scala 98:28]
  wire  out_switch_5_io_sel; // @[Benes.scala 98:28]
  wire [31:0] out_switch_6_io_y; // @[Benes.scala 98:28]
  wire [31:0] out_switch_6_io_in0; // @[Benes.scala 98:28]
  wire [31:0] out_switch_6_io_in1; // @[Benes.scala 98:28]
  wire  out_switch_6_io_sel; // @[Benes.scala 98:28]
  wire [31:0] out_switch_7_io_y; // @[Benes.scala 98:28]
  wire [31:0] out_switch_7_io_in0; // @[Benes.scala 98:28]
  wire [31:0] out_switch_7_io_in1; // @[Benes.scala 98:28]
  wire  out_switch_7_io_sel; // @[Benes.scala 98:28]
  wire [31:0] out_switch_8_io_y; // @[Benes.scala 98:28]
  wire [31:0] out_switch_8_io_in0; // @[Benes.scala 98:28]
  wire [31:0] out_switch_8_io_in1; // @[Benes.scala 98:28]
  wire  out_switch_8_io_sel; // @[Benes.scala 98:28]
  wire [31:0] out_switch_9_io_y; // @[Benes.scala 98:28]
  wire [31:0] out_switch_9_io_in0; // @[Benes.scala 98:28]
  wire [31:0] out_switch_9_io_in1; // @[Benes.scala 98:28]
  wire  out_switch_9_io_sel; // @[Benes.scala 98:28]
  wire [31:0] out_switch_10_io_y; // @[Benes.scala 98:28]
  wire [31:0] out_switch_10_io_in0; // @[Benes.scala 98:28]
  wire [31:0] out_switch_10_io_in1; // @[Benes.scala 98:28]
  wire  out_switch_10_io_sel; // @[Benes.scala 98:28]
  wire [31:0] out_switch_11_io_y; // @[Benes.scala 98:28]
  wire [31:0] out_switch_11_io_in0; // @[Benes.scala 98:28]
  wire [31:0] out_switch_11_io_in1; // @[Benes.scala 98:28]
  wire  out_switch_11_io_sel; // @[Benes.scala 98:28]
  wire [31:0] out_switch_12_io_y; // @[Benes.scala 98:28]
  wire [31:0] out_switch_12_io_in0; // @[Benes.scala 98:28]
  wire [31:0] out_switch_12_io_in1; // @[Benes.scala 98:28]
  wire  out_switch_12_io_sel; // @[Benes.scala 98:28]
  wire [31:0] out_switch_13_io_y; // @[Benes.scala 98:28]
  wire [31:0] out_switch_13_io_in0; // @[Benes.scala 98:28]
  wire [31:0] out_switch_13_io_in1; // @[Benes.scala 98:28]
  wire  out_switch_13_io_sel; // @[Benes.scala 98:28]
  wire [31:0] out_switch_14_io_y; // @[Benes.scala 98:28]
  wire [31:0] out_switch_14_io_in0; // @[Benes.scala 98:28]
  wire [31:0] out_switch_14_io_in1; // @[Benes.scala 98:28]
  wire  out_switch_14_io_sel; // @[Benes.scala 98:28]
  wire [31:0] out_switch_15_io_y; // @[Benes.scala 98:28]
  wire [31:0] out_switch_15_io_in0; // @[Benes.scala 98:28]
  wire [31:0] out_switch_15_io_in1; // @[Benes.scala 98:28]
  wire  out_switch_15_io_sel; // @[Benes.scala 98:28]
  wire [31:0] out_switch_16_io_y; // @[Benes.scala 98:28]
  wire [31:0] out_switch_16_io_in0; // @[Benes.scala 98:28]
  wire [31:0] out_switch_16_io_in1; // @[Benes.scala 98:28]
  wire  out_switch_16_io_sel; // @[Benes.scala 98:28]
  wire [31:0] out_switch_17_io_y; // @[Benes.scala 98:28]
  wire [31:0] out_switch_17_io_in0; // @[Benes.scala 98:28]
  wire [31:0] out_switch_17_io_in1; // @[Benes.scala 98:28]
  wire  out_switch_17_io_sel; // @[Benes.scala 98:28]
  wire [31:0] out_switch_18_io_y; // @[Benes.scala 98:28]
  wire [31:0] out_switch_18_io_in0; // @[Benes.scala 98:28]
  wire [31:0] out_switch_18_io_in1; // @[Benes.scala 98:28]
  wire  out_switch_18_io_sel; // @[Benes.scala 98:28]
  wire [31:0] out_switch_19_io_y; // @[Benes.scala 98:28]
  wire [31:0] out_switch_19_io_in0; // @[Benes.scala 98:28]
  wire [31:0] out_switch_19_io_in1; // @[Benes.scala 98:28]
  wire  out_switch_19_io_sel; // @[Benes.scala 98:28]
  wire [31:0] out_switch_20_io_y; // @[Benes.scala 98:28]
  wire [31:0] out_switch_20_io_in0; // @[Benes.scala 98:28]
  wire [31:0] out_switch_20_io_in1; // @[Benes.scala 98:28]
  wire  out_switch_20_io_sel; // @[Benes.scala 98:28]
  wire [31:0] out_switch_21_io_y; // @[Benes.scala 98:28]
  wire [31:0] out_switch_21_io_in0; // @[Benes.scala 98:28]
  wire [31:0] out_switch_21_io_in1; // @[Benes.scala 98:28]
  wire  out_switch_21_io_sel; // @[Benes.scala 98:28]
  wire [31:0] out_switch_22_io_y; // @[Benes.scala 98:28]
  wire [31:0] out_switch_22_io_in0; // @[Benes.scala 98:28]
  wire [31:0] out_switch_22_io_in1; // @[Benes.scala 98:28]
  wire  out_switch_22_io_sel; // @[Benes.scala 98:28]
  wire [31:0] out_switch_23_io_y; // @[Benes.scala 98:28]
  wire [31:0] out_switch_23_io_in0; // @[Benes.scala 98:28]
  wire [31:0] out_switch_23_io_in1; // @[Benes.scala 98:28]
  wire  out_switch_23_io_sel; // @[Benes.scala 98:28]
  wire [31:0] out_switch_24_io_y; // @[Benes.scala 98:28]
  wire [31:0] out_switch_24_io_in0; // @[Benes.scala 98:28]
  wire [31:0] out_switch_24_io_in1; // @[Benes.scala 98:28]
  wire  out_switch_24_io_sel; // @[Benes.scala 98:28]
  wire [31:0] out_switch_25_io_y; // @[Benes.scala 98:28]
  wire [31:0] out_switch_25_io_in0; // @[Benes.scala 98:28]
  wire [31:0] out_switch_25_io_in1; // @[Benes.scala 98:28]
  wire  out_switch_25_io_sel; // @[Benes.scala 98:28]
  wire [31:0] out_switch_26_io_y; // @[Benes.scala 98:28]
  wire [31:0] out_switch_26_io_in0; // @[Benes.scala 98:28]
  wire [31:0] out_switch_26_io_in1; // @[Benes.scala 98:28]
  wire  out_switch_26_io_sel; // @[Benes.scala 98:28]
  wire [31:0] out_switch_27_io_y; // @[Benes.scala 98:28]
  wire [31:0] out_switch_27_io_in0; // @[Benes.scala 98:28]
  wire [31:0] out_switch_27_io_in1; // @[Benes.scala 98:28]
  wire  out_switch_27_io_sel; // @[Benes.scala 98:28]
  wire [31:0] out_switch_28_io_y; // @[Benes.scala 98:28]
  wire [31:0] out_switch_28_io_in0; // @[Benes.scala 98:28]
  wire [31:0] out_switch_28_io_in1; // @[Benes.scala 98:28]
  wire  out_switch_28_io_sel; // @[Benes.scala 98:28]
  wire [31:0] out_switch_29_io_y; // @[Benes.scala 98:28]
  wire [31:0] out_switch_29_io_in0; // @[Benes.scala 98:28]
  wire [31:0] out_switch_29_io_in1; // @[Benes.scala 98:28]
  wire  out_switch_29_io_sel; // @[Benes.scala 98:28]
  wire [31:0] out_switch_30_io_y; // @[Benes.scala 98:28]
  wire [31:0] out_switch_30_io_in0; // @[Benes.scala 98:28]
  wire [31:0] out_switch_30_io_in1; // @[Benes.scala 98:28]
  wire  out_switch_30_io_sel; // @[Benes.scala 98:28]
  wire [31:0] out_switch_31_io_y; // @[Benes.scala 98:28]
  wire [31:0] out_switch_31_io_in0; // @[Benes.scala 98:28]
  wire [31:0] out_switch_31_io_in1; // @[Benes.scala 98:28]
  wire  out_switch_31_io_sel; // @[Benes.scala 98:28]
  wire [31:0] imm_switch_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_1_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_1_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_1_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_1_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_1_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_1_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_2_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_2_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_2_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_2_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_2_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_2_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_3_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_3_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_3_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_3_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_3_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_3_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_4_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_4_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_4_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_4_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_4_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_4_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_5_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_5_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_5_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_5_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_5_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_5_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_6_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_6_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_6_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_6_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_6_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_6_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_7_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_7_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_7_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_7_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_7_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_7_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_8_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_8_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_8_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_8_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_8_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_8_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_9_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_9_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_9_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_9_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_9_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_9_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_10_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_10_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_10_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_10_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_10_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_10_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_11_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_11_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_11_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_11_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_11_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_11_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_12_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_12_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_12_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_12_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_12_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_12_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_13_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_13_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_13_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_13_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_13_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_13_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_14_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_14_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_14_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_14_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_14_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_14_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_15_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_15_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_15_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_15_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_15_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_15_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_16_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_16_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_16_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_16_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_16_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_16_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_17_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_17_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_17_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_17_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_17_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_17_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_18_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_18_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_18_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_18_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_18_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_18_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_19_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_19_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_19_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_19_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_19_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_19_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_20_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_20_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_20_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_20_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_20_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_20_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_21_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_21_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_21_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_21_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_21_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_21_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_22_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_22_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_22_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_22_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_22_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_22_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_23_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_23_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_23_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_23_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_23_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_23_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_24_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_24_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_24_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_24_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_24_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_24_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_25_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_25_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_25_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_25_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_25_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_25_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_26_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_26_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_26_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_26_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_26_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_26_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_27_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_27_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_27_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_27_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_27_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_27_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_28_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_28_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_28_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_28_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_28_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_28_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_29_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_29_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_29_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_29_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_29_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_29_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_30_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_30_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_30_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_30_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_30_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_30_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_31_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_31_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_31_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_31_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_31_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_31_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_32_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_32_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_32_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_32_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_32_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_32_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_33_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_33_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_33_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_33_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_33_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_33_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_34_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_34_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_34_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_34_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_34_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_34_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_35_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_35_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_35_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_35_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_35_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_35_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_36_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_36_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_36_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_36_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_36_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_36_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_37_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_37_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_37_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_37_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_37_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_37_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_38_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_38_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_38_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_38_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_38_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_38_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_39_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_39_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_39_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_39_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_39_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_39_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_40_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_40_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_40_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_40_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_40_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_40_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_41_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_41_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_41_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_41_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_41_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_41_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_42_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_42_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_42_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_42_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_42_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_42_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_43_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_43_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_43_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_43_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_43_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_43_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_44_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_44_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_44_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_44_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_44_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_44_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_45_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_45_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_45_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_45_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_45_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_45_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_46_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_46_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_46_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_46_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_46_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_46_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_47_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_47_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_47_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_47_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_47_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_47_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_48_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_48_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_48_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_48_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_48_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_48_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_49_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_49_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_49_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_49_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_49_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_49_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_50_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_50_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_50_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_50_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_50_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_50_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_51_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_51_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_51_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_51_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_51_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_51_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_52_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_52_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_52_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_52_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_52_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_52_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_53_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_53_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_53_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_53_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_53_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_53_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_54_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_54_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_54_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_54_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_54_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_54_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_55_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_55_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_55_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_55_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_55_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_55_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_56_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_56_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_56_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_56_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_56_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_56_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_57_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_57_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_57_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_57_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_57_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_57_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_58_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_58_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_58_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_58_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_58_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_58_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_59_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_59_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_59_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_59_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_59_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_59_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_60_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_60_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_60_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_60_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_60_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_60_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_61_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_61_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_61_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_61_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_61_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_61_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_62_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_62_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_62_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_62_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_62_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_62_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_63_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_63_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_63_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_63_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_63_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_63_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_64_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_64_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_64_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_64_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_64_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_64_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_65_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_65_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_65_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_65_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_65_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_65_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_66_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_66_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_66_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_66_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_66_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_66_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_67_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_67_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_67_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_67_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_67_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_67_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_68_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_68_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_68_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_68_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_68_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_68_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_69_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_69_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_69_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_69_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_69_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_69_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_70_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_70_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_70_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_70_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_70_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_70_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_71_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_71_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_71_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_71_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_71_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_71_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_72_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_72_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_72_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_72_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_72_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_72_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_73_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_73_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_73_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_73_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_73_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_73_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_74_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_74_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_74_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_74_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_74_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_74_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_75_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_75_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_75_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_75_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_75_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_75_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_76_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_76_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_76_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_76_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_76_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_76_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_77_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_77_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_77_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_77_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_77_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_77_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_78_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_78_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_78_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_78_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_78_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_78_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_79_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_79_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_79_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_79_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_79_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_79_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_80_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_80_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_80_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_80_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_80_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_80_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_81_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_81_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_81_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_81_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_81_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_81_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_82_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_82_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_82_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_82_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_82_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_82_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_83_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_83_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_83_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_83_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_83_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_83_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_84_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_84_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_84_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_84_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_84_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_84_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_85_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_85_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_85_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_85_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_85_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_85_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_86_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_86_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_86_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_86_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_86_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_86_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_87_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_87_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_87_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_87_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_87_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_87_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_88_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_88_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_88_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_88_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_88_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_88_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_89_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_89_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_89_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_89_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_89_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_89_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_90_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_90_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_90_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_90_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_90_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_90_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_91_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_91_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_91_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_91_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_91_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_91_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_92_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_92_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_92_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_92_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_92_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_92_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_93_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_93_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_93_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_93_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_93_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_93_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_94_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_94_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_94_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_94_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_94_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_94_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_95_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_95_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_95_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_95_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_95_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_95_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_96_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_96_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_96_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_96_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_96_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_96_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_97_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_97_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_97_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_97_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_97_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_97_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_98_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_98_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_98_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_98_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_98_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_98_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_99_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_99_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_99_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_99_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_99_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_99_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_100_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_100_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_100_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_100_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_100_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_100_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_101_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_101_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_101_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_101_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_101_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_101_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_102_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_102_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_102_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_102_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_102_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_102_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_103_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_103_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_103_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_103_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_103_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_103_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_104_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_104_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_104_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_104_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_104_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_104_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_105_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_105_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_105_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_105_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_105_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_105_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_106_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_106_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_106_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_106_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_106_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_106_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_107_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_107_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_107_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_107_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_107_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_107_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_108_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_108_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_108_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_108_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_108_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_108_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_109_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_109_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_109_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_109_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_109_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_109_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_110_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_110_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_110_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_110_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_110_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_110_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_111_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_111_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_111_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_111_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_111_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_111_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_112_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_112_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_112_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_112_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_112_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_112_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_113_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_113_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_113_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_113_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_113_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_113_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_114_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_114_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_114_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_114_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_114_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_114_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_115_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_115_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_115_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_115_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_115_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_115_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_116_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_116_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_116_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_116_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_116_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_116_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_117_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_117_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_117_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_117_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_117_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_117_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_118_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_118_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_118_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_118_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_118_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_118_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_119_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_119_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_119_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_119_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_119_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_119_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_120_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_120_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_120_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_120_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_120_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_120_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_121_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_121_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_121_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_121_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_121_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_121_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_122_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_122_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_122_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_122_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_122_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_122_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_123_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_123_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_123_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_123_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_123_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_123_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_124_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_124_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_124_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_124_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_124_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_124_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_125_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_125_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_125_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_125_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_125_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_125_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_126_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_126_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_126_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_126_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_126_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_126_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_127_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_127_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_127_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_127_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_127_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_127_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_128_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_128_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_128_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_128_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_128_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_128_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_129_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_129_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_129_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_129_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_129_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_129_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_130_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_130_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_130_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_130_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_130_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_130_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_131_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_131_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_131_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_131_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_131_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_131_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_132_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_132_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_132_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_132_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_132_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_132_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_133_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_133_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_133_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_133_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_133_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_133_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_134_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_134_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_134_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_134_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_134_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_134_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_135_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_135_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_135_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_135_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_135_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_135_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_136_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_136_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_136_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_136_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_136_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_136_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_137_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_137_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_137_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_137_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_137_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_137_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_138_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_138_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_138_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_138_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_138_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_138_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_139_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_139_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_139_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_139_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_139_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_139_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_140_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_140_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_140_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_140_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_140_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_140_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_141_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_141_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_141_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_141_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_141_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_141_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_142_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_142_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_142_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_142_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_142_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_142_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_143_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_143_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_143_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_143_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_143_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_143_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_144_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_144_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_144_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_144_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_144_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_144_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_145_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_145_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_145_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_145_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_145_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_145_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_146_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_146_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_146_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_146_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_146_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_146_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_147_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_147_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_147_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_147_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_147_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_147_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_148_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_148_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_148_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_148_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_148_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_148_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_149_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_149_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_149_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_149_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_149_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_149_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_150_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_150_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_150_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_150_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_150_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_150_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_151_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_151_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_151_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_151_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_151_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_151_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_152_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_152_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_152_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_152_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_152_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_152_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_153_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_153_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_153_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_153_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_153_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_153_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_154_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_154_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_154_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_154_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_154_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_154_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_155_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_155_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_155_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_155_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_155_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_155_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_156_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_156_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_156_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_156_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_156_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_156_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_157_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_157_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_157_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_157_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_157_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_157_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_158_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_158_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_158_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_158_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_158_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_158_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_159_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_159_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_159_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_159_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_159_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_159_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_160_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_160_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_160_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_160_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_160_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_160_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_161_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_161_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_161_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_161_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_161_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_161_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_162_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_162_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_162_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_162_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_162_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_162_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_163_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_163_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_163_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_163_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_163_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_163_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_164_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_164_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_164_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_164_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_164_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_164_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_165_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_165_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_165_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_165_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_165_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_165_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_166_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_166_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_166_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_166_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_166_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_166_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_167_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_167_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_167_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_167_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_167_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_167_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_168_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_168_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_168_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_168_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_168_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_168_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_169_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_169_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_169_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_169_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_169_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_169_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_170_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_170_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_170_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_170_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_170_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_170_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_171_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_171_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_171_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_171_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_171_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_171_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_172_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_172_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_172_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_172_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_172_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_172_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_173_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_173_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_173_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_173_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_173_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_173_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_174_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_174_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_174_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_174_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_174_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_174_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_175_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_175_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_175_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_175_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_175_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_175_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_176_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_176_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_176_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_176_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_176_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_176_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_177_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_177_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_177_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_177_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_177_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_177_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_178_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_178_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_178_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_178_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_178_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_178_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_179_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_179_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_179_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_179_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_179_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_179_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_180_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_180_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_180_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_180_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_180_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_180_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_181_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_181_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_181_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_181_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_181_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_181_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_182_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_182_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_182_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_182_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_182_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_182_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_183_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_183_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_183_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_183_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_183_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_183_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_184_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_184_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_184_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_184_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_184_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_184_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_185_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_185_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_185_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_185_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_185_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_185_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_186_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_186_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_186_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_186_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_186_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_186_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_187_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_187_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_187_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_187_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_187_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_187_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_188_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_188_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_188_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_188_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_188_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_188_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_189_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_189_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_189_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_189_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_189_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_189_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_190_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_190_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_190_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_190_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_190_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_190_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_191_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_191_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_191_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_191_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_191_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_191_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_192_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_192_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_192_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_192_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_192_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_192_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_193_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_193_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_193_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_193_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_193_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_193_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_194_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_194_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_194_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_194_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_194_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_194_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_195_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_195_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_195_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_195_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_195_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_195_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_196_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_196_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_196_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_196_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_196_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_196_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_197_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_197_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_197_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_197_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_197_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_197_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_198_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_198_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_198_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_198_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_198_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_198_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_199_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_199_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_199_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_199_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_199_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_199_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_200_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_200_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_200_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_200_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_200_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_200_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_201_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_201_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_201_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_201_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_201_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_201_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_202_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_202_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_202_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_202_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_202_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_202_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_203_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_203_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_203_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_203_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_203_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_203_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_204_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_204_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_204_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_204_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_204_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_204_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_205_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_205_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_205_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_205_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_205_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_205_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_206_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_206_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_206_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_206_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_206_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_206_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_207_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_207_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_207_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_207_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_207_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_207_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_208_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_208_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_208_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_208_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_208_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_208_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_209_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_209_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_209_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_209_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_209_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_209_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_210_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_210_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_210_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_210_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_210_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_210_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_211_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_211_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_211_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_211_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_211_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_211_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_212_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_212_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_212_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_212_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_212_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_212_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_213_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_213_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_213_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_213_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_213_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_213_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_214_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_214_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_214_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_214_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_214_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_214_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_215_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_215_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_215_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_215_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_215_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_215_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_216_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_216_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_216_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_216_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_216_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_216_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_217_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_217_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_217_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_217_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_217_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_217_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_218_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_218_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_218_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_218_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_218_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_218_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_219_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_219_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_219_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_219_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_219_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_219_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_220_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_220_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_220_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_220_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_220_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_220_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_221_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_221_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_221_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_221_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_221_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_221_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_222_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_222_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_222_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_222_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_222_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_222_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_223_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_223_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_223_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_223_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_223_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_223_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_224_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_224_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_224_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_224_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_224_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_224_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_225_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_225_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_225_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_225_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_225_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_225_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_226_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_226_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_226_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_226_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_226_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_226_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_227_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_227_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_227_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_227_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_227_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_227_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_228_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_228_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_228_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_228_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_228_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_228_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_229_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_229_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_229_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_229_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_229_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_229_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_230_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_230_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_230_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_230_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_230_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_230_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_231_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_231_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_231_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_231_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_231_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_231_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_232_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_232_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_232_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_232_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_232_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_232_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_233_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_233_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_233_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_233_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_233_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_233_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_234_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_234_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_234_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_234_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_234_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_234_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_235_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_235_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_235_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_235_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_235_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_235_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_236_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_236_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_236_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_236_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_236_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_236_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_237_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_237_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_237_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_237_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_237_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_237_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_238_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_238_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_238_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_238_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_238_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_238_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_239_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_239_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_239_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_239_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_239_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_239_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_240_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_240_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_240_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_240_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_240_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_240_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_241_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_241_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_241_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_241_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_241_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_241_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_242_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_242_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_242_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_242_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_242_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_242_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_243_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_243_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_243_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_243_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_243_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_243_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_244_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_244_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_244_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_244_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_244_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_244_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_245_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_245_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_245_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_245_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_245_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_245_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_246_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_246_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_246_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_246_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_246_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_246_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_247_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_247_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_247_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_247_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_247_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_247_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_248_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_248_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_248_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_248_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_248_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_248_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_249_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_249_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_249_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_249_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_249_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_249_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_250_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_250_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_250_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_250_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_250_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_250_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_251_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_251_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_251_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_251_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_251_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_251_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_252_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_252_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_252_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_252_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_252_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_252_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_253_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_253_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_253_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_253_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_253_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_253_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_254_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_254_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_254_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_254_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_254_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_254_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_255_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_255_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_255_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_255_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_255_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_255_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_256_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_256_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_256_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_256_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_256_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_256_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_257_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_257_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_257_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_257_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_257_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_257_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_258_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_258_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_258_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_258_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_258_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_258_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_259_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_259_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_259_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_259_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_259_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_259_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_260_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_260_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_260_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_260_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_260_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_260_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_261_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_261_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_261_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_261_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_261_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_261_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_262_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_262_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_262_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_262_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_262_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_262_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_263_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_263_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_263_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_263_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_263_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_263_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_264_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_264_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_264_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_264_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_264_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_264_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_265_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_265_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_265_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_265_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_265_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_265_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_266_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_266_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_266_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_266_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_266_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_266_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_267_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_267_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_267_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_267_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_267_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_267_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_268_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_268_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_268_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_268_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_268_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_268_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_269_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_269_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_269_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_269_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_269_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_269_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_270_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_270_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_270_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_270_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_270_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_270_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_271_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_271_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_271_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_271_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_271_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_271_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_272_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_272_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_272_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_272_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_272_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_272_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_273_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_273_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_273_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_273_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_273_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_273_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_274_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_274_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_274_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_274_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_274_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_274_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_275_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_275_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_275_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_275_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_275_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_275_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_276_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_276_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_276_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_276_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_276_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_276_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_277_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_277_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_277_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_277_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_277_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_277_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_278_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_278_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_278_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_278_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_278_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_278_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_279_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_279_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_279_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_279_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_279_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_279_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_280_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_280_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_280_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_280_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_280_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_280_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_281_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_281_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_281_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_281_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_281_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_281_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_282_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_282_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_282_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_282_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_282_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_282_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_283_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_283_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_283_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_283_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_283_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_283_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_284_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_284_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_284_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_284_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_284_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_284_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_285_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_285_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_285_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_285_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_285_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_285_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_286_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_286_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_286_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_286_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_286_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_286_io_sel1; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_287_io_y; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_287_io_z; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_287_io_in0; // @[Benes.scala 108:30]
  wire [31:0] imm_switch_287_io_in1; // @[Benes.scala 108:30]
  wire  imm_switch_287_io_sel0; // @[Benes.scala 108:30]
  wire  imm_switch_287_io_sel1; // @[Benes.scala 108:30]
  reg [31:0] r_data_bus_ff_0; // @[Benes.scala 76:32]
  reg [31:0] r_data_bus_ff_1; // @[Benes.scala 76:32]
  reg [31:0] r_data_bus_ff_2; // @[Benes.scala 76:32]
  reg [31:0] r_data_bus_ff_3; // @[Benes.scala 76:32]
  reg [31:0] r_data_bus_ff_4; // @[Benes.scala 76:32]
  reg [31:0] r_data_bus_ff_5; // @[Benes.scala 76:32]
  reg [31:0] r_data_bus_ff_6; // @[Benes.scala 76:32]
  reg [31:0] r_data_bus_ff_7; // @[Benes.scala 76:32]
  reg [31:0] r_data_bus_ff_8; // @[Benes.scala 76:32]
  reg [31:0] r_data_bus_ff_9; // @[Benes.scala 76:32]
  reg [31:0] r_data_bus_ff_10; // @[Benes.scala 76:32]
  reg [31:0] r_data_bus_ff_11; // @[Benes.scala 76:32]
  reg [31:0] r_data_bus_ff_12; // @[Benes.scala 76:32]
  reg [31:0] r_data_bus_ff_13; // @[Benes.scala 76:32]
  reg [31:0] r_data_bus_ff_14; // @[Benes.scala 76:32]
  reg [31:0] r_data_bus_ff_15; // @[Benes.scala 76:32]
  reg [31:0] r_data_bus_ff_16; // @[Benes.scala 76:32]
  reg [31:0] r_data_bus_ff_17; // @[Benes.scala 76:32]
  reg [31:0] r_data_bus_ff_18; // @[Benes.scala 76:32]
  reg [31:0] r_data_bus_ff_19; // @[Benes.scala 76:32]
  reg [31:0] r_data_bus_ff_20; // @[Benes.scala 76:32]
  reg [31:0] r_data_bus_ff_21; // @[Benes.scala 76:32]
  reg [31:0] r_data_bus_ff_22; // @[Benes.scala 76:32]
  reg [31:0] r_data_bus_ff_23; // @[Benes.scala 76:32]
  reg [31:0] r_data_bus_ff_24; // @[Benes.scala 76:32]
  reg [31:0] r_data_bus_ff_25; // @[Benes.scala 76:32]
  reg [31:0] r_data_bus_ff_26; // @[Benes.scala 76:32]
  reg [31:0] r_data_bus_ff_27; // @[Benes.scala 76:32]
  reg [31:0] r_data_bus_ff_28; // @[Benes.scala 76:32]
  reg [31:0] r_data_bus_ff_29; // @[Benes.scala 76:32]
  reg [31:0] r_data_bus_ff_30; // @[Benes.scala 76:32]
  reg [31:0] r_data_bus_ff_31; // @[Benes.scala 76:32]
  reg  r_mux_bus_ff_0; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_1; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_2; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_3; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_4; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_5; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_6; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_7; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_8; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_9; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_10; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_11; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_12; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_13; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_14; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_15; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_16; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_17; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_18; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_19; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_20; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_21; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_22; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_23; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_24; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_25; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_26; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_27; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_28; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_29; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_30; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_31; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_32; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_33; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_34; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_35; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_36; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_37; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_38; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_39; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_40; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_41; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_42; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_43; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_44; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_45; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_46; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_47; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_48; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_49; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_50; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_51; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_52; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_53; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_54; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_55; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_56; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_57; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_58; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_59; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_60; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_61; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_62; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_63; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_64; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_65; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_66; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_67; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_68; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_69; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_70; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_71; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_72; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_73; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_74; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_75; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_76; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_77; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_78; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_79; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_80; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_81; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_82; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_83; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_84; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_85; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_86; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_87; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_88; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_89; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_90; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_91; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_92; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_93; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_94; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_95; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_96; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_97; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_98; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_99; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_100; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_101; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_102; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_103; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_104; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_105; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_106; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_107; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_108; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_109; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_110; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_111; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_112; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_113; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_114; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_115; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_116; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_117; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_118; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_119; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_120; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_121; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_122; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_123; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_124; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_125; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_126; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_127; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_128; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_129; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_130; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_131; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_132; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_133; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_134; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_135; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_136; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_137; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_138; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_139; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_140; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_141; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_142; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_143; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_144; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_145; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_146; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_147; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_148; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_149; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_150; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_151; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_152; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_153; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_154; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_155; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_156; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_157; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_158; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_159; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_160; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_161; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_162; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_163; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_164; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_165; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_166; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_167; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_168; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_169; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_170; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_171; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_172; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_173; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_174; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_175; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_176; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_177; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_178; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_179; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_180; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_181; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_182; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_183; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_184; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_185; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_186; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_187; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_188; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_189; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_190; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_191; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_192; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_193; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_194; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_195; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_196; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_197; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_198; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_199; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_200; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_201; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_202; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_203; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_204; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_205; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_206; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_207; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_208; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_209; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_210; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_211; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_212; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_213; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_214; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_215; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_216; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_217; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_218; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_219; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_220; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_221; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_222; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_223; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_224; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_225; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_226; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_227; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_228; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_229; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_230; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_231; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_232; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_233; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_234; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_235; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_236; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_237; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_238; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_239; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_240; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_241; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_242; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_243; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_244; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_245; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_246; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_247; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_248; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_249; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_250; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_251; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_252; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_253; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_254; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_255; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_256; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_257; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_258; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_259; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_260; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_261; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_262; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_263; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_264; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_265; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_266; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_267; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_268; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_269; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_270; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_271; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_272; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_273; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_274; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_275; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_276; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_277; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_278; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_279; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_280; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_281; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_282; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_283; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_284; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_285; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_286; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_287; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_288; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_289; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_290; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_291; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_292; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_293; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_294; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_295; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_296; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_297; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_298; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_299; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_300; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_301; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_302; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_303; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_304; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_305; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_306; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_307; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_308; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_309; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_310; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_311; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_312; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_313; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_314; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_315; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_316; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_317; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_318; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_319; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_320; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_321; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_322; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_323; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_324; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_325; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_326; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_327; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_328; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_329; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_330; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_331; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_332; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_333; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_334; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_335; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_336; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_337; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_338; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_339; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_340; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_341; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_342; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_343; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_344; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_345; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_346; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_347; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_348; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_349; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_350; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_351; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_352; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_353; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_354; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_355; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_356; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_357; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_358; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_359; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_360; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_361; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_362; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_363; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_364; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_365; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_366; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_367; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_368; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_369; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_370; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_371; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_372; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_373; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_374; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_375; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_376; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_377; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_378; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_379; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_380; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_381; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_382; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_383; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_384; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_385; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_386; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_387; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_388; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_389; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_390; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_391; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_392; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_393; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_394; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_395; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_396; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_397; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_398; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_399; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_400; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_401; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_402; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_403; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_404; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_405; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_406; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_407; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_408; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_409; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_410; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_411; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_412; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_413; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_414; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_415; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_416; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_417; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_418; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_419; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_420; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_421; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_422; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_423; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_424; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_425; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_426; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_427; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_428; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_429; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_430; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_431; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_432; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_433; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_434; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_435; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_436; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_437; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_438; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_439; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_440; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_441; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_442; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_443; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_444; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_445; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_446; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_447; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_448; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_449; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_450; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_451; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_452; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_453; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_454; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_455; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_456; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_457; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_458; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_459; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_460; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_461; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_462; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_463; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_464; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_465; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_466; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_467; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_468; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_469; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_470; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_471; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_472; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_473; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_474; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_475; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_476; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_477; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_478; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_479; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_480; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_481; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_482; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_483; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_484; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_485; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_486; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_487; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_488; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_489; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_490; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_491; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_492; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_493; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_494; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_495; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_496; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_497; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_498; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_499; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_500; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_501; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_502; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_503; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_504; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_505; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_506; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_507; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_508; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_509; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_510; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_511; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_512; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_513; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_514; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_515; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_516; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_517; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_518; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_519; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_520; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_521; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_522; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_523; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_524; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_525; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_526; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_527; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_528; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_529; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_530; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_531; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_532; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_533; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_534; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_535; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_536; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_537; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_538; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_539; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_540; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_541; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_542; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_543; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_544; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_545; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_546; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_547; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_548; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_549; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_550; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_551; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_552; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_553; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_554; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_555; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_556; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_557; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_558; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_559; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_560; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_561; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_562; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_563; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_564; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_565; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_566; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_567; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_568; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_569; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_570; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_571; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_572; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_573; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_574; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_575; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_576; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_577; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_578; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_579; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_580; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_581; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_582; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_583; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_584; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_585; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_586; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_587; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_588; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_589; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_590; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_591; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_592; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_593; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_594; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_595; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_596; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_597; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_598; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_599; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_600; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_601; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_602; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_603; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_604; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_605; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_606; // @[Benes.scala 77:32]
  reg  r_mux_bus_ff_607; // @[Benes.scala 77:32]
  wire [31:0] w_dist_bus_0 = out_switch_io_y; // @[Benes.scala 102:23 78:29]
  wire [31:0] w_dist_bus_1 = out_switch_1_io_y; // @[Benes.scala 102:23 78:29]
  wire [31:0] w_dist_bus_2 = out_switch_2_io_y; // @[Benes.scala 102:23 78:29]
  wire [31:0] w_dist_bus_3 = out_switch_3_io_y; // @[Benes.scala 102:23 78:29]
  wire [31:0] w_dist_bus_4 = out_switch_4_io_y; // @[Benes.scala 102:23 78:29]
  wire [31:0] w_dist_bus_5 = out_switch_5_io_y; // @[Benes.scala 102:23 78:29]
  wire [31:0] w_dist_bus_6 = out_switch_6_io_y; // @[Benes.scala 102:23 78:29]
  wire [31:0] w_dist_bus_7 = out_switch_7_io_y; // @[Benes.scala 102:23 78:29]
  wire [31:0] w_dist_bus_8 = out_switch_8_io_y; // @[Benes.scala 102:23 78:29]
  wire [31:0] w_dist_bus_9 = out_switch_9_io_y; // @[Benes.scala 102:23 78:29]
  wire [31:0] w_dist_bus_10 = out_switch_10_io_y; // @[Benes.scala 102:23 78:29]
  wire [31:0] w_dist_bus_11 = out_switch_11_io_y; // @[Benes.scala 102:23 78:29]
  wire [31:0] w_dist_bus_12 = out_switch_12_io_y; // @[Benes.scala 102:23 78:29]
  wire [31:0] w_dist_bus_13 = out_switch_13_io_y; // @[Benes.scala 102:23 78:29]
  wire [31:0] w_dist_bus_14 = out_switch_14_io_y; // @[Benes.scala 102:23 78:29]
  wire [31:0] w_dist_bus_15 = out_switch_15_io_y; // @[Benes.scala 102:23 78:29]
  wire [31:0] w_dist_bus_16 = out_switch_16_io_y; // @[Benes.scala 102:23 78:29]
  wire [31:0] w_dist_bus_17 = out_switch_17_io_y; // @[Benes.scala 102:23 78:29]
  wire [31:0] w_dist_bus_18 = out_switch_18_io_y; // @[Benes.scala 102:23 78:29]
  wire [31:0] w_dist_bus_19 = out_switch_19_io_y; // @[Benes.scala 102:23 78:29]
  wire [31:0] w_dist_bus_20 = out_switch_20_io_y; // @[Benes.scala 102:23 78:29]
  wire [31:0] w_dist_bus_21 = out_switch_21_io_y; // @[Benes.scala 102:23 78:29]
  wire [31:0] w_dist_bus_22 = out_switch_22_io_y; // @[Benes.scala 102:23 78:29]
  wire [31:0] w_dist_bus_23 = out_switch_23_io_y; // @[Benes.scala 102:23 78:29]
  wire [31:0] w_dist_bus_24 = out_switch_24_io_y; // @[Benes.scala 102:23 78:29]
  wire [31:0] w_dist_bus_25 = out_switch_25_io_y; // @[Benes.scala 102:23 78:29]
  wire [31:0] w_dist_bus_26 = out_switch_26_io_y; // @[Benes.scala 102:23 78:29]
  wire [31:0] w_dist_bus_27 = out_switch_27_io_y; // @[Benes.scala 102:23 78:29]
  wire [31:0] w_dist_bus_28 = out_switch_28_io_y; // @[Benes.scala 102:23 78:29]
  wire [31:0] w_dist_bus_29 = out_switch_29_io_y; // @[Benes.scala 102:23 78:29]
  wire [31:0] w_dist_bus_30 = out_switch_30_io_y; // @[Benes.scala 102:23 78:29]
  wire [31:0] w_dist_bus_31 = out_switch_31_io_y; // @[Benes.scala 102:23 78:29]
  wire [31:0] w_internal_0 = in_switch_io_y; // @[Benes.scala 79:29 91:43]
  wire [31:0] w_internal_1 = in_switch_io_z; // @[Benes.scala 79:29 92:43]
  wire [31:0] w_internal_2 = imm_switch_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_3 = imm_switch_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_4 = imm_switch_1_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_5 = imm_switch_1_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_6 = imm_switch_2_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_7 = imm_switch_2_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_8 = imm_switch_3_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_9 = imm_switch_3_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_10 = imm_switch_4_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_11 = imm_switch_4_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_12 = imm_switch_5_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_13 = imm_switch_5_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_14 = imm_switch_6_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_15 = imm_switch_6_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_16 = imm_switch_7_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_17 = imm_switch_7_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_18 = imm_switch_8_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_19 = imm_switch_8_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_20 = in_switch_1_io_y; // @[Benes.scala 79:29 91:43]
  wire [31:0] w_internal_21 = in_switch_1_io_z; // @[Benes.scala 79:29 92:43]
  wire [31:0] w_internal_22 = imm_switch_9_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_23 = imm_switch_9_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_24 = imm_switch_10_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_25 = imm_switch_10_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_26 = imm_switch_11_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_27 = imm_switch_11_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_28 = imm_switch_12_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_29 = imm_switch_12_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_30 = imm_switch_13_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_31 = imm_switch_13_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_32 = imm_switch_14_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_33 = imm_switch_14_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_34 = imm_switch_15_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_35 = imm_switch_15_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_36 = imm_switch_16_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_37 = imm_switch_16_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_38 = imm_switch_17_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_39 = imm_switch_17_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_40 = in_switch_2_io_y; // @[Benes.scala 79:29 91:43]
  wire [31:0] w_internal_41 = in_switch_2_io_z; // @[Benes.scala 79:29 92:43]
  wire [31:0] w_internal_42 = imm_switch_18_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_43 = imm_switch_18_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_44 = imm_switch_19_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_45 = imm_switch_19_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_46 = imm_switch_20_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_47 = imm_switch_20_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_48 = imm_switch_21_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_49 = imm_switch_21_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_50 = imm_switch_22_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_51 = imm_switch_22_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_52 = imm_switch_23_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_53 = imm_switch_23_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_54 = imm_switch_24_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_55 = imm_switch_24_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_56 = imm_switch_25_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_57 = imm_switch_25_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_58 = imm_switch_26_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_59 = imm_switch_26_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_60 = in_switch_3_io_y; // @[Benes.scala 79:29 91:43]
  wire [31:0] w_internal_61 = in_switch_3_io_z; // @[Benes.scala 79:29 92:43]
  wire [31:0] w_internal_62 = imm_switch_27_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_63 = imm_switch_27_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_64 = imm_switch_28_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_65 = imm_switch_28_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_66 = imm_switch_29_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_67 = imm_switch_29_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_68 = imm_switch_30_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_69 = imm_switch_30_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_70 = imm_switch_31_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_71 = imm_switch_31_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_72 = imm_switch_32_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_73 = imm_switch_32_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_74 = imm_switch_33_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_75 = imm_switch_33_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_76 = imm_switch_34_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_77 = imm_switch_34_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_78 = imm_switch_35_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_79 = imm_switch_35_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_80 = in_switch_4_io_y; // @[Benes.scala 79:29 91:43]
  wire [31:0] w_internal_81 = in_switch_4_io_z; // @[Benes.scala 79:29 92:43]
  wire [31:0] w_internal_82 = imm_switch_36_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_83 = imm_switch_36_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_84 = imm_switch_37_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_85 = imm_switch_37_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_86 = imm_switch_38_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_87 = imm_switch_38_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_88 = imm_switch_39_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_89 = imm_switch_39_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_90 = imm_switch_40_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_91 = imm_switch_40_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_92 = imm_switch_41_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_93 = imm_switch_41_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_94 = imm_switch_42_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_95 = imm_switch_42_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_96 = imm_switch_43_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_97 = imm_switch_43_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_98 = imm_switch_44_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_99 = imm_switch_44_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_100 = in_switch_5_io_y; // @[Benes.scala 79:29 91:43]
  wire [31:0] w_internal_101 = in_switch_5_io_z; // @[Benes.scala 79:29 92:43]
  wire [31:0] w_internal_102 = imm_switch_45_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_103 = imm_switch_45_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_104 = imm_switch_46_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_105 = imm_switch_46_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_106 = imm_switch_47_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_107 = imm_switch_47_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_108 = imm_switch_48_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_109 = imm_switch_48_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_110 = imm_switch_49_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_111 = imm_switch_49_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_112 = imm_switch_50_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_113 = imm_switch_50_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_114 = imm_switch_51_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_115 = imm_switch_51_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_116 = imm_switch_52_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_117 = imm_switch_52_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_118 = imm_switch_53_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_119 = imm_switch_53_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_120 = in_switch_6_io_y; // @[Benes.scala 79:29 91:43]
  wire [31:0] w_internal_121 = in_switch_6_io_z; // @[Benes.scala 79:29 92:43]
  wire [31:0] w_internal_122 = imm_switch_54_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_123 = imm_switch_54_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_124 = imm_switch_55_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_125 = imm_switch_55_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_126 = imm_switch_56_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_127 = imm_switch_56_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_128 = imm_switch_57_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_129 = imm_switch_57_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_130 = imm_switch_58_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_131 = imm_switch_58_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_132 = imm_switch_59_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_133 = imm_switch_59_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_134 = imm_switch_60_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_135 = imm_switch_60_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_136 = imm_switch_61_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_137 = imm_switch_61_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_138 = imm_switch_62_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_139 = imm_switch_62_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_140 = in_switch_7_io_y; // @[Benes.scala 79:29 91:43]
  wire [31:0] w_internal_141 = in_switch_7_io_z; // @[Benes.scala 79:29 92:43]
  wire [31:0] w_internal_142 = imm_switch_63_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_143 = imm_switch_63_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_144 = imm_switch_64_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_145 = imm_switch_64_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_146 = imm_switch_65_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_147 = imm_switch_65_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_148 = imm_switch_66_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_149 = imm_switch_66_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_150 = imm_switch_67_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_151 = imm_switch_67_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_152 = imm_switch_68_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_153 = imm_switch_68_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_154 = imm_switch_69_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_155 = imm_switch_69_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_156 = imm_switch_70_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_157 = imm_switch_70_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_158 = imm_switch_71_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_159 = imm_switch_71_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_160 = in_switch_8_io_y; // @[Benes.scala 79:29 91:43]
  wire [31:0] w_internal_161 = in_switch_8_io_z; // @[Benes.scala 79:29 92:43]
  wire [31:0] w_internal_162 = imm_switch_72_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_163 = imm_switch_72_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_164 = imm_switch_73_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_165 = imm_switch_73_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_166 = imm_switch_74_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_167 = imm_switch_74_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_168 = imm_switch_75_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_169 = imm_switch_75_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_170 = imm_switch_76_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_171 = imm_switch_76_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_172 = imm_switch_77_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_173 = imm_switch_77_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_174 = imm_switch_78_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_175 = imm_switch_78_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_176 = imm_switch_79_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_177 = imm_switch_79_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_178 = imm_switch_80_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_179 = imm_switch_80_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_180 = in_switch_9_io_y; // @[Benes.scala 79:29 91:43]
  wire [31:0] w_internal_181 = in_switch_9_io_z; // @[Benes.scala 79:29 92:43]
  wire [31:0] w_internal_182 = imm_switch_81_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_183 = imm_switch_81_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_184 = imm_switch_82_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_185 = imm_switch_82_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_186 = imm_switch_83_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_187 = imm_switch_83_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_188 = imm_switch_84_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_189 = imm_switch_84_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_190 = imm_switch_85_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_191 = imm_switch_85_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_192 = imm_switch_86_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_193 = imm_switch_86_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_194 = imm_switch_87_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_195 = imm_switch_87_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_196 = imm_switch_88_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_197 = imm_switch_88_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_198 = imm_switch_89_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_199 = imm_switch_89_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_200 = in_switch_10_io_y; // @[Benes.scala 79:29 91:43]
  wire [31:0] w_internal_201 = in_switch_10_io_z; // @[Benes.scala 79:29 92:43]
  wire [31:0] w_internal_202 = imm_switch_90_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_203 = imm_switch_90_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_204 = imm_switch_91_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_205 = imm_switch_91_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_206 = imm_switch_92_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_207 = imm_switch_92_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_208 = imm_switch_93_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_209 = imm_switch_93_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_210 = imm_switch_94_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_211 = imm_switch_94_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_212 = imm_switch_95_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_213 = imm_switch_95_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_214 = imm_switch_96_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_215 = imm_switch_96_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_216 = imm_switch_97_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_217 = imm_switch_97_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_218 = imm_switch_98_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_219 = imm_switch_98_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_220 = in_switch_11_io_y; // @[Benes.scala 79:29 91:43]
  wire [31:0] w_internal_221 = in_switch_11_io_z; // @[Benes.scala 79:29 92:43]
  wire [31:0] w_internal_222 = imm_switch_99_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_223 = imm_switch_99_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_224 = imm_switch_100_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_225 = imm_switch_100_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_226 = imm_switch_101_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_227 = imm_switch_101_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_228 = imm_switch_102_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_229 = imm_switch_102_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_230 = imm_switch_103_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_231 = imm_switch_103_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_232 = imm_switch_104_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_233 = imm_switch_104_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_234 = imm_switch_105_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_235 = imm_switch_105_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_236 = imm_switch_106_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_237 = imm_switch_106_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_238 = imm_switch_107_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_239 = imm_switch_107_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_240 = in_switch_12_io_y; // @[Benes.scala 79:29 91:43]
  wire [31:0] w_internal_241 = in_switch_12_io_z; // @[Benes.scala 79:29 92:43]
  wire [31:0] w_internal_242 = imm_switch_108_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_243 = imm_switch_108_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_244 = imm_switch_109_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_245 = imm_switch_109_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_246 = imm_switch_110_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_247 = imm_switch_110_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_248 = imm_switch_111_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_249 = imm_switch_111_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_250 = imm_switch_112_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_251 = imm_switch_112_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_252 = imm_switch_113_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_253 = imm_switch_113_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_254 = imm_switch_114_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_255 = imm_switch_114_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_256 = imm_switch_115_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_257 = imm_switch_115_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_258 = imm_switch_116_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_259 = imm_switch_116_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_260 = in_switch_13_io_y; // @[Benes.scala 79:29 91:43]
  wire [31:0] w_internal_261 = in_switch_13_io_z; // @[Benes.scala 79:29 92:43]
  wire [31:0] w_internal_262 = imm_switch_117_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_263 = imm_switch_117_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_264 = imm_switch_118_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_265 = imm_switch_118_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_266 = imm_switch_119_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_267 = imm_switch_119_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_268 = imm_switch_120_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_269 = imm_switch_120_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_270 = imm_switch_121_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_271 = imm_switch_121_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_272 = imm_switch_122_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_273 = imm_switch_122_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_274 = imm_switch_123_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_275 = imm_switch_123_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_276 = imm_switch_124_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_277 = imm_switch_124_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_278 = imm_switch_125_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_279 = imm_switch_125_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_280 = in_switch_14_io_y; // @[Benes.scala 79:29 91:43]
  wire [31:0] w_internal_281 = in_switch_14_io_z; // @[Benes.scala 79:29 92:43]
  wire [31:0] w_internal_282 = imm_switch_126_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_283 = imm_switch_126_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_284 = imm_switch_127_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_285 = imm_switch_127_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_286 = imm_switch_128_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_287 = imm_switch_128_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_288 = imm_switch_129_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_289 = imm_switch_129_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_290 = imm_switch_130_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_291 = imm_switch_130_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_292 = imm_switch_131_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_293 = imm_switch_131_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_294 = imm_switch_132_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_295 = imm_switch_132_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_296 = imm_switch_133_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_297 = imm_switch_133_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_298 = imm_switch_134_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_299 = imm_switch_134_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_300 = in_switch_15_io_y; // @[Benes.scala 79:29 91:43]
  wire [31:0] w_internal_301 = in_switch_15_io_z; // @[Benes.scala 79:29 92:43]
  wire [31:0] w_internal_302 = imm_switch_135_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_303 = imm_switch_135_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_304 = imm_switch_136_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_305 = imm_switch_136_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_306 = imm_switch_137_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_307 = imm_switch_137_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_308 = imm_switch_138_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_309 = imm_switch_138_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_310 = imm_switch_139_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_311 = imm_switch_139_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_312 = imm_switch_140_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_313 = imm_switch_140_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_314 = imm_switch_141_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_315 = imm_switch_141_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_316 = imm_switch_142_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_317 = imm_switch_142_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_318 = imm_switch_143_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_319 = imm_switch_143_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_320 = in_switch_16_io_y; // @[Benes.scala 79:29 91:43]
  wire [31:0] w_internal_321 = in_switch_16_io_z; // @[Benes.scala 79:29 92:43]
  wire [31:0] w_internal_322 = imm_switch_144_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_323 = imm_switch_144_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_324 = imm_switch_145_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_325 = imm_switch_145_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_326 = imm_switch_146_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_327 = imm_switch_146_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_328 = imm_switch_147_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_329 = imm_switch_147_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_330 = imm_switch_148_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_331 = imm_switch_148_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_332 = imm_switch_149_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_333 = imm_switch_149_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_334 = imm_switch_150_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_335 = imm_switch_150_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_336 = imm_switch_151_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_337 = imm_switch_151_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_338 = imm_switch_152_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_339 = imm_switch_152_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_340 = in_switch_17_io_y; // @[Benes.scala 79:29 91:43]
  wire [31:0] w_internal_341 = in_switch_17_io_z; // @[Benes.scala 79:29 92:43]
  wire [31:0] w_internal_342 = imm_switch_153_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_343 = imm_switch_153_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_344 = imm_switch_154_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_345 = imm_switch_154_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_346 = imm_switch_155_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_347 = imm_switch_155_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_348 = imm_switch_156_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_349 = imm_switch_156_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_350 = imm_switch_157_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_351 = imm_switch_157_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_352 = imm_switch_158_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_353 = imm_switch_158_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_354 = imm_switch_159_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_355 = imm_switch_159_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_356 = imm_switch_160_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_357 = imm_switch_160_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_358 = imm_switch_161_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_359 = imm_switch_161_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_360 = in_switch_18_io_y; // @[Benes.scala 79:29 91:43]
  wire [31:0] w_internal_361 = in_switch_18_io_z; // @[Benes.scala 79:29 92:43]
  wire [31:0] w_internal_362 = imm_switch_162_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_363 = imm_switch_162_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_364 = imm_switch_163_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_365 = imm_switch_163_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_366 = imm_switch_164_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_367 = imm_switch_164_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_368 = imm_switch_165_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_369 = imm_switch_165_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_370 = imm_switch_166_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_371 = imm_switch_166_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_372 = imm_switch_167_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_373 = imm_switch_167_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_374 = imm_switch_168_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_375 = imm_switch_168_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_376 = imm_switch_169_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_377 = imm_switch_169_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_378 = imm_switch_170_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_379 = imm_switch_170_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_380 = in_switch_19_io_y; // @[Benes.scala 79:29 91:43]
  wire [31:0] w_internal_381 = in_switch_19_io_z; // @[Benes.scala 79:29 92:43]
  wire [31:0] w_internal_382 = imm_switch_171_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_383 = imm_switch_171_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_384 = imm_switch_172_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_385 = imm_switch_172_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_386 = imm_switch_173_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_387 = imm_switch_173_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_388 = imm_switch_174_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_389 = imm_switch_174_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_390 = imm_switch_175_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_391 = imm_switch_175_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_392 = imm_switch_176_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_393 = imm_switch_176_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_394 = imm_switch_177_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_395 = imm_switch_177_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_396 = imm_switch_178_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_397 = imm_switch_178_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_398 = imm_switch_179_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_399 = imm_switch_179_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_400 = in_switch_20_io_y; // @[Benes.scala 79:29 91:43]
  wire [31:0] w_internal_401 = in_switch_20_io_z; // @[Benes.scala 79:29 92:43]
  wire [31:0] w_internal_402 = imm_switch_180_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_403 = imm_switch_180_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_404 = imm_switch_181_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_405 = imm_switch_181_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_406 = imm_switch_182_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_407 = imm_switch_182_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_408 = imm_switch_183_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_409 = imm_switch_183_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_410 = imm_switch_184_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_411 = imm_switch_184_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_412 = imm_switch_185_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_413 = imm_switch_185_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_414 = imm_switch_186_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_415 = imm_switch_186_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_416 = imm_switch_187_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_417 = imm_switch_187_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_418 = imm_switch_188_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_419 = imm_switch_188_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_420 = in_switch_21_io_y; // @[Benes.scala 79:29 91:43]
  wire [31:0] w_internal_421 = in_switch_21_io_z; // @[Benes.scala 79:29 92:43]
  wire [31:0] w_internal_422 = imm_switch_189_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_423 = imm_switch_189_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_424 = imm_switch_190_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_425 = imm_switch_190_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_426 = imm_switch_191_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_427 = imm_switch_191_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_428 = imm_switch_192_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_429 = imm_switch_192_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_430 = imm_switch_193_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_431 = imm_switch_193_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_432 = imm_switch_194_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_433 = imm_switch_194_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_434 = imm_switch_195_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_435 = imm_switch_195_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_436 = imm_switch_196_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_437 = imm_switch_196_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_438 = imm_switch_197_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_439 = imm_switch_197_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_440 = in_switch_22_io_y; // @[Benes.scala 79:29 91:43]
  wire [31:0] w_internal_441 = in_switch_22_io_z; // @[Benes.scala 79:29 92:43]
  wire [31:0] w_internal_442 = imm_switch_198_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_443 = imm_switch_198_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_444 = imm_switch_199_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_445 = imm_switch_199_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_446 = imm_switch_200_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_447 = imm_switch_200_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_448 = imm_switch_201_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_449 = imm_switch_201_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_450 = imm_switch_202_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_451 = imm_switch_202_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_452 = imm_switch_203_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_453 = imm_switch_203_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_454 = imm_switch_204_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_455 = imm_switch_204_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_456 = imm_switch_205_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_457 = imm_switch_205_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_458 = imm_switch_206_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_459 = imm_switch_206_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_460 = in_switch_23_io_y; // @[Benes.scala 79:29 91:43]
  wire [31:0] w_internal_461 = in_switch_23_io_z; // @[Benes.scala 79:29 92:43]
  wire [31:0] w_internal_462 = imm_switch_207_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_463 = imm_switch_207_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_464 = imm_switch_208_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_465 = imm_switch_208_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_466 = imm_switch_209_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_467 = imm_switch_209_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_468 = imm_switch_210_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_469 = imm_switch_210_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_470 = imm_switch_211_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_471 = imm_switch_211_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_472 = imm_switch_212_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_473 = imm_switch_212_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_474 = imm_switch_213_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_475 = imm_switch_213_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_476 = imm_switch_214_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_477 = imm_switch_214_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_478 = imm_switch_215_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_479 = imm_switch_215_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_480 = in_switch_24_io_y; // @[Benes.scala 79:29 91:43]
  wire [31:0] w_internal_481 = in_switch_24_io_z; // @[Benes.scala 79:29 92:43]
  wire [31:0] w_internal_482 = imm_switch_216_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_483 = imm_switch_216_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_484 = imm_switch_217_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_485 = imm_switch_217_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_486 = imm_switch_218_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_487 = imm_switch_218_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_488 = imm_switch_219_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_489 = imm_switch_219_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_490 = imm_switch_220_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_491 = imm_switch_220_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_492 = imm_switch_221_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_493 = imm_switch_221_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_494 = imm_switch_222_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_495 = imm_switch_222_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_496 = imm_switch_223_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_497 = imm_switch_223_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_498 = imm_switch_224_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_499 = imm_switch_224_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_500 = in_switch_25_io_y; // @[Benes.scala 79:29 91:43]
  wire [31:0] w_internal_501 = in_switch_25_io_z; // @[Benes.scala 79:29 92:43]
  wire [31:0] w_internal_502 = imm_switch_225_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_503 = imm_switch_225_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_504 = imm_switch_226_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_505 = imm_switch_226_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_506 = imm_switch_227_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_507 = imm_switch_227_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_508 = imm_switch_228_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_509 = imm_switch_228_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_510 = imm_switch_229_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_511 = imm_switch_229_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_512 = imm_switch_230_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_513 = imm_switch_230_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_514 = imm_switch_231_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_515 = imm_switch_231_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_516 = imm_switch_232_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_517 = imm_switch_232_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_518 = imm_switch_233_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_519 = imm_switch_233_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_520 = in_switch_26_io_y; // @[Benes.scala 79:29 91:43]
  wire [31:0] w_internal_521 = in_switch_26_io_z; // @[Benes.scala 79:29 92:43]
  wire [31:0] w_internal_522 = imm_switch_234_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_523 = imm_switch_234_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_524 = imm_switch_235_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_525 = imm_switch_235_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_526 = imm_switch_236_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_527 = imm_switch_236_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_528 = imm_switch_237_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_529 = imm_switch_237_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_530 = imm_switch_238_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_531 = imm_switch_238_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_532 = imm_switch_239_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_533 = imm_switch_239_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_534 = imm_switch_240_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_535 = imm_switch_240_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_536 = imm_switch_241_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_537 = imm_switch_241_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_538 = imm_switch_242_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_539 = imm_switch_242_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_540 = in_switch_27_io_y; // @[Benes.scala 79:29 91:43]
  wire [31:0] w_internal_541 = in_switch_27_io_z; // @[Benes.scala 79:29 92:43]
  wire [31:0] w_internal_542 = imm_switch_243_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_543 = imm_switch_243_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_544 = imm_switch_244_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_545 = imm_switch_244_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_546 = imm_switch_245_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_547 = imm_switch_245_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_548 = imm_switch_246_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_549 = imm_switch_246_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_550 = imm_switch_247_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_551 = imm_switch_247_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_552 = imm_switch_248_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_553 = imm_switch_248_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_554 = imm_switch_249_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_555 = imm_switch_249_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_556 = imm_switch_250_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_557 = imm_switch_250_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_558 = imm_switch_251_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_559 = imm_switch_251_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_560 = in_switch_28_io_y; // @[Benes.scala 79:29 91:43]
  wire [31:0] w_internal_561 = in_switch_28_io_z; // @[Benes.scala 79:29 92:43]
  wire [31:0] w_internal_562 = imm_switch_252_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_563 = imm_switch_252_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_564 = imm_switch_253_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_565 = imm_switch_253_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_566 = imm_switch_254_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_567 = imm_switch_254_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_568 = imm_switch_255_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_569 = imm_switch_255_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_570 = imm_switch_256_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_571 = imm_switch_256_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_572 = imm_switch_257_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_573 = imm_switch_257_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_574 = imm_switch_258_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_575 = imm_switch_258_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_576 = imm_switch_259_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_577 = imm_switch_259_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_578 = imm_switch_260_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_579 = imm_switch_260_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_580 = in_switch_29_io_y; // @[Benes.scala 79:29 91:43]
  wire [31:0] w_internal_581 = in_switch_29_io_z; // @[Benes.scala 79:29 92:43]
  wire [31:0] w_internal_582 = imm_switch_261_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_583 = imm_switch_261_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_584 = imm_switch_262_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_585 = imm_switch_262_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_586 = imm_switch_263_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_587 = imm_switch_263_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_588 = imm_switch_264_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_589 = imm_switch_264_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_590 = imm_switch_265_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_591 = imm_switch_265_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_592 = imm_switch_266_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_593 = imm_switch_266_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_594 = imm_switch_267_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_595 = imm_switch_267_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_596 = imm_switch_268_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_597 = imm_switch_268_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_598 = imm_switch_269_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_599 = imm_switch_269_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_600 = in_switch_30_io_y; // @[Benes.scala 79:29 91:43]
  wire [31:0] w_internal_601 = in_switch_30_io_z; // @[Benes.scala 79:29 92:43]
  wire [31:0] w_internal_602 = imm_switch_270_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_603 = imm_switch_270_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_604 = imm_switch_271_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_605 = imm_switch_271_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_606 = imm_switch_272_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_607 = imm_switch_272_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_608 = imm_switch_273_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_609 = imm_switch_273_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_610 = imm_switch_274_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_611 = imm_switch_274_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_612 = imm_switch_275_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_613 = imm_switch_275_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_614 = imm_switch_276_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_615 = imm_switch_276_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_616 = imm_switch_277_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_617 = imm_switch_277_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_618 = imm_switch_278_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_619 = imm_switch_278_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_620 = in_switch_31_io_y; // @[Benes.scala 79:29 91:43]
  wire [31:0] w_internal_621 = in_switch_31_io_z; // @[Benes.scala 79:29 92:43]
  wire [31:0] w_internal_622 = imm_switch_279_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_623 = imm_switch_279_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_624 = imm_switch_280_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_625 = imm_switch_280_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_626 = imm_switch_281_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_627 = imm_switch_281_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_628 = imm_switch_282_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_629 = imm_switch_282_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_630 = imm_switch_283_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_631 = imm_switch_283_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_632 = imm_switch_284_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_633 = imm_switch_284_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_634 = imm_switch_285_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_635 = imm_switch_285_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_636 = imm_switch_286_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_637 = imm_switch_286_io_z; // @[Benes.scala 79:29 126:53]
  wire [31:0] w_internal_638 = imm_switch_287_io_y; // @[Benes.scala 79:29 125:53]
  wire [31:0] w_internal_639 = imm_switch_287_io_z; // @[Benes.scala 79:29 126:53]
  InputSwitch in_switch ( // @[Benes.scala 89:27]
    .io_y(in_switch_io_y),
    .io_z(in_switch_io_z),
    .io_in(in_switch_io_in)
  );
  InputSwitch in_switch_1 ( // @[Benes.scala 89:27]
    .io_y(in_switch_1_io_y),
    .io_z(in_switch_1_io_z),
    .io_in(in_switch_1_io_in)
  );
  InputSwitch in_switch_2 ( // @[Benes.scala 89:27]
    .io_y(in_switch_2_io_y),
    .io_z(in_switch_2_io_z),
    .io_in(in_switch_2_io_in)
  );
  InputSwitch in_switch_3 ( // @[Benes.scala 89:27]
    .io_y(in_switch_3_io_y),
    .io_z(in_switch_3_io_z),
    .io_in(in_switch_3_io_in)
  );
  InputSwitch in_switch_4 ( // @[Benes.scala 89:27]
    .io_y(in_switch_4_io_y),
    .io_z(in_switch_4_io_z),
    .io_in(in_switch_4_io_in)
  );
  InputSwitch in_switch_5 ( // @[Benes.scala 89:27]
    .io_y(in_switch_5_io_y),
    .io_z(in_switch_5_io_z),
    .io_in(in_switch_5_io_in)
  );
  InputSwitch in_switch_6 ( // @[Benes.scala 89:27]
    .io_y(in_switch_6_io_y),
    .io_z(in_switch_6_io_z),
    .io_in(in_switch_6_io_in)
  );
  InputSwitch in_switch_7 ( // @[Benes.scala 89:27]
    .io_y(in_switch_7_io_y),
    .io_z(in_switch_7_io_z),
    .io_in(in_switch_7_io_in)
  );
  InputSwitch in_switch_8 ( // @[Benes.scala 89:27]
    .io_y(in_switch_8_io_y),
    .io_z(in_switch_8_io_z),
    .io_in(in_switch_8_io_in)
  );
  InputSwitch in_switch_9 ( // @[Benes.scala 89:27]
    .io_y(in_switch_9_io_y),
    .io_z(in_switch_9_io_z),
    .io_in(in_switch_9_io_in)
  );
  InputSwitch in_switch_10 ( // @[Benes.scala 89:27]
    .io_y(in_switch_10_io_y),
    .io_z(in_switch_10_io_z),
    .io_in(in_switch_10_io_in)
  );
  InputSwitch in_switch_11 ( // @[Benes.scala 89:27]
    .io_y(in_switch_11_io_y),
    .io_z(in_switch_11_io_z),
    .io_in(in_switch_11_io_in)
  );
  InputSwitch in_switch_12 ( // @[Benes.scala 89:27]
    .io_y(in_switch_12_io_y),
    .io_z(in_switch_12_io_z),
    .io_in(in_switch_12_io_in)
  );
  InputSwitch in_switch_13 ( // @[Benes.scala 89:27]
    .io_y(in_switch_13_io_y),
    .io_z(in_switch_13_io_z),
    .io_in(in_switch_13_io_in)
  );
  InputSwitch in_switch_14 ( // @[Benes.scala 89:27]
    .io_y(in_switch_14_io_y),
    .io_z(in_switch_14_io_z),
    .io_in(in_switch_14_io_in)
  );
  InputSwitch in_switch_15 ( // @[Benes.scala 89:27]
    .io_y(in_switch_15_io_y),
    .io_z(in_switch_15_io_z),
    .io_in(in_switch_15_io_in)
  );
  InputSwitch in_switch_16 ( // @[Benes.scala 89:27]
    .io_y(in_switch_16_io_y),
    .io_z(in_switch_16_io_z),
    .io_in(in_switch_16_io_in)
  );
  InputSwitch in_switch_17 ( // @[Benes.scala 89:27]
    .io_y(in_switch_17_io_y),
    .io_z(in_switch_17_io_z),
    .io_in(in_switch_17_io_in)
  );
  InputSwitch in_switch_18 ( // @[Benes.scala 89:27]
    .io_y(in_switch_18_io_y),
    .io_z(in_switch_18_io_z),
    .io_in(in_switch_18_io_in)
  );
  InputSwitch in_switch_19 ( // @[Benes.scala 89:27]
    .io_y(in_switch_19_io_y),
    .io_z(in_switch_19_io_z),
    .io_in(in_switch_19_io_in)
  );
  InputSwitch in_switch_20 ( // @[Benes.scala 89:27]
    .io_y(in_switch_20_io_y),
    .io_z(in_switch_20_io_z),
    .io_in(in_switch_20_io_in)
  );
  InputSwitch in_switch_21 ( // @[Benes.scala 89:27]
    .io_y(in_switch_21_io_y),
    .io_z(in_switch_21_io_z),
    .io_in(in_switch_21_io_in)
  );
  InputSwitch in_switch_22 ( // @[Benes.scala 89:27]
    .io_y(in_switch_22_io_y),
    .io_z(in_switch_22_io_z),
    .io_in(in_switch_22_io_in)
  );
  InputSwitch in_switch_23 ( // @[Benes.scala 89:27]
    .io_y(in_switch_23_io_y),
    .io_z(in_switch_23_io_z),
    .io_in(in_switch_23_io_in)
  );
  InputSwitch in_switch_24 ( // @[Benes.scala 89:27]
    .io_y(in_switch_24_io_y),
    .io_z(in_switch_24_io_z),
    .io_in(in_switch_24_io_in)
  );
  InputSwitch in_switch_25 ( // @[Benes.scala 89:27]
    .io_y(in_switch_25_io_y),
    .io_z(in_switch_25_io_z),
    .io_in(in_switch_25_io_in)
  );
  InputSwitch in_switch_26 ( // @[Benes.scala 89:27]
    .io_y(in_switch_26_io_y),
    .io_z(in_switch_26_io_z),
    .io_in(in_switch_26_io_in)
  );
  InputSwitch in_switch_27 ( // @[Benes.scala 89:27]
    .io_y(in_switch_27_io_y),
    .io_z(in_switch_27_io_z),
    .io_in(in_switch_27_io_in)
  );
  InputSwitch in_switch_28 ( // @[Benes.scala 89:27]
    .io_y(in_switch_28_io_y),
    .io_z(in_switch_28_io_z),
    .io_in(in_switch_28_io_in)
  );
  InputSwitch in_switch_29 ( // @[Benes.scala 89:27]
    .io_y(in_switch_29_io_y),
    .io_z(in_switch_29_io_z),
    .io_in(in_switch_29_io_in)
  );
  InputSwitch in_switch_30 ( // @[Benes.scala 89:27]
    .io_y(in_switch_30_io_y),
    .io_z(in_switch_30_io_z),
    .io_in(in_switch_30_io_in)
  );
  InputSwitch in_switch_31 ( // @[Benes.scala 89:27]
    .io_y(in_switch_31_io_y),
    .io_z(in_switch_31_io_z),
    .io_in(in_switch_31_io_in)
  );
  OutputSwitch out_switch ( // @[Benes.scala 98:28]
    .io_y(out_switch_io_y),
    .io_in0(out_switch_io_in0),
    .io_in1(out_switch_io_in1),
    .io_sel(out_switch_io_sel)
  );
  OutputSwitch out_switch_1 ( // @[Benes.scala 98:28]
    .io_y(out_switch_1_io_y),
    .io_in0(out_switch_1_io_in0),
    .io_in1(out_switch_1_io_in1),
    .io_sel(out_switch_1_io_sel)
  );
  OutputSwitch out_switch_2 ( // @[Benes.scala 98:28]
    .io_y(out_switch_2_io_y),
    .io_in0(out_switch_2_io_in0),
    .io_in1(out_switch_2_io_in1),
    .io_sel(out_switch_2_io_sel)
  );
  OutputSwitch out_switch_3 ( // @[Benes.scala 98:28]
    .io_y(out_switch_3_io_y),
    .io_in0(out_switch_3_io_in0),
    .io_in1(out_switch_3_io_in1),
    .io_sel(out_switch_3_io_sel)
  );
  OutputSwitch out_switch_4 ( // @[Benes.scala 98:28]
    .io_y(out_switch_4_io_y),
    .io_in0(out_switch_4_io_in0),
    .io_in1(out_switch_4_io_in1),
    .io_sel(out_switch_4_io_sel)
  );
  OutputSwitch out_switch_5 ( // @[Benes.scala 98:28]
    .io_y(out_switch_5_io_y),
    .io_in0(out_switch_5_io_in0),
    .io_in1(out_switch_5_io_in1),
    .io_sel(out_switch_5_io_sel)
  );
  OutputSwitch out_switch_6 ( // @[Benes.scala 98:28]
    .io_y(out_switch_6_io_y),
    .io_in0(out_switch_6_io_in0),
    .io_in1(out_switch_6_io_in1),
    .io_sel(out_switch_6_io_sel)
  );
  OutputSwitch out_switch_7 ( // @[Benes.scala 98:28]
    .io_y(out_switch_7_io_y),
    .io_in0(out_switch_7_io_in0),
    .io_in1(out_switch_7_io_in1),
    .io_sel(out_switch_7_io_sel)
  );
  OutputSwitch out_switch_8 ( // @[Benes.scala 98:28]
    .io_y(out_switch_8_io_y),
    .io_in0(out_switch_8_io_in0),
    .io_in1(out_switch_8_io_in1),
    .io_sel(out_switch_8_io_sel)
  );
  OutputSwitch out_switch_9 ( // @[Benes.scala 98:28]
    .io_y(out_switch_9_io_y),
    .io_in0(out_switch_9_io_in0),
    .io_in1(out_switch_9_io_in1),
    .io_sel(out_switch_9_io_sel)
  );
  OutputSwitch out_switch_10 ( // @[Benes.scala 98:28]
    .io_y(out_switch_10_io_y),
    .io_in0(out_switch_10_io_in0),
    .io_in1(out_switch_10_io_in1),
    .io_sel(out_switch_10_io_sel)
  );
  OutputSwitch out_switch_11 ( // @[Benes.scala 98:28]
    .io_y(out_switch_11_io_y),
    .io_in0(out_switch_11_io_in0),
    .io_in1(out_switch_11_io_in1),
    .io_sel(out_switch_11_io_sel)
  );
  OutputSwitch out_switch_12 ( // @[Benes.scala 98:28]
    .io_y(out_switch_12_io_y),
    .io_in0(out_switch_12_io_in0),
    .io_in1(out_switch_12_io_in1),
    .io_sel(out_switch_12_io_sel)
  );
  OutputSwitch out_switch_13 ( // @[Benes.scala 98:28]
    .io_y(out_switch_13_io_y),
    .io_in0(out_switch_13_io_in0),
    .io_in1(out_switch_13_io_in1),
    .io_sel(out_switch_13_io_sel)
  );
  OutputSwitch out_switch_14 ( // @[Benes.scala 98:28]
    .io_y(out_switch_14_io_y),
    .io_in0(out_switch_14_io_in0),
    .io_in1(out_switch_14_io_in1),
    .io_sel(out_switch_14_io_sel)
  );
  OutputSwitch out_switch_15 ( // @[Benes.scala 98:28]
    .io_y(out_switch_15_io_y),
    .io_in0(out_switch_15_io_in0),
    .io_in1(out_switch_15_io_in1),
    .io_sel(out_switch_15_io_sel)
  );
  OutputSwitch out_switch_16 ( // @[Benes.scala 98:28]
    .io_y(out_switch_16_io_y),
    .io_in0(out_switch_16_io_in0),
    .io_in1(out_switch_16_io_in1),
    .io_sel(out_switch_16_io_sel)
  );
  OutputSwitch out_switch_17 ( // @[Benes.scala 98:28]
    .io_y(out_switch_17_io_y),
    .io_in0(out_switch_17_io_in0),
    .io_in1(out_switch_17_io_in1),
    .io_sel(out_switch_17_io_sel)
  );
  OutputSwitch out_switch_18 ( // @[Benes.scala 98:28]
    .io_y(out_switch_18_io_y),
    .io_in0(out_switch_18_io_in0),
    .io_in1(out_switch_18_io_in1),
    .io_sel(out_switch_18_io_sel)
  );
  OutputSwitch out_switch_19 ( // @[Benes.scala 98:28]
    .io_y(out_switch_19_io_y),
    .io_in0(out_switch_19_io_in0),
    .io_in1(out_switch_19_io_in1),
    .io_sel(out_switch_19_io_sel)
  );
  OutputSwitch out_switch_20 ( // @[Benes.scala 98:28]
    .io_y(out_switch_20_io_y),
    .io_in0(out_switch_20_io_in0),
    .io_in1(out_switch_20_io_in1),
    .io_sel(out_switch_20_io_sel)
  );
  OutputSwitch out_switch_21 ( // @[Benes.scala 98:28]
    .io_y(out_switch_21_io_y),
    .io_in0(out_switch_21_io_in0),
    .io_in1(out_switch_21_io_in1),
    .io_sel(out_switch_21_io_sel)
  );
  OutputSwitch out_switch_22 ( // @[Benes.scala 98:28]
    .io_y(out_switch_22_io_y),
    .io_in0(out_switch_22_io_in0),
    .io_in1(out_switch_22_io_in1),
    .io_sel(out_switch_22_io_sel)
  );
  OutputSwitch out_switch_23 ( // @[Benes.scala 98:28]
    .io_y(out_switch_23_io_y),
    .io_in0(out_switch_23_io_in0),
    .io_in1(out_switch_23_io_in1),
    .io_sel(out_switch_23_io_sel)
  );
  OutputSwitch out_switch_24 ( // @[Benes.scala 98:28]
    .io_y(out_switch_24_io_y),
    .io_in0(out_switch_24_io_in0),
    .io_in1(out_switch_24_io_in1),
    .io_sel(out_switch_24_io_sel)
  );
  OutputSwitch out_switch_25 ( // @[Benes.scala 98:28]
    .io_y(out_switch_25_io_y),
    .io_in0(out_switch_25_io_in0),
    .io_in1(out_switch_25_io_in1),
    .io_sel(out_switch_25_io_sel)
  );
  OutputSwitch out_switch_26 ( // @[Benes.scala 98:28]
    .io_y(out_switch_26_io_y),
    .io_in0(out_switch_26_io_in0),
    .io_in1(out_switch_26_io_in1),
    .io_sel(out_switch_26_io_sel)
  );
  OutputSwitch out_switch_27 ( // @[Benes.scala 98:28]
    .io_y(out_switch_27_io_y),
    .io_in0(out_switch_27_io_in0),
    .io_in1(out_switch_27_io_in1),
    .io_sel(out_switch_27_io_sel)
  );
  OutputSwitch out_switch_28 ( // @[Benes.scala 98:28]
    .io_y(out_switch_28_io_y),
    .io_in0(out_switch_28_io_in0),
    .io_in1(out_switch_28_io_in1),
    .io_sel(out_switch_28_io_sel)
  );
  OutputSwitch out_switch_29 ( // @[Benes.scala 98:28]
    .io_y(out_switch_29_io_y),
    .io_in0(out_switch_29_io_in0),
    .io_in1(out_switch_29_io_in1),
    .io_sel(out_switch_29_io_sel)
  );
  OutputSwitch out_switch_30 ( // @[Benes.scala 98:28]
    .io_y(out_switch_30_io_y),
    .io_in0(out_switch_30_io_in0),
    .io_in1(out_switch_30_io_in1),
    .io_sel(out_switch_30_io_sel)
  );
  OutputSwitch out_switch_31 ( // @[Benes.scala 98:28]
    .io_y(out_switch_31_io_y),
    .io_in0(out_switch_31_io_in0),
    .io_in1(out_switch_31_io_in1),
    .io_sel(out_switch_31_io_sel)
  );
  Switch imm_switch ( // @[Benes.scala 108:30]
    .io_y(imm_switch_io_y),
    .io_z(imm_switch_io_z),
    .io_in0(imm_switch_io_in0),
    .io_in1(imm_switch_io_in1),
    .io_sel0(imm_switch_io_sel0),
    .io_sel1(imm_switch_io_sel1)
  );
  Switch imm_switch_1 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_1_io_y),
    .io_z(imm_switch_1_io_z),
    .io_in0(imm_switch_1_io_in0),
    .io_in1(imm_switch_1_io_in1),
    .io_sel0(imm_switch_1_io_sel0),
    .io_sel1(imm_switch_1_io_sel1)
  );
  Switch imm_switch_2 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_2_io_y),
    .io_z(imm_switch_2_io_z),
    .io_in0(imm_switch_2_io_in0),
    .io_in1(imm_switch_2_io_in1),
    .io_sel0(imm_switch_2_io_sel0),
    .io_sel1(imm_switch_2_io_sel1)
  );
  Switch imm_switch_3 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_3_io_y),
    .io_z(imm_switch_3_io_z),
    .io_in0(imm_switch_3_io_in0),
    .io_in1(imm_switch_3_io_in1),
    .io_sel0(imm_switch_3_io_sel0),
    .io_sel1(imm_switch_3_io_sel1)
  );
  Switch imm_switch_4 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_4_io_y),
    .io_z(imm_switch_4_io_z),
    .io_in0(imm_switch_4_io_in0),
    .io_in1(imm_switch_4_io_in1),
    .io_sel0(imm_switch_4_io_sel0),
    .io_sel1(imm_switch_4_io_sel1)
  );
  Switch imm_switch_5 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_5_io_y),
    .io_z(imm_switch_5_io_z),
    .io_in0(imm_switch_5_io_in0),
    .io_in1(imm_switch_5_io_in1),
    .io_sel0(imm_switch_5_io_sel0),
    .io_sel1(imm_switch_5_io_sel1)
  );
  Switch imm_switch_6 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_6_io_y),
    .io_z(imm_switch_6_io_z),
    .io_in0(imm_switch_6_io_in0),
    .io_in1(imm_switch_6_io_in1),
    .io_sel0(imm_switch_6_io_sel0),
    .io_sel1(imm_switch_6_io_sel1)
  );
  Switch imm_switch_7 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_7_io_y),
    .io_z(imm_switch_7_io_z),
    .io_in0(imm_switch_7_io_in0),
    .io_in1(imm_switch_7_io_in1),
    .io_sel0(imm_switch_7_io_sel0),
    .io_sel1(imm_switch_7_io_sel1)
  );
  Switch imm_switch_8 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_8_io_y),
    .io_z(imm_switch_8_io_z),
    .io_in0(imm_switch_8_io_in0),
    .io_in1(imm_switch_8_io_in1),
    .io_sel0(imm_switch_8_io_sel0),
    .io_sel1(imm_switch_8_io_sel1)
  );
  Switch imm_switch_9 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_9_io_y),
    .io_z(imm_switch_9_io_z),
    .io_in0(imm_switch_9_io_in0),
    .io_in1(imm_switch_9_io_in1),
    .io_sel0(imm_switch_9_io_sel0),
    .io_sel1(imm_switch_9_io_sel1)
  );
  Switch imm_switch_10 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_10_io_y),
    .io_z(imm_switch_10_io_z),
    .io_in0(imm_switch_10_io_in0),
    .io_in1(imm_switch_10_io_in1),
    .io_sel0(imm_switch_10_io_sel0),
    .io_sel1(imm_switch_10_io_sel1)
  );
  Switch imm_switch_11 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_11_io_y),
    .io_z(imm_switch_11_io_z),
    .io_in0(imm_switch_11_io_in0),
    .io_in1(imm_switch_11_io_in1),
    .io_sel0(imm_switch_11_io_sel0),
    .io_sel1(imm_switch_11_io_sel1)
  );
  Switch imm_switch_12 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_12_io_y),
    .io_z(imm_switch_12_io_z),
    .io_in0(imm_switch_12_io_in0),
    .io_in1(imm_switch_12_io_in1),
    .io_sel0(imm_switch_12_io_sel0),
    .io_sel1(imm_switch_12_io_sel1)
  );
  Switch imm_switch_13 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_13_io_y),
    .io_z(imm_switch_13_io_z),
    .io_in0(imm_switch_13_io_in0),
    .io_in1(imm_switch_13_io_in1),
    .io_sel0(imm_switch_13_io_sel0),
    .io_sel1(imm_switch_13_io_sel1)
  );
  Switch imm_switch_14 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_14_io_y),
    .io_z(imm_switch_14_io_z),
    .io_in0(imm_switch_14_io_in0),
    .io_in1(imm_switch_14_io_in1),
    .io_sel0(imm_switch_14_io_sel0),
    .io_sel1(imm_switch_14_io_sel1)
  );
  Switch imm_switch_15 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_15_io_y),
    .io_z(imm_switch_15_io_z),
    .io_in0(imm_switch_15_io_in0),
    .io_in1(imm_switch_15_io_in1),
    .io_sel0(imm_switch_15_io_sel0),
    .io_sel1(imm_switch_15_io_sel1)
  );
  Switch imm_switch_16 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_16_io_y),
    .io_z(imm_switch_16_io_z),
    .io_in0(imm_switch_16_io_in0),
    .io_in1(imm_switch_16_io_in1),
    .io_sel0(imm_switch_16_io_sel0),
    .io_sel1(imm_switch_16_io_sel1)
  );
  Switch imm_switch_17 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_17_io_y),
    .io_z(imm_switch_17_io_z),
    .io_in0(imm_switch_17_io_in0),
    .io_in1(imm_switch_17_io_in1),
    .io_sel0(imm_switch_17_io_sel0),
    .io_sel1(imm_switch_17_io_sel1)
  );
  Switch imm_switch_18 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_18_io_y),
    .io_z(imm_switch_18_io_z),
    .io_in0(imm_switch_18_io_in0),
    .io_in1(imm_switch_18_io_in1),
    .io_sel0(imm_switch_18_io_sel0),
    .io_sel1(imm_switch_18_io_sel1)
  );
  Switch imm_switch_19 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_19_io_y),
    .io_z(imm_switch_19_io_z),
    .io_in0(imm_switch_19_io_in0),
    .io_in1(imm_switch_19_io_in1),
    .io_sel0(imm_switch_19_io_sel0),
    .io_sel1(imm_switch_19_io_sel1)
  );
  Switch imm_switch_20 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_20_io_y),
    .io_z(imm_switch_20_io_z),
    .io_in0(imm_switch_20_io_in0),
    .io_in1(imm_switch_20_io_in1),
    .io_sel0(imm_switch_20_io_sel0),
    .io_sel1(imm_switch_20_io_sel1)
  );
  Switch imm_switch_21 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_21_io_y),
    .io_z(imm_switch_21_io_z),
    .io_in0(imm_switch_21_io_in0),
    .io_in1(imm_switch_21_io_in1),
    .io_sel0(imm_switch_21_io_sel0),
    .io_sel1(imm_switch_21_io_sel1)
  );
  Switch imm_switch_22 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_22_io_y),
    .io_z(imm_switch_22_io_z),
    .io_in0(imm_switch_22_io_in0),
    .io_in1(imm_switch_22_io_in1),
    .io_sel0(imm_switch_22_io_sel0),
    .io_sel1(imm_switch_22_io_sel1)
  );
  Switch imm_switch_23 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_23_io_y),
    .io_z(imm_switch_23_io_z),
    .io_in0(imm_switch_23_io_in0),
    .io_in1(imm_switch_23_io_in1),
    .io_sel0(imm_switch_23_io_sel0),
    .io_sel1(imm_switch_23_io_sel1)
  );
  Switch imm_switch_24 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_24_io_y),
    .io_z(imm_switch_24_io_z),
    .io_in0(imm_switch_24_io_in0),
    .io_in1(imm_switch_24_io_in1),
    .io_sel0(imm_switch_24_io_sel0),
    .io_sel1(imm_switch_24_io_sel1)
  );
  Switch imm_switch_25 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_25_io_y),
    .io_z(imm_switch_25_io_z),
    .io_in0(imm_switch_25_io_in0),
    .io_in1(imm_switch_25_io_in1),
    .io_sel0(imm_switch_25_io_sel0),
    .io_sel1(imm_switch_25_io_sel1)
  );
  Switch imm_switch_26 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_26_io_y),
    .io_z(imm_switch_26_io_z),
    .io_in0(imm_switch_26_io_in0),
    .io_in1(imm_switch_26_io_in1),
    .io_sel0(imm_switch_26_io_sel0),
    .io_sel1(imm_switch_26_io_sel1)
  );
  Switch imm_switch_27 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_27_io_y),
    .io_z(imm_switch_27_io_z),
    .io_in0(imm_switch_27_io_in0),
    .io_in1(imm_switch_27_io_in1),
    .io_sel0(imm_switch_27_io_sel0),
    .io_sel1(imm_switch_27_io_sel1)
  );
  Switch imm_switch_28 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_28_io_y),
    .io_z(imm_switch_28_io_z),
    .io_in0(imm_switch_28_io_in0),
    .io_in1(imm_switch_28_io_in1),
    .io_sel0(imm_switch_28_io_sel0),
    .io_sel1(imm_switch_28_io_sel1)
  );
  Switch imm_switch_29 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_29_io_y),
    .io_z(imm_switch_29_io_z),
    .io_in0(imm_switch_29_io_in0),
    .io_in1(imm_switch_29_io_in1),
    .io_sel0(imm_switch_29_io_sel0),
    .io_sel1(imm_switch_29_io_sel1)
  );
  Switch imm_switch_30 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_30_io_y),
    .io_z(imm_switch_30_io_z),
    .io_in0(imm_switch_30_io_in0),
    .io_in1(imm_switch_30_io_in1),
    .io_sel0(imm_switch_30_io_sel0),
    .io_sel1(imm_switch_30_io_sel1)
  );
  Switch imm_switch_31 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_31_io_y),
    .io_z(imm_switch_31_io_z),
    .io_in0(imm_switch_31_io_in0),
    .io_in1(imm_switch_31_io_in1),
    .io_sel0(imm_switch_31_io_sel0),
    .io_sel1(imm_switch_31_io_sel1)
  );
  Switch imm_switch_32 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_32_io_y),
    .io_z(imm_switch_32_io_z),
    .io_in0(imm_switch_32_io_in0),
    .io_in1(imm_switch_32_io_in1),
    .io_sel0(imm_switch_32_io_sel0),
    .io_sel1(imm_switch_32_io_sel1)
  );
  Switch imm_switch_33 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_33_io_y),
    .io_z(imm_switch_33_io_z),
    .io_in0(imm_switch_33_io_in0),
    .io_in1(imm_switch_33_io_in1),
    .io_sel0(imm_switch_33_io_sel0),
    .io_sel1(imm_switch_33_io_sel1)
  );
  Switch imm_switch_34 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_34_io_y),
    .io_z(imm_switch_34_io_z),
    .io_in0(imm_switch_34_io_in0),
    .io_in1(imm_switch_34_io_in1),
    .io_sel0(imm_switch_34_io_sel0),
    .io_sel1(imm_switch_34_io_sel1)
  );
  Switch imm_switch_35 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_35_io_y),
    .io_z(imm_switch_35_io_z),
    .io_in0(imm_switch_35_io_in0),
    .io_in1(imm_switch_35_io_in1),
    .io_sel0(imm_switch_35_io_sel0),
    .io_sel1(imm_switch_35_io_sel1)
  );
  Switch imm_switch_36 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_36_io_y),
    .io_z(imm_switch_36_io_z),
    .io_in0(imm_switch_36_io_in0),
    .io_in1(imm_switch_36_io_in1),
    .io_sel0(imm_switch_36_io_sel0),
    .io_sel1(imm_switch_36_io_sel1)
  );
  Switch imm_switch_37 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_37_io_y),
    .io_z(imm_switch_37_io_z),
    .io_in0(imm_switch_37_io_in0),
    .io_in1(imm_switch_37_io_in1),
    .io_sel0(imm_switch_37_io_sel0),
    .io_sel1(imm_switch_37_io_sel1)
  );
  Switch imm_switch_38 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_38_io_y),
    .io_z(imm_switch_38_io_z),
    .io_in0(imm_switch_38_io_in0),
    .io_in1(imm_switch_38_io_in1),
    .io_sel0(imm_switch_38_io_sel0),
    .io_sel1(imm_switch_38_io_sel1)
  );
  Switch imm_switch_39 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_39_io_y),
    .io_z(imm_switch_39_io_z),
    .io_in0(imm_switch_39_io_in0),
    .io_in1(imm_switch_39_io_in1),
    .io_sel0(imm_switch_39_io_sel0),
    .io_sel1(imm_switch_39_io_sel1)
  );
  Switch imm_switch_40 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_40_io_y),
    .io_z(imm_switch_40_io_z),
    .io_in0(imm_switch_40_io_in0),
    .io_in1(imm_switch_40_io_in1),
    .io_sel0(imm_switch_40_io_sel0),
    .io_sel1(imm_switch_40_io_sel1)
  );
  Switch imm_switch_41 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_41_io_y),
    .io_z(imm_switch_41_io_z),
    .io_in0(imm_switch_41_io_in0),
    .io_in1(imm_switch_41_io_in1),
    .io_sel0(imm_switch_41_io_sel0),
    .io_sel1(imm_switch_41_io_sel1)
  );
  Switch imm_switch_42 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_42_io_y),
    .io_z(imm_switch_42_io_z),
    .io_in0(imm_switch_42_io_in0),
    .io_in1(imm_switch_42_io_in1),
    .io_sel0(imm_switch_42_io_sel0),
    .io_sel1(imm_switch_42_io_sel1)
  );
  Switch imm_switch_43 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_43_io_y),
    .io_z(imm_switch_43_io_z),
    .io_in0(imm_switch_43_io_in0),
    .io_in1(imm_switch_43_io_in1),
    .io_sel0(imm_switch_43_io_sel0),
    .io_sel1(imm_switch_43_io_sel1)
  );
  Switch imm_switch_44 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_44_io_y),
    .io_z(imm_switch_44_io_z),
    .io_in0(imm_switch_44_io_in0),
    .io_in1(imm_switch_44_io_in1),
    .io_sel0(imm_switch_44_io_sel0),
    .io_sel1(imm_switch_44_io_sel1)
  );
  Switch imm_switch_45 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_45_io_y),
    .io_z(imm_switch_45_io_z),
    .io_in0(imm_switch_45_io_in0),
    .io_in1(imm_switch_45_io_in1),
    .io_sel0(imm_switch_45_io_sel0),
    .io_sel1(imm_switch_45_io_sel1)
  );
  Switch imm_switch_46 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_46_io_y),
    .io_z(imm_switch_46_io_z),
    .io_in0(imm_switch_46_io_in0),
    .io_in1(imm_switch_46_io_in1),
    .io_sel0(imm_switch_46_io_sel0),
    .io_sel1(imm_switch_46_io_sel1)
  );
  Switch imm_switch_47 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_47_io_y),
    .io_z(imm_switch_47_io_z),
    .io_in0(imm_switch_47_io_in0),
    .io_in1(imm_switch_47_io_in1),
    .io_sel0(imm_switch_47_io_sel0),
    .io_sel1(imm_switch_47_io_sel1)
  );
  Switch imm_switch_48 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_48_io_y),
    .io_z(imm_switch_48_io_z),
    .io_in0(imm_switch_48_io_in0),
    .io_in1(imm_switch_48_io_in1),
    .io_sel0(imm_switch_48_io_sel0),
    .io_sel1(imm_switch_48_io_sel1)
  );
  Switch imm_switch_49 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_49_io_y),
    .io_z(imm_switch_49_io_z),
    .io_in0(imm_switch_49_io_in0),
    .io_in1(imm_switch_49_io_in1),
    .io_sel0(imm_switch_49_io_sel0),
    .io_sel1(imm_switch_49_io_sel1)
  );
  Switch imm_switch_50 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_50_io_y),
    .io_z(imm_switch_50_io_z),
    .io_in0(imm_switch_50_io_in0),
    .io_in1(imm_switch_50_io_in1),
    .io_sel0(imm_switch_50_io_sel0),
    .io_sel1(imm_switch_50_io_sel1)
  );
  Switch imm_switch_51 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_51_io_y),
    .io_z(imm_switch_51_io_z),
    .io_in0(imm_switch_51_io_in0),
    .io_in1(imm_switch_51_io_in1),
    .io_sel0(imm_switch_51_io_sel0),
    .io_sel1(imm_switch_51_io_sel1)
  );
  Switch imm_switch_52 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_52_io_y),
    .io_z(imm_switch_52_io_z),
    .io_in0(imm_switch_52_io_in0),
    .io_in1(imm_switch_52_io_in1),
    .io_sel0(imm_switch_52_io_sel0),
    .io_sel1(imm_switch_52_io_sel1)
  );
  Switch imm_switch_53 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_53_io_y),
    .io_z(imm_switch_53_io_z),
    .io_in0(imm_switch_53_io_in0),
    .io_in1(imm_switch_53_io_in1),
    .io_sel0(imm_switch_53_io_sel0),
    .io_sel1(imm_switch_53_io_sel1)
  );
  Switch imm_switch_54 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_54_io_y),
    .io_z(imm_switch_54_io_z),
    .io_in0(imm_switch_54_io_in0),
    .io_in1(imm_switch_54_io_in1),
    .io_sel0(imm_switch_54_io_sel0),
    .io_sel1(imm_switch_54_io_sel1)
  );
  Switch imm_switch_55 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_55_io_y),
    .io_z(imm_switch_55_io_z),
    .io_in0(imm_switch_55_io_in0),
    .io_in1(imm_switch_55_io_in1),
    .io_sel0(imm_switch_55_io_sel0),
    .io_sel1(imm_switch_55_io_sel1)
  );
  Switch imm_switch_56 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_56_io_y),
    .io_z(imm_switch_56_io_z),
    .io_in0(imm_switch_56_io_in0),
    .io_in1(imm_switch_56_io_in1),
    .io_sel0(imm_switch_56_io_sel0),
    .io_sel1(imm_switch_56_io_sel1)
  );
  Switch imm_switch_57 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_57_io_y),
    .io_z(imm_switch_57_io_z),
    .io_in0(imm_switch_57_io_in0),
    .io_in1(imm_switch_57_io_in1),
    .io_sel0(imm_switch_57_io_sel0),
    .io_sel1(imm_switch_57_io_sel1)
  );
  Switch imm_switch_58 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_58_io_y),
    .io_z(imm_switch_58_io_z),
    .io_in0(imm_switch_58_io_in0),
    .io_in1(imm_switch_58_io_in1),
    .io_sel0(imm_switch_58_io_sel0),
    .io_sel1(imm_switch_58_io_sel1)
  );
  Switch imm_switch_59 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_59_io_y),
    .io_z(imm_switch_59_io_z),
    .io_in0(imm_switch_59_io_in0),
    .io_in1(imm_switch_59_io_in1),
    .io_sel0(imm_switch_59_io_sel0),
    .io_sel1(imm_switch_59_io_sel1)
  );
  Switch imm_switch_60 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_60_io_y),
    .io_z(imm_switch_60_io_z),
    .io_in0(imm_switch_60_io_in0),
    .io_in1(imm_switch_60_io_in1),
    .io_sel0(imm_switch_60_io_sel0),
    .io_sel1(imm_switch_60_io_sel1)
  );
  Switch imm_switch_61 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_61_io_y),
    .io_z(imm_switch_61_io_z),
    .io_in0(imm_switch_61_io_in0),
    .io_in1(imm_switch_61_io_in1),
    .io_sel0(imm_switch_61_io_sel0),
    .io_sel1(imm_switch_61_io_sel1)
  );
  Switch imm_switch_62 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_62_io_y),
    .io_z(imm_switch_62_io_z),
    .io_in0(imm_switch_62_io_in0),
    .io_in1(imm_switch_62_io_in1),
    .io_sel0(imm_switch_62_io_sel0),
    .io_sel1(imm_switch_62_io_sel1)
  );
  Switch imm_switch_63 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_63_io_y),
    .io_z(imm_switch_63_io_z),
    .io_in0(imm_switch_63_io_in0),
    .io_in1(imm_switch_63_io_in1),
    .io_sel0(imm_switch_63_io_sel0),
    .io_sel1(imm_switch_63_io_sel1)
  );
  Switch imm_switch_64 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_64_io_y),
    .io_z(imm_switch_64_io_z),
    .io_in0(imm_switch_64_io_in0),
    .io_in1(imm_switch_64_io_in1),
    .io_sel0(imm_switch_64_io_sel0),
    .io_sel1(imm_switch_64_io_sel1)
  );
  Switch imm_switch_65 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_65_io_y),
    .io_z(imm_switch_65_io_z),
    .io_in0(imm_switch_65_io_in0),
    .io_in1(imm_switch_65_io_in1),
    .io_sel0(imm_switch_65_io_sel0),
    .io_sel1(imm_switch_65_io_sel1)
  );
  Switch imm_switch_66 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_66_io_y),
    .io_z(imm_switch_66_io_z),
    .io_in0(imm_switch_66_io_in0),
    .io_in1(imm_switch_66_io_in1),
    .io_sel0(imm_switch_66_io_sel0),
    .io_sel1(imm_switch_66_io_sel1)
  );
  Switch imm_switch_67 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_67_io_y),
    .io_z(imm_switch_67_io_z),
    .io_in0(imm_switch_67_io_in0),
    .io_in1(imm_switch_67_io_in1),
    .io_sel0(imm_switch_67_io_sel0),
    .io_sel1(imm_switch_67_io_sel1)
  );
  Switch imm_switch_68 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_68_io_y),
    .io_z(imm_switch_68_io_z),
    .io_in0(imm_switch_68_io_in0),
    .io_in1(imm_switch_68_io_in1),
    .io_sel0(imm_switch_68_io_sel0),
    .io_sel1(imm_switch_68_io_sel1)
  );
  Switch imm_switch_69 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_69_io_y),
    .io_z(imm_switch_69_io_z),
    .io_in0(imm_switch_69_io_in0),
    .io_in1(imm_switch_69_io_in1),
    .io_sel0(imm_switch_69_io_sel0),
    .io_sel1(imm_switch_69_io_sel1)
  );
  Switch imm_switch_70 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_70_io_y),
    .io_z(imm_switch_70_io_z),
    .io_in0(imm_switch_70_io_in0),
    .io_in1(imm_switch_70_io_in1),
    .io_sel0(imm_switch_70_io_sel0),
    .io_sel1(imm_switch_70_io_sel1)
  );
  Switch imm_switch_71 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_71_io_y),
    .io_z(imm_switch_71_io_z),
    .io_in0(imm_switch_71_io_in0),
    .io_in1(imm_switch_71_io_in1),
    .io_sel0(imm_switch_71_io_sel0),
    .io_sel1(imm_switch_71_io_sel1)
  );
  Switch imm_switch_72 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_72_io_y),
    .io_z(imm_switch_72_io_z),
    .io_in0(imm_switch_72_io_in0),
    .io_in1(imm_switch_72_io_in1),
    .io_sel0(imm_switch_72_io_sel0),
    .io_sel1(imm_switch_72_io_sel1)
  );
  Switch imm_switch_73 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_73_io_y),
    .io_z(imm_switch_73_io_z),
    .io_in0(imm_switch_73_io_in0),
    .io_in1(imm_switch_73_io_in1),
    .io_sel0(imm_switch_73_io_sel0),
    .io_sel1(imm_switch_73_io_sel1)
  );
  Switch imm_switch_74 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_74_io_y),
    .io_z(imm_switch_74_io_z),
    .io_in0(imm_switch_74_io_in0),
    .io_in1(imm_switch_74_io_in1),
    .io_sel0(imm_switch_74_io_sel0),
    .io_sel1(imm_switch_74_io_sel1)
  );
  Switch imm_switch_75 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_75_io_y),
    .io_z(imm_switch_75_io_z),
    .io_in0(imm_switch_75_io_in0),
    .io_in1(imm_switch_75_io_in1),
    .io_sel0(imm_switch_75_io_sel0),
    .io_sel1(imm_switch_75_io_sel1)
  );
  Switch imm_switch_76 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_76_io_y),
    .io_z(imm_switch_76_io_z),
    .io_in0(imm_switch_76_io_in0),
    .io_in1(imm_switch_76_io_in1),
    .io_sel0(imm_switch_76_io_sel0),
    .io_sel1(imm_switch_76_io_sel1)
  );
  Switch imm_switch_77 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_77_io_y),
    .io_z(imm_switch_77_io_z),
    .io_in0(imm_switch_77_io_in0),
    .io_in1(imm_switch_77_io_in1),
    .io_sel0(imm_switch_77_io_sel0),
    .io_sel1(imm_switch_77_io_sel1)
  );
  Switch imm_switch_78 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_78_io_y),
    .io_z(imm_switch_78_io_z),
    .io_in0(imm_switch_78_io_in0),
    .io_in1(imm_switch_78_io_in1),
    .io_sel0(imm_switch_78_io_sel0),
    .io_sel1(imm_switch_78_io_sel1)
  );
  Switch imm_switch_79 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_79_io_y),
    .io_z(imm_switch_79_io_z),
    .io_in0(imm_switch_79_io_in0),
    .io_in1(imm_switch_79_io_in1),
    .io_sel0(imm_switch_79_io_sel0),
    .io_sel1(imm_switch_79_io_sel1)
  );
  Switch imm_switch_80 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_80_io_y),
    .io_z(imm_switch_80_io_z),
    .io_in0(imm_switch_80_io_in0),
    .io_in1(imm_switch_80_io_in1),
    .io_sel0(imm_switch_80_io_sel0),
    .io_sel1(imm_switch_80_io_sel1)
  );
  Switch imm_switch_81 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_81_io_y),
    .io_z(imm_switch_81_io_z),
    .io_in0(imm_switch_81_io_in0),
    .io_in1(imm_switch_81_io_in1),
    .io_sel0(imm_switch_81_io_sel0),
    .io_sel1(imm_switch_81_io_sel1)
  );
  Switch imm_switch_82 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_82_io_y),
    .io_z(imm_switch_82_io_z),
    .io_in0(imm_switch_82_io_in0),
    .io_in1(imm_switch_82_io_in1),
    .io_sel0(imm_switch_82_io_sel0),
    .io_sel1(imm_switch_82_io_sel1)
  );
  Switch imm_switch_83 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_83_io_y),
    .io_z(imm_switch_83_io_z),
    .io_in0(imm_switch_83_io_in0),
    .io_in1(imm_switch_83_io_in1),
    .io_sel0(imm_switch_83_io_sel0),
    .io_sel1(imm_switch_83_io_sel1)
  );
  Switch imm_switch_84 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_84_io_y),
    .io_z(imm_switch_84_io_z),
    .io_in0(imm_switch_84_io_in0),
    .io_in1(imm_switch_84_io_in1),
    .io_sel0(imm_switch_84_io_sel0),
    .io_sel1(imm_switch_84_io_sel1)
  );
  Switch imm_switch_85 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_85_io_y),
    .io_z(imm_switch_85_io_z),
    .io_in0(imm_switch_85_io_in0),
    .io_in1(imm_switch_85_io_in1),
    .io_sel0(imm_switch_85_io_sel0),
    .io_sel1(imm_switch_85_io_sel1)
  );
  Switch imm_switch_86 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_86_io_y),
    .io_z(imm_switch_86_io_z),
    .io_in0(imm_switch_86_io_in0),
    .io_in1(imm_switch_86_io_in1),
    .io_sel0(imm_switch_86_io_sel0),
    .io_sel1(imm_switch_86_io_sel1)
  );
  Switch imm_switch_87 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_87_io_y),
    .io_z(imm_switch_87_io_z),
    .io_in0(imm_switch_87_io_in0),
    .io_in1(imm_switch_87_io_in1),
    .io_sel0(imm_switch_87_io_sel0),
    .io_sel1(imm_switch_87_io_sel1)
  );
  Switch imm_switch_88 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_88_io_y),
    .io_z(imm_switch_88_io_z),
    .io_in0(imm_switch_88_io_in0),
    .io_in1(imm_switch_88_io_in1),
    .io_sel0(imm_switch_88_io_sel0),
    .io_sel1(imm_switch_88_io_sel1)
  );
  Switch imm_switch_89 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_89_io_y),
    .io_z(imm_switch_89_io_z),
    .io_in0(imm_switch_89_io_in0),
    .io_in1(imm_switch_89_io_in1),
    .io_sel0(imm_switch_89_io_sel0),
    .io_sel1(imm_switch_89_io_sel1)
  );
  Switch imm_switch_90 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_90_io_y),
    .io_z(imm_switch_90_io_z),
    .io_in0(imm_switch_90_io_in0),
    .io_in1(imm_switch_90_io_in1),
    .io_sel0(imm_switch_90_io_sel0),
    .io_sel1(imm_switch_90_io_sel1)
  );
  Switch imm_switch_91 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_91_io_y),
    .io_z(imm_switch_91_io_z),
    .io_in0(imm_switch_91_io_in0),
    .io_in1(imm_switch_91_io_in1),
    .io_sel0(imm_switch_91_io_sel0),
    .io_sel1(imm_switch_91_io_sel1)
  );
  Switch imm_switch_92 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_92_io_y),
    .io_z(imm_switch_92_io_z),
    .io_in0(imm_switch_92_io_in0),
    .io_in1(imm_switch_92_io_in1),
    .io_sel0(imm_switch_92_io_sel0),
    .io_sel1(imm_switch_92_io_sel1)
  );
  Switch imm_switch_93 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_93_io_y),
    .io_z(imm_switch_93_io_z),
    .io_in0(imm_switch_93_io_in0),
    .io_in1(imm_switch_93_io_in1),
    .io_sel0(imm_switch_93_io_sel0),
    .io_sel1(imm_switch_93_io_sel1)
  );
  Switch imm_switch_94 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_94_io_y),
    .io_z(imm_switch_94_io_z),
    .io_in0(imm_switch_94_io_in0),
    .io_in1(imm_switch_94_io_in1),
    .io_sel0(imm_switch_94_io_sel0),
    .io_sel1(imm_switch_94_io_sel1)
  );
  Switch imm_switch_95 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_95_io_y),
    .io_z(imm_switch_95_io_z),
    .io_in0(imm_switch_95_io_in0),
    .io_in1(imm_switch_95_io_in1),
    .io_sel0(imm_switch_95_io_sel0),
    .io_sel1(imm_switch_95_io_sel1)
  );
  Switch imm_switch_96 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_96_io_y),
    .io_z(imm_switch_96_io_z),
    .io_in0(imm_switch_96_io_in0),
    .io_in1(imm_switch_96_io_in1),
    .io_sel0(imm_switch_96_io_sel0),
    .io_sel1(imm_switch_96_io_sel1)
  );
  Switch imm_switch_97 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_97_io_y),
    .io_z(imm_switch_97_io_z),
    .io_in0(imm_switch_97_io_in0),
    .io_in1(imm_switch_97_io_in1),
    .io_sel0(imm_switch_97_io_sel0),
    .io_sel1(imm_switch_97_io_sel1)
  );
  Switch imm_switch_98 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_98_io_y),
    .io_z(imm_switch_98_io_z),
    .io_in0(imm_switch_98_io_in0),
    .io_in1(imm_switch_98_io_in1),
    .io_sel0(imm_switch_98_io_sel0),
    .io_sel1(imm_switch_98_io_sel1)
  );
  Switch imm_switch_99 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_99_io_y),
    .io_z(imm_switch_99_io_z),
    .io_in0(imm_switch_99_io_in0),
    .io_in1(imm_switch_99_io_in1),
    .io_sel0(imm_switch_99_io_sel0),
    .io_sel1(imm_switch_99_io_sel1)
  );
  Switch imm_switch_100 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_100_io_y),
    .io_z(imm_switch_100_io_z),
    .io_in0(imm_switch_100_io_in0),
    .io_in1(imm_switch_100_io_in1),
    .io_sel0(imm_switch_100_io_sel0),
    .io_sel1(imm_switch_100_io_sel1)
  );
  Switch imm_switch_101 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_101_io_y),
    .io_z(imm_switch_101_io_z),
    .io_in0(imm_switch_101_io_in0),
    .io_in1(imm_switch_101_io_in1),
    .io_sel0(imm_switch_101_io_sel0),
    .io_sel1(imm_switch_101_io_sel1)
  );
  Switch imm_switch_102 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_102_io_y),
    .io_z(imm_switch_102_io_z),
    .io_in0(imm_switch_102_io_in0),
    .io_in1(imm_switch_102_io_in1),
    .io_sel0(imm_switch_102_io_sel0),
    .io_sel1(imm_switch_102_io_sel1)
  );
  Switch imm_switch_103 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_103_io_y),
    .io_z(imm_switch_103_io_z),
    .io_in0(imm_switch_103_io_in0),
    .io_in1(imm_switch_103_io_in1),
    .io_sel0(imm_switch_103_io_sel0),
    .io_sel1(imm_switch_103_io_sel1)
  );
  Switch imm_switch_104 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_104_io_y),
    .io_z(imm_switch_104_io_z),
    .io_in0(imm_switch_104_io_in0),
    .io_in1(imm_switch_104_io_in1),
    .io_sel0(imm_switch_104_io_sel0),
    .io_sel1(imm_switch_104_io_sel1)
  );
  Switch imm_switch_105 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_105_io_y),
    .io_z(imm_switch_105_io_z),
    .io_in0(imm_switch_105_io_in0),
    .io_in1(imm_switch_105_io_in1),
    .io_sel0(imm_switch_105_io_sel0),
    .io_sel1(imm_switch_105_io_sel1)
  );
  Switch imm_switch_106 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_106_io_y),
    .io_z(imm_switch_106_io_z),
    .io_in0(imm_switch_106_io_in0),
    .io_in1(imm_switch_106_io_in1),
    .io_sel0(imm_switch_106_io_sel0),
    .io_sel1(imm_switch_106_io_sel1)
  );
  Switch imm_switch_107 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_107_io_y),
    .io_z(imm_switch_107_io_z),
    .io_in0(imm_switch_107_io_in0),
    .io_in1(imm_switch_107_io_in1),
    .io_sel0(imm_switch_107_io_sel0),
    .io_sel1(imm_switch_107_io_sel1)
  );
  Switch imm_switch_108 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_108_io_y),
    .io_z(imm_switch_108_io_z),
    .io_in0(imm_switch_108_io_in0),
    .io_in1(imm_switch_108_io_in1),
    .io_sel0(imm_switch_108_io_sel0),
    .io_sel1(imm_switch_108_io_sel1)
  );
  Switch imm_switch_109 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_109_io_y),
    .io_z(imm_switch_109_io_z),
    .io_in0(imm_switch_109_io_in0),
    .io_in1(imm_switch_109_io_in1),
    .io_sel0(imm_switch_109_io_sel0),
    .io_sel1(imm_switch_109_io_sel1)
  );
  Switch imm_switch_110 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_110_io_y),
    .io_z(imm_switch_110_io_z),
    .io_in0(imm_switch_110_io_in0),
    .io_in1(imm_switch_110_io_in1),
    .io_sel0(imm_switch_110_io_sel0),
    .io_sel1(imm_switch_110_io_sel1)
  );
  Switch imm_switch_111 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_111_io_y),
    .io_z(imm_switch_111_io_z),
    .io_in0(imm_switch_111_io_in0),
    .io_in1(imm_switch_111_io_in1),
    .io_sel0(imm_switch_111_io_sel0),
    .io_sel1(imm_switch_111_io_sel1)
  );
  Switch imm_switch_112 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_112_io_y),
    .io_z(imm_switch_112_io_z),
    .io_in0(imm_switch_112_io_in0),
    .io_in1(imm_switch_112_io_in1),
    .io_sel0(imm_switch_112_io_sel0),
    .io_sel1(imm_switch_112_io_sel1)
  );
  Switch imm_switch_113 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_113_io_y),
    .io_z(imm_switch_113_io_z),
    .io_in0(imm_switch_113_io_in0),
    .io_in1(imm_switch_113_io_in1),
    .io_sel0(imm_switch_113_io_sel0),
    .io_sel1(imm_switch_113_io_sel1)
  );
  Switch imm_switch_114 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_114_io_y),
    .io_z(imm_switch_114_io_z),
    .io_in0(imm_switch_114_io_in0),
    .io_in1(imm_switch_114_io_in1),
    .io_sel0(imm_switch_114_io_sel0),
    .io_sel1(imm_switch_114_io_sel1)
  );
  Switch imm_switch_115 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_115_io_y),
    .io_z(imm_switch_115_io_z),
    .io_in0(imm_switch_115_io_in0),
    .io_in1(imm_switch_115_io_in1),
    .io_sel0(imm_switch_115_io_sel0),
    .io_sel1(imm_switch_115_io_sel1)
  );
  Switch imm_switch_116 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_116_io_y),
    .io_z(imm_switch_116_io_z),
    .io_in0(imm_switch_116_io_in0),
    .io_in1(imm_switch_116_io_in1),
    .io_sel0(imm_switch_116_io_sel0),
    .io_sel1(imm_switch_116_io_sel1)
  );
  Switch imm_switch_117 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_117_io_y),
    .io_z(imm_switch_117_io_z),
    .io_in0(imm_switch_117_io_in0),
    .io_in1(imm_switch_117_io_in1),
    .io_sel0(imm_switch_117_io_sel0),
    .io_sel1(imm_switch_117_io_sel1)
  );
  Switch imm_switch_118 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_118_io_y),
    .io_z(imm_switch_118_io_z),
    .io_in0(imm_switch_118_io_in0),
    .io_in1(imm_switch_118_io_in1),
    .io_sel0(imm_switch_118_io_sel0),
    .io_sel1(imm_switch_118_io_sel1)
  );
  Switch imm_switch_119 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_119_io_y),
    .io_z(imm_switch_119_io_z),
    .io_in0(imm_switch_119_io_in0),
    .io_in1(imm_switch_119_io_in1),
    .io_sel0(imm_switch_119_io_sel0),
    .io_sel1(imm_switch_119_io_sel1)
  );
  Switch imm_switch_120 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_120_io_y),
    .io_z(imm_switch_120_io_z),
    .io_in0(imm_switch_120_io_in0),
    .io_in1(imm_switch_120_io_in1),
    .io_sel0(imm_switch_120_io_sel0),
    .io_sel1(imm_switch_120_io_sel1)
  );
  Switch imm_switch_121 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_121_io_y),
    .io_z(imm_switch_121_io_z),
    .io_in0(imm_switch_121_io_in0),
    .io_in1(imm_switch_121_io_in1),
    .io_sel0(imm_switch_121_io_sel0),
    .io_sel1(imm_switch_121_io_sel1)
  );
  Switch imm_switch_122 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_122_io_y),
    .io_z(imm_switch_122_io_z),
    .io_in0(imm_switch_122_io_in0),
    .io_in1(imm_switch_122_io_in1),
    .io_sel0(imm_switch_122_io_sel0),
    .io_sel1(imm_switch_122_io_sel1)
  );
  Switch imm_switch_123 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_123_io_y),
    .io_z(imm_switch_123_io_z),
    .io_in0(imm_switch_123_io_in0),
    .io_in1(imm_switch_123_io_in1),
    .io_sel0(imm_switch_123_io_sel0),
    .io_sel1(imm_switch_123_io_sel1)
  );
  Switch imm_switch_124 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_124_io_y),
    .io_z(imm_switch_124_io_z),
    .io_in0(imm_switch_124_io_in0),
    .io_in1(imm_switch_124_io_in1),
    .io_sel0(imm_switch_124_io_sel0),
    .io_sel1(imm_switch_124_io_sel1)
  );
  Switch imm_switch_125 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_125_io_y),
    .io_z(imm_switch_125_io_z),
    .io_in0(imm_switch_125_io_in0),
    .io_in1(imm_switch_125_io_in1),
    .io_sel0(imm_switch_125_io_sel0),
    .io_sel1(imm_switch_125_io_sel1)
  );
  Switch imm_switch_126 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_126_io_y),
    .io_z(imm_switch_126_io_z),
    .io_in0(imm_switch_126_io_in0),
    .io_in1(imm_switch_126_io_in1),
    .io_sel0(imm_switch_126_io_sel0),
    .io_sel1(imm_switch_126_io_sel1)
  );
  Switch imm_switch_127 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_127_io_y),
    .io_z(imm_switch_127_io_z),
    .io_in0(imm_switch_127_io_in0),
    .io_in1(imm_switch_127_io_in1),
    .io_sel0(imm_switch_127_io_sel0),
    .io_sel1(imm_switch_127_io_sel1)
  );
  Switch imm_switch_128 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_128_io_y),
    .io_z(imm_switch_128_io_z),
    .io_in0(imm_switch_128_io_in0),
    .io_in1(imm_switch_128_io_in1),
    .io_sel0(imm_switch_128_io_sel0),
    .io_sel1(imm_switch_128_io_sel1)
  );
  Switch imm_switch_129 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_129_io_y),
    .io_z(imm_switch_129_io_z),
    .io_in0(imm_switch_129_io_in0),
    .io_in1(imm_switch_129_io_in1),
    .io_sel0(imm_switch_129_io_sel0),
    .io_sel1(imm_switch_129_io_sel1)
  );
  Switch imm_switch_130 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_130_io_y),
    .io_z(imm_switch_130_io_z),
    .io_in0(imm_switch_130_io_in0),
    .io_in1(imm_switch_130_io_in1),
    .io_sel0(imm_switch_130_io_sel0),
    .io_sel1(imm_switch_130_io_sel1)
  );
  Switch imm_switch_131 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_131_io_y),
    .io_z(imm_switch_131_io_z),
    .io_in0(imm_switch_131_io_in0),
    .io_in1(imm_switch_131_io_in1),
    .io_sel0(imm_switch_131_io_sel0),
    .io_sel1(imm_switch_131_io_sel1)
  );
  Switch imm_switch_132 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_132_io_y),
    .io_z(imm_switch_132_io_z),
    .io_in0(imm_switch_132_io_in0),
    .io_in1(imm_switch_132_io_in1),
    .io_sel0(imm_switch_132_io_sel0),
    .io_sel1(imm_switch_132_io_sel1)
  );
  Switch imm_switch_133 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_133_io_y),
    .io_z(imm_switch_133_io_z),
    .io_in0(imm_switch_133_io_in0),
    .io_in1(imm_switch_133_io_in1),
    .io_sel0(imm_switch_133_io_sel0),
    .io_sel1(imm_switch_133_io_sel1)
  );
  Switch imm_switch_134 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_134_io_y),
    .io_z(imm_switch_134_io_z),
    .io_in0(imm_switch_134_io_in0),
    .io_in1(imm_switch_134_io_in1),
    .io_sel0(imm_switch_134_io_sel0),
    .io_sel1(imm_switch_134_io_sel1)
  );
  Switch imm_switch_135 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_135_io_y),
    .io_z(imm_switch_135_io_z),
    .io_in0(imm_switch_135_io_in0),
    .io_in1(imm_switch_135_io_in1),
    .io_sel0(imm_switch_135_io_sel0),
    .io_sel1(imm_switch_135_io_sel1)
  );
  Switch imm_switch_136 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_136_io_y),
    .io_z(imm_switch_136_io_z),
    .io_in0(imm_switch_136_io_in0),
    .io_in1(imm_switch_136_io_in1),
    .io_sel0(imm_switch_136_io_sel0),
    .io_sel1(imm_switch_136_io_sel1)
  );
  Switch imm_switch_137 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_137_io_y),
    .io_z(imm_switch_137_io_z),
    .io_in0(imm_switch_137_io_in0),
    .io_in1(imm_switch_137_io_in1),
    .io_sel0(imm_switch_137_io_sel0),
    .io_sel1(imm_switch_137_io_sel1)
  );
  Switch imm_switch_138 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_138_io_y),
    .io_z(imm_switch_138_io_z),
    .io_in0(imm_switch_138_io_in0),
    .io_in1(imm_switch_138_io_in1),
    .io_sel0(imm_switch_138_io_sel0),
    .io_sel1(imm_switch_138_io_sel1)
  );
  Switch imm_switch_139 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_139_io_y),
    .io_z(imm_switch_139_io_z),
    .io_in0(imm_switch_139_io_in0),
    .io_in1(imm_switch_139_io_in1),
    .io_sel0(imm_switch_139_io_sel0),
    .io_sel1(imm_switch_139_io_sel1)
  );
  Switch imm_switch_140 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_140_io_y),
    .io_z(imm_switch_140_io_z),
    .io_in0(imm_switch_140_io_in0),
    .io_in1(imm_switch_140_io_in1),
    .io_sel0(imm_switch_140_io_sel0),
    .io_sel1(imm_switch_140_io_sel1)
  );
  Switch imm_switch_141 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_141_io_y),
    .io_z(imm_switch_141_io_z),
    .io_in0(imm_switch_141_io_in0),
    .io_in1(imm_switch_141_io_in1),
    .io_sel0(imm_switch_141_io_sel0),
    .io_sel1(imm_switch_141_io_sel1)
  );
  Switch imm_switch_142 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_142_io_y),
    .io_z(imm_switch_142_io_z),
    .io_in0(imm_switch_142_io_in0),
    .io_in1(imm_switch_142_io_in1),
    .io_sel0(imm_switch_142_io_sel0),
    .io_sel1(imm_switch_142_io_sel1)
  );
  Switch imm_switch_143 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_143_io_y),
    .io_z(imm_switch_143_io_z),
    .io_in0(imm_switch_143_io_in0),
    .io_in1(imm_switch_143_io_in1),
    .io_sel0(imm_switch_143_io_sel0),
    .io_sel1(imm_switch_143_io_sel1)
  );
  Switch imm_switch_144 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_144_io_y),
    .io_z(imm_switch_144_io_z),
    .io_in0(imm_switch_144_io_in0),
    .io_in1(imm_switch_144_io_in1),
    .io_sel0(imm_switch_144_io_sel0),
    .io_sel1(imm_switch_144_io_sel1)
  );
  Switch imm_switch_145 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_145_io_y),
    .io_z(imm_switch_145_io_z),
    .io_in0(imm_switch_145_io_in0),
    .io_in1(imm_switch_145_io_in1),
    .io_sel0(imm_switch_145_io_sel0),
    .io_sel1(imm_switch_145_io_sel1)
  );
  Switch imm_switch_146 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_146_io_y),
    .io_z(imm_switch_146_io_z),
    .io_in0(imm_switch_146_io_in0),
    .io_in1(imm_switch_146_io_in1),
    .io_sel0(imm_switch_146_io_sel0),
    .io_sel1(imm_switch_146_io_sel1)
  );
  Switch imm_switch_147 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_147_io_y),
    .io_z(imm_switch_147_io_z),
    .io_in0(imm_switch_147_io_in0),
    .io_in1(imm_switch_147_io_in1),
    .io_sel0(imm_switch_147_io_sel0),
    .io_sel1(imm_switch_147_io_sel1)
  );
  Switch imm_switch_148 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_148_io_y),
    .io_z(imm_switch_148_io_z),
    .io_in0(imm_switch_148_io_in0),
    .io_in1(imm_switch_148_io_in1),
    .io_sel0(imm_switch_148_io_sel0),
    .io_sel1(imm_switch_148_io_sel1)
  );
  Switch imm_switch_149 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_149_io_y),
    .io_z(imm_switch_149_io_z),
    .io_in0(imm_switch_149_io_in0),
    .io_in1(imm_switch_149_io_in1),
    .io_sel0(imm_switch_149_io_sel0),
    .io_sel1(imm_switch_149_io_sel1)
  );
  Switch imm_switch_150 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_150_io_y),
    .io_z(imm_switch_150_io_z),
    .io_in0(imm_switch_150_io_in0),
    .io_in1(imm_switch_150_io_in1),
    .io_sel0(imm_switch_150_io_sel0),
    .io_sel1(imm_switch_150_io_sel1)
  );
  Switch imm_switch_151 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_151_io_y),
    .io_z(imm_switch_151_io_z),
    .io_in0(imm_switch_151_io_in0),
    .io_in1(imm_switch_151_io_in1),
    .io_sel0(imm_switch_151_io_sel0),
    .io_sel1(imm_switch_151_io_sel1)
  );
  Switch imm_switch_152 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_152_io_y),
    .io_z(imm_switch_152_io_z),
    .io_in0(imm_switch_152_io_in0),
    .io_in1(imm_switch_152_io_in1),
    .io_sel0(imm_switch_152_io_sel0),
    .io_sel1(imm_switch_152_io_sel1)
  );
  Switch imm_switch_153 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_153_io_y),
    .io_z(imm_switch_153_io_z),
    .io_in0(imm_switch_153_io_in0),
    .io_in1(imm_switch_153_io_in1),
    .io_sel0(imm_switch_153_io_sel0),
    .io_sel1(imm_switch_153_io_sel1)
  );
  Switch imm_switch_154 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_154_io_y),
    .io_z(imm_switch_154_io_z),
    .io_in0(imm_switch_154_io_in0),
    .io_in1(imm_switch_154_io_in1),
    .io_sel0(imm_switch_154_io_sel0),
    .io_sel1(imm_switch_154_io_sel1)
  );
  Switch imm_switch_155 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_155_io_y),
    .io_z(imm_switch_155_io_z),
    .io_in0(imm_switch_155_io_in0),
    .io_in1(imm_switch_155_io_in1),
    .io_sel0(imm_switch_155_io_sel0),
    .io_sel1(imm_switch_155_io_sel1)
  );
  Switch imm_switch_156 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_156_io_y),
    .io_z(imm_switch_156_io_z),
    .io_in0(imm_switch_156_io_in0),
    .io_in1(imm_switch_156_io_in1),
    .io_sel0(imm_switch_156_io_sel0),
    .io_sel1(imm_switch_156_io_sel1)
  );
  Switch imm_switch_157 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_157_io_y),
    .io_z(imm_switch_157_io_z),
    .io_in0(imm_switch_157_io_in0),
    .io_in1(imm_switch_157_io_in1),
    .io_sel0(imm_switch_157_io_sel0),
    .io_sel1(imm_switch_157_io_sel1)
  );
  Switch imm_switch_158 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_158_io_y),
    .io_z(imm_switch_158_io_z),
    .io_in0(imm_switch_158_io_in0),
    .io_in1(imm_switch_158_io_in1),
    .io_sel0(imm_switch_158_io_sel0),
    .io_sel1(imm_switch_158_io_sel1)
  );
  Switch imm_switch_159 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_159_io_y),
    .io_z(imm_switch_159_io_z),
    .io_in0(imm_switch_159_io_in0),
    .io_in1(imm_switch_159_io_in1),
    .io_sel0(imm_switch_159_io_sel0),
    .io_sel1(imm_switch_159_io_sel1)
  );
  Switch imm_switch_160 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_160_io_y),
    .io_z(imm_switch_160_io_z),
    .io_in0(imm_switch_160_io_in0),
    .io_in1(imm_switch_160_io_in1),
    .io_sel0(imm_switch_160_io_sel0),
    .io_sel1(imm_switch_160_io_sel1)
  );
  Switch imm_switch_161 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_161_io_y),
    .io_z(imm_switch_161_io_z),
    .io_in0(imm_switch_161_io_in0),
    .io_in1(imm_switch_161_io_in1),
    .io_sel0(imm_switch_161_io_sel0),
    .io_sel1(imm_switch_161_io_sel1)
  );
  Switch imm_switch_162 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_162_io_y),
    .io_z(imm_switch_162_io_z),
    .io_in0(imm_switch_162_io_in0),
    .io_in1(imm_switch_162_io_in1),
    .io_sel0(imm_switch_162_io_sel0),
    .io_sel1(imm_switch_162_io_sel1)
  );
  Switch imm_switch_163 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_163_io_y),
    .io_z(imm_switch_163_io_z),
    .io_in0(imm_switch_163_io_in0),
    .io_in1(imm_switch_163_io_in1),
    .io_sel0(imm_switch_163_io_sel0),
    .io_sel1(imm_switch_163_io_sel1)
  );
  Switch imm_switch_164 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_164_io_y),
    .io_z(imm_switch_164_io_z),
    .io_in0(imm_switch_164_io_in0),
    .io_in1(imm_switch_164_io_in1),
    .io_sel0(imm_switch_164_io_sel0),
    .io_sel1(imm_switch_164_io_sel1)
  );
  Switch imm_switch_165 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_165_io_y),
    .io_z(imm_switch_165_io_z),
    .io_in0(imm_switch_165_io_in0),
    .io_in1(imm_switch_165_io_in1),
    .io_sel0(imm_switch_165_io_sel0),
    .io_sel1(imm_switch_165_io_sel1)
  );
  Switch imm_switch_166 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_166_io_y),
    .io_z(imm_switch_166_io_z),
    .io_in0(imm_switch_166_io_in0),
    .io_in1(imm_switch_166_io_in1),
    .io_sel0(imm_switch_166_io_sel0),
    .io_sel1(imm_switch_166_io_sel1)
  );
  Switch imm_switch_167 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_167_io_y),
    .io_z(imm_switch_167_io_z),
    .io_in0(imm_switch_167_io_in0),
    .io_in1(imm_switch_167_io_in1),
    .io_sel0(imm_switch_167_io_sel0),
    .io_sel1(imm_switch_167_io_sel1)
  );
  Switch imm_switch_168 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_168_io_y),
    .io_z(imm_switch_168_io_z),
    .io_in0(imm_switch_168_io_in0),
    .io_in1(imm_switch_168_io_in1),
    .io_sel0(imm_switch_168_io_sel0),
    .io_sel1(imm_switch_168_io_sel1)
  );
  Switch imm_switch_169 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_169_io_y),
    .io_z(imm_switch_169_io_z),
    .io_in0(imm_switch_169_io_in0),
    .io_in1(imm_switch_169_io_in1),
    .io_sel0(imm_switch_169_io_sel0),
    .io_sel1(imm_switch_169_io_sel1)
  );
  Switch imm_switch_170 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_170_io_y),
    .io_z(imm_switch_170_io_z),
    .io_in0(imm_switch_170_io_in0),
    .io_in1(imm_switch_170_io_in1),
    .io_sel0(imm_switch_170_io_sel0),
    .io_sel1(imm_switch_170_io_sel1)
  );
  Switch imm_switch_171 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_171_io_y),
    .io_z(imm_switch_171_io_z),
    .io_in0(imm_switch_171_io_in0),
    .io_in1(imm_switch_171_io_in1),
    .io_sel0(imm_switch_171_io_sel0),
    .io_sel1(imm_switch_171_io_sel1)
  );
  Switch imm_switch_172 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_172_io_y),
    .io_z(imm_switch_172_io_z),
    .io_in0(imm_switch_172_io_in0),
    .io_in1(imm_switch_172_io_in1),
    .io_sel0(imm_switch_172_io_sel0),
    .io_sel1(imm_switch_172_io_sel1)
  );
  Switch imm_switch_173 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_173_io_y),
    .io_z(imm_switch_173_io_z),
    .io_in0(imm_switch_173_io_in0),
    .io_in1(imm_switch_173_io_in1),
    .io_sel0(imm_switch_173_io_sel0),
    .io_sel1(imm_switch_173_io_sel1)
  );
  Switch imm_switch_174 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_174_io_y),
    .io_z(imm_switch_174_io_z),
    .io_in0(imm_switch_174_io_in0),
    .io_in1(imm_switch_174_io_in1),
    .io_sel0(imm_switch_174_io_sel0),
    .io_sel1(imm_switch_174_io_sel1)
  );
  Switch imm_switch_175 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_175_io_y),
    .io_z(imm_switch_175_io_z),
    .io_in0(imm_switch_175_io_in0),
    .io_in1(imm_switch_175_io_in1),
    .io_sel0(imm_switch_175_io_sel0),
    .io_sel1(imm_switch_175_io_sel1)
  );
  Switch imm_switch_176 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_176_io_y),
    .io_z(imm_switch_176_io_z),
    .io_in0(imm_switch_176_io_in0),
    .io_in1(imm_switch_176_io_in1),
    .io_sel0(imm_switch_176_io_sel0),
    .io_sel1(imm_switch_176_io_sel1)
  );
  Switch imm_switch_177 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_177_io_y),
    .io_z(imm_switch_177_io_z),
    .io_in0(imm_switch_177_io_in0),
    .io_in1(imm_switch_177_io_in1),
    .io_sel0(imm_switch_177_io_sel0),
    .io_sel1(imm_switch_177_io_sel1)
  );
  Switch imm_switch_178 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_178_io_y),
    .io_z(imm_switch_178_io_z),
    .io_in0(imm_switch_178_io_in0),
    .io_in1(imm_switch_178_io_in1),
    .io_sel0(imm_switch_178_io_sel0),
    .io_sel1(imm_switch_178_io_sel1)
  );
  Switch imm_switch_179 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_179_io_y),
    .io_z(imm_switch_179_io_z),
    .io_in0(imm_switch_179_io_in0),
    .io_in1(imm_switch_179_io_in1),
    .io_sel0(imm_switch_179_io_sel0),
    .io_sel1(imm_switch_179_io_sel1)
  );
  Switch imm_switch_180 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_180_io_y),
    .io_z(imm_switch_180_io_z),
    .io_in0(imm_switch_180_io_in0),
    .io_in1(imm_switch_180_io_in1),
    .io_sel0(imm_switch_180_io_sel0),
    .io_sel1(imm_switch_180_io_sel1)
  );
  Switch imm_switch_181 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_181_io_y),
    .io_z(imm_switch_181_io_z),
    .io_in0(imm_switch_181_io_in0),
    .io_in1(imm_switch_181_io_in1),
    .io_sel0(imm_switch_181_io_sel0),
    .io_sel1(imm_switch_181_io_sel1)
  );
  Switch imm_switch_182 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_182_io_y),
    .io_z(imm_switch_182_io_z),
    .io_in0(imm_switch_182_io_in0),
    .io_in1(imm_switch_182_io_in1),
    .io_sel0(imm_switch_182_io_sel0),
    .io_sel1(imm_switch_182_io_sel1)
  );
  Switch imm_switch_183 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_183_io_y),
    .io_z(imm_switch_183_io_z),
    .io_in0(imm_switch_183_io_in0),
    .io_in1(imm_switch_183_io_in1),
    .io_sel0(imm_switch_183_io_sel0),
    .io_sel1(imm_switch_183_io_sel1)
  );
  Switch imm_switch_184 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_184_io_y),
    .io_z(imm_switch_184_io_z),
    .io_in0(imm_switch_184_io_in0),
    .io_in1(imm_switch_184_io_in1),
    .io_sel0(imm_switch_184_io_sel0),
    .io_sel1(imm_switch_184_io_sel1)
  );
  Switch imm_switch_185 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_185_io_y),
    .io_z(imm_switch_185_io_z),
    .io_in0(imm_switch_185_io_in0),
    .io_in1(imm_switch_185_io_in1),
    .io_sel0(imm_switch_185_io_sel0),
    .io_sel1(imm_switch_185_io_sel1)
  );
  Switch imm_switch_186 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_186_io_y),
    .io_z(imm_switch_186_io_z),
    .io_in0(imm_switch_186_io_in0),
    .io_in1(imm_switch_186_io_in1),
    .io_sel0(imm_switch_186_io_sel0),
    .io_sel1(imm_switch_186_io_sel1)
  );
  Switch imm_switch_187 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_187_io_y),
    .io_z(imm_switch_187_io_z),
    .io_in0(imm_switch_187_io_in0),
    .io_in1(imm_switch_187_io_in1),
    .io_sel0(imm_switch_187_io_sel0),
    .io_sel1(imm_switch_187_io_sel1)
  );
  Switch imm_switch_188 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_188_io_y),
    .io_z(imm_switch_188_io_z),
    .io_in0(imm_switch_188_io_in0),
    .io_in1(imm_switch_188_io_in1),
    .io_sel0(imm_switch_188_io_sel0),
    .io_sel1(imm_switch_188_io_sel1)
  );
  Switch imm_switch_189 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_189_io_y),
    .io_z(imm_switch_189_io_z),
    .io_in0(imm_switch_189_io_in0),
    .io_in1(imm_switch_189_io_in1),
    .io_sel0(imm_switch_189_io_sel0),
    .io_sel1(imm_switch_189_io_sel1)
  );
  Switch imm_switch_190 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_190_io_y),
    .io_z(imm_switch_190_io_z),
    .io_in0(imm_switch_190_io_in0),
    .io_in1(imm_switch_190_io_in1),
    .io_sel0(imm_switch_190_io_sel0),
    .io_sel1(imm_switch_190_io_sel1)
  );
  Switch imm_switch_191 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_191_io_y),
    .io_z(imm_switch_191_io_z),
    .io_in0(imm_switch_191_io_in0),
    .io_in1(imm_switch_191_io_in1),
    .io_sel0(imm_switch_191_io_sel0),
    .io_sel1(imm_switch_191_io_sel1)
  );
  Switch imm_switch_192 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_192_io_y),
    .io_z(imm_switch_192_io_z),
    .io_in0(imm_switch_192_io_in0),
    .io_in1(imm_switch_192_io_in1),
    .io_sel0(imm_switch_192_io_sel0),
    .io_sel1(imm_switch_192_io_sel1)
  );
  Switch imm_switch_193 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_193_io_y),
    .io_z(imm_switch_193_io_z),
    .io_in0(imm_switch_193_io_in0),
    .io_in1(imm_switch_193_io_in1),
    .io_sel0(imm_switch_193_io_sel0),
    .io_sel1(imm_switch_193_io_sel1)
  );
  Switch imm_switch_194 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_194_io_y),
    .io_z(imm_switch_194_io_z),
    .io_in0(imm_switch_194_io_in0),
    .io_in1(imm_switch_194_io_in1),
    .io_sel0(imm_switch_194_io_sel0),
    .io_sel1(imm_switch_194_io_sel1)
  );
  Switch imm_switch_195 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_195_io_y),
    .io_z(imm_switch_195_io_z),
    .io_in0(imm_switch_195_io_in0),
    .io_in1(imm_switch_195_io_in1),
    .io_sel0(imm_switch_195_io_sel0),
    .io_sel1(imm_switch_195_io_sel1)
  );
  Switch imm_switch_196 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_196_io_y),
    .io_z(imm_switch_196_io_z),
    .io_in0(imm_switch_196_io_in0),
    .io_in1(imm_switch_196_io_in1),
    .io_sel0(imm_switch_196_io_sel0),
    .io_sel1(imm_switch_196_io_sel1)
  );
  Switch imm_switch_197 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_197_io_y),
    .io_z(imm_switch_197_io_z),
    .io_in0(imm_switch_197_io_in0),
    .io_in1(imm_switch_197_io_in1),
    .io_sel0(imm_switch_197_io_sel0),
    .io_sel1(imm_switch_197_io_sel1)
  );
  Switch imm_switch_198 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_198_io_y),
    .io_z(imm_switch_198_io_z),
    .io_in0(imm_switch_198_io_in0),
    .io_in1(imm_switch_198_io_in1),
    .io_sel0(imm_switch_198_io_sel0),
    .io_sel1(imm_switch_198_io_sel1)
  );
  Switch imm_switch_199 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_199_io_y),
    .io_z(imm_switch_199_io_z),
    .io_in0(imm_switch_199_io_in0),
    .io_in1(imm_switch_199_io_in1),
    .io_sel0(imm_switch_199_io_sel0),
    .io_sel1(imm_switch_199_io_sel1)
  );
  Switch imm_switch_200 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_200_io_y),
    .io_z(imm_switch_200_io_z),
    .io_in0(imm_switch_200_io_in0),
    .io_in1(imm_switch_200_io_in1),
    .io_sel0(imm_switch_200_io_sel0),
    .io_sel1(imm_switch_200_io_sel1)
  );
  Switch imm_switch_201 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_201_io_y),
    .io_z(imm_switch_201_io_z),
    .io_in0(imm_switch_201_io_in0),
    .io_in1(imm_switch_201_io_in1),
    .io_sel0(imm_switch_201_io_sel0),
    .io_sel1(imm_switch_201_io_sel1)
  );
  Switch imm_switch_202 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_202_io_y),
    .io_z(imm_switch_202_io_z),
    .io_in0(imm_switch_202_io_in0),
    .io_in1(imm_switch_202_io_in1),
    .io_sel0(imm_switch_202_io_sel0),
    .io_sel1(imm_switch_202_io_sel1)
  );
  Switch imm_switch_203 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_203_io_y),
    .io_z(imm_switch_203_io_z),
    .io_in0(imm_switch_203_io_in0),
    .io_in1(imm_switch_203_io_in1),
    .io_sel0(imm_switch_203_io_sel0),
    .io_sel1(imm_switch_203_io_sel1)
  );
  Switch imm_switch_204 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_204_io_y),
    .io_z(imm_switch_204_io_z),
    .io_in0(imm_switch_204_io_in0),
    .io_in1(imm_switch_204_io_in1),
    .io_sel0(imm_switch_204_io_sel0),
    .io_sel1(imm_switch_204_io_sel1)
  );
  Switch imm_switch_205 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_205_io_y),
    .io_z(imm_switch_205_io_z),
    .io_in0(imm_switch_205_io_in0),
    .io_in1(imm_switch_205_io_in1),
    .io_sel0(imm_switch_205_io_sel0),
    .io_sel1(imm_switch_205_io_sel1)
  );
  Switch imm_switch_206 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_206_io_y),
    .io_z(imm_switch_206_io_z),
    .io_in0(imm_switch_206_io_in0),
    .io_in1(imm_switch_206_io_in1),
    .io_sel0(imm_switch_206_io_sel0),
    .io_sel1(imm_switch_206_io_sel1)
  );
  Switch imm_switch_207 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_207_io_y),
    .io_z(imm_switch_207_io_z),
    .io_in0(imm_switch_207_io_in0),
    .io_in1(imm_switch_207_io_in1),
    .io_sel0(imm_switch_207_io_sel0),
    .io_sel1(imm_switch_207_io_sel1)
  );
  Switch imm_switch_208 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_208_io_y),
    .io_z(imm_switch_208_io_z),
    .io_in0(imm_switch_208_io_in0),
    .io_in1(imm_switch_208_io_in1),
    .io_sel0(imm_switch_208_io_sel0),
    .io_sel1(imm_switch_208_io_sel1)
  );
  Switch imm_switch_209 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_209_io_y),
    .io_z(imm_switch_209_io_z),
    .io_in0(imm_switch_209_io_in0),
    .io_in1(imm_switch_209_io_in1),
    .io_sel0(imm_switch_209_io_sel0),
    .io_sel1(imm_switch_209_io_sel1)
  );
  Switch imm_switch_210 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_210_io_y),
    .io_z(imm_switch_210_io_z),
    .io_in0(imm_switch_210_io_in0),
    .io_in1(imm_switch_210_io_in1),
    .io_sel0(imm_switch_210_io_sel0),
    .io_sel1(imm_switch_210_io_sel1)
  );
  Switch imm_switch_211 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_211_io_y),
    .io_z(imm_switch_211_io_z),
    .io_in0(imm_switch_211_io_in0),
    .io_in1(imm_switch_211_io_in1),
    .io_sel0(imm_switch_211_io_sel0),
    .io_sel1(imm_switch_211_io_sel1)
  );
  Switch imm_switch_212 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_212_io_y),
    .io_z(imm_switch_212_io_z),
    .io_in0(imm_switch_212_io_in0),
    .io_in1(imm_switch_212_io_in1),
    .io_sel0(imm_switch_212_io_sel0),
    .io_sel1(imm_switch_212_io_sel1)
  );
  Switch imm_switch_213 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_213_io_y),
    .io_z(imm_switch_213_io_z),
    .io_in0(imm_switch_213_io_in0),
    .io_in1(imm_switch_213_io_in1),
    .io_sel0(imm_switch_213_io_sel0),
    .io_sel1(imm_switch_213_io_sel1)
  );
  Switch imm_switch_214 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_214_io_y),
    .io_z(imm_switch_214_io_z),
    .io_in0(imm_switch_214_io_in0),
    .io_in1(imm_switch_214_io_in1),
    .io_sel0(imm_switch_214_io_sel0),
    .io_sel1(imm_switch_214_io_sel1)
  );
  Switch imm_switch_215 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_215_io_y),
    .io_z(imm_switch_215_io_z),
    .io_in0(imm_switch_215_io_in0),
    .io_in1(imm_switch_215_io_in1),
    .io_sel0(imm_switch_215_io_sel0),
    .io_sel1(imm_switch_215_io_sel1)
  );
  Switch imm_switch_216 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_216_io_y),
    .io_z(imm_switch_216_io_z),
    .io_in0(imm_switch_216_io_in0),
    .io_in1(imm_switch_216_io_in1),
    .io_sel0(imm_switch_216_io_sel0),
    .io_sel1(imm_switch_216_io_sel1)
  );
  Switch imm_switch_217 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_217_io_y),
    .io_z(imm_switch_217_io_z),
    .io_in0(imm_switch_217_io_in0),
    .io_in1(imm_switch_217_io_in1),
    .io_sel0(imm_switch_217_io_sel0),
    .io_sel1(imm_switch_217_io_sel1)
  );
  Switch imm_switch_218 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_218_io_y),
    .io_z(imm_switch_218_io_z),
    .io_in0(imm_switch_218_io_in0),
    .io_in1(imm_switch_218_io_in1),
    .io_sel0(imm_switch_218_io_sel0),
    .io_sel1(imm_switch_218_io_sel1)
  );
  Switch imm_switch_219 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_219_io_y),
    .io_z(imm_switch_219_io_z),
    .io_in0(imm_switch_219_io_in0),
    .io_in1(imm_switch_219_io_in1),
    .io_sel0(imm_switch_219_io_sel0),
    .io_sel1(imm_switch_219_io_sel1)
  );
  Switch imm_switch_220 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_220_io_y),
    .io_z(imm_switch_220_io_z),
    .io_in0(imm_switch_220_io_in0),
    .io_in1(imm_switch_220_io_in1),
    .io_sel0(imm_switch_220_io_sel0),
    .io_sel1(imm_switch_220_io_sel1)
  );
  Switch imm_switch_221 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_221_io_y),
    .io_z(imm_switch_221_io_z),
    .io_in0(imm_switch_221_io_in0),
    .io_in1(imm_switch_221_io_in1),
    .io_sel0(imm_switch_221_io_sel0),
    .io_sel1(imm_switch_221_io_sel1)
  );
  Switch imm_switch_222 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_222_io_y),
    .io_z(imm_switch_222_io_z),
    .io_in0(imm_switch_222_io_in0),
    .io_in1(imm_switch_222_io_in1),
    .io_sel0(imm_switch_222_io_sel0),
    .io_sel1(imm_switch_222_io_sel1)
  );
  Switch imm_switch_223 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_223_io_y),
    .io_z(imm_switch_223_io_z),
    .io_in0(imm_switch_223_io_in0),
    .io_in1(imm_switch_223_io_in1),
    .io_sel0(imm_switch_223_io_sel0),
    .io_sel1(imm_switch_223_io_sel1)
  );
  Switch imm_switch_224 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_224_io_y),
    .io_z(imm_switch_224_io_z),
    .io_in0(imm_switch_224_io_in0),
    .io_in1(imm_switch_224_io_in1),
    .io_sel0(imm_switch_224_io_sel0),
    .io_sel1(imm_switch_224_io_sel1)
  );
  Switch imm_switch_225 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_225_io_y),
    .io_z(imm_switch_225_io_z),
    .io_in0(imm_switch_225_io_in0),
    .io_in1(imm_switch_225_io_in1),
    .io_sel0(imm_switch_225_io_sel0),
    .io_sel1(imm_switch_225_io_sel1)
  );
  Switch imm_switch_226 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_226_io_y),
    .io_z(imm_switch_226_io_z),
    .io_in0(imm_switch_226_io_in0),
    .io_in1(imm_switch_226_io_in1),
    .io_sel0(imm_switch_226_io_sel0),
    .io_sel1(imm_switch_226_io_sel1)
  );
  Switch imm_switch_227 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_227_io_y),
    .io_z(imm_switch_227_io_z),
    .io_in0(imm_switch_227_io_in0),
    .io_in1(imm_switch_227_io_in1),
    .io_sel0(imm_switch_227_io_sel0),
    .io_sel1(imm_switch_227_io_sel1)
  );
  Switch imm_switch_228 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_228_io_y),
    .io_z(imm_switch_228_io_z),
    .io_in0(imm_switch_228_io_in0),
    .io_in1(imm_switch_228_io_in1),
    .io_sel0(imm_switch_228_io_sel0),
    .io_sel1(imm_switch_228_io_sel1)
  );
  Switch imm_switch_229 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_229_io_y),
    .io_z(imm_switch_229_io_z),
    .io_in0(imm_switch_229_io_in0),
    .io_in1(imm_switch_229_io_in1),
    .io_sel0(imm_switch_229_io_sel0),
    .io_sel1(imm_switch_229_io_sel1)
  );
  Switch imm_switch_230 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_230_io_y),
    .io_z(imm_switch_230_io_z),
    .io_in0(imm_switch_230_io_in0),
    .io_in1(imm_switch_230_io_in1),
    .io_sel0(imm_switch_230_io_sel0),
    .io_sel1(imm_switch_230_io_sel1)
  );
  Switch imm_switch_231 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_231_io_y),
    .io_z(imm_switch_231_io_z),
    .io_in0(imm_switch_231_io_in0),
    .io_in1(imm_switch_231_io_in1),
    .io_sel0(imm_switch_231_io_sel0),
    .io_sel1(imm_switch_231_io_sel1)
  );
  Switch imm_switch_232 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_232_io_y),
    .io_z(imm_switch_232_io_z),
    .io_in0(imm_switch_232_io_in0),
    .io_in1(imm_switch_232_io_in1),
    .io_sel0(imm_switch_232_io_sel0),
    .io_sel1(imm_switch_232_io_sel1)
  );
  Switch imm_switch_233 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_233_io_y),
    .io_z(imm_switch_233_io_z),
    .io_in0(imm_switch_233_io_in0),
    .io_in1(imm_switch_233_io_in1),
    .io_sel0(imm_switch_233_io_sel0),
    .io_sel1(imm_switch_233_io_sel1)
  );
  Switch imm_switch_234 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_234_io_y),
    .io_z(imm_switch_234_io_z),
    .io_in0(imm_switch_234_io_in0),
    .io_in1(imm_switch_234_io_in1),
    .io_sel0(imm_switch_234_io_sel0),
    .io_sel1(imm_switch_234_io_sel1)
  );
  Switch imm_switch_235 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_235_io_y),
    .io_z(imm_switch_235_io_z),
    .io_in0(imm_switch_235_io_in0),
    .io_in1(imm_switch_235_io_in1),
    .io_sel0(imm_switch_235_io_sel0),
    .io_sel1(imm_switch_235_io_sel1)
  );
  Switch imm_switch_236 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_236_io_y),
    .io_z(imm_switch_236_io_z),
    .io_in0(imm_switch_236_io_in0),
    .io_in1(imm_switch_236_io_in1),
    .io_sel0(imm_switch_236_io_sel0),
    .io_sel1(imm_switch_236_io_sel1)
  );
  Switch imm_switch_237 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_237_io_y),
    .io_z(imm_switch_237_io_z),
    .io_in0(imm_switch_237_io_in0),
    .io_in1(imm_switch_237_io_in1),
    .io_sel0(imm_switch_237_io_sel0),
    .io_sel1(imm_switch_237_io_sel1)
  );
  Switch imm_switch_238 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_238_io_y),
    .io_z(imm_switch_238_io_z),
    .io_in0(imm_switch_238_io_in0),
    .io_in1(imm_switch_238_io_in1),
    .io_sel0(imm_switch_238_io_sel0),
    .io_sel1(imm_switch_238_io_sel1)
  );
  Switch imm_switch_239 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_239_io_y),
    .io_z(imm_switch_239_io_z),
    .io_in0(imm_switch_239_io_in0),
    .io_in1(imm_switch_239_io_in1),
    .io_sel0(imm_switch_239_io_sel0),
    .io_sel1(imm_switch_239_io_sel1)
  );
  Switch imm_switch_240 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_240_io_y),
    .io_z(imm_switch_240_io_z),
    .io_in0(imm_switch_240_io_in0),
    .io_in1(imm_switch_240_io_in1),
    .io_sel0(imm_switch_240_io_sel0),
    .io_sel1(imm_switch_240_io_sel1)
  );
  Switch imm_switch_241 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_241_io_y),
    .io_z(imm_switch_241_io_z),
    .io_in0(imm_switch_241_io_in0),
    .io_in1(imm_switch_241_io_in1),
    .io_sel0(imm_switch_241_io_sel0),
    .io_sel1(imm_switch_241_io_sel1)
  );
  Switch imm_switch_242 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_242_io_y),
    .io_z(imm_switch_242_io_z),
    .io_in0(imm_switch_242_io_in0),
    .io_in1(imm_switch_242_io_in1),
    .io_sel0(imm_switch_242_io_sel0),
    .io_sel1(imm_switch_242_io_sel1)
  );
  Switch imm_switch_243 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_243_io_y),
    .io_z(imm_switch_243_io_z),
    .io_in0(imm_switch_243_io_in0),
    .io_in1(imm_switch_243_io_in1),
    .io_sel0(imm_switch_243_io_sel0),
    .io_sel1(imm_switch_243_io_sel1)
  );
  Switch imm_switch_244 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_244_io_y),
    .io_z(imm_switch_244_io_z),
    .io_in0(imm_switch_244_io_in0),
    .io_in1(imm_switch_244_io_in1),
    .io_sel0(imm_switch_244_io_sel0),
    .io_sel1(imm_switch_244_io_sel1)
  );
  Switch imm_switch_245 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_245_io_y),
    .io_z(imm_switch_245_io_z),
    .io_in0(imm_switch_245_io_in0),
    .io_in1(imm_switch_245_io_in1),
    .io_sel0(imm_switch_245_io_sel0),
    .io_sel1(imm_switch_245_io_sel1)
  );
  Switch imm_switch_246 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_246_io_y),
    .io_z(imm_switch_246_io_z),
    .io_in0(imm_switch_246_io_in0),
    .io_in1(imm_switch_246_io_in1),
    .io_sel0(imm_switch_246_io_sel0),
    .io_sel1(imm_switch_246_io_sel1)
  );
  Switch imm_switch_247 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_247_io_y),
    .io_z(imm_switch_247_io_z),
    .io_in0(imm_switch_247_io_in0),
    .io_in1(imm_switch_247_io_in1),
    .io_sel0(imm_switch_247_io_sel0),
    .io_sel1(imm_switch_247_io_sel1)
  );
  Switch imm_switch_248 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_248_io_y),
    .io_z(imm_switch_248_io_z),
    .io_in0(imm_switch_248_io_in0),
    .io_in1(imm_switch_248_io_in1),
    .io_sel0(imm_switch_248_io_sel0),
    .io_sel1(imm_switch_248_io_sel1)
  );
  Switch imm_switch_249 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_249_io_y),
    .io_z(imm_switch_249_io_z),
    .io_in0(imm_switch_249_io_in0),
    .io_in1(imm_switch_249_io_in1),
    .io_sel0(imm_switch_249_io_sel0),
    .io_sel1(imm_switch_249_io_sel1)
  );
  Switch imm_switch_250 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_250_io_y),
    .io_z(imm_switch_250_io_z),
    .io_in0(imm_switch_250_io_in0),
    .io_in1(imm_switch_250_io_in1),
    .io_sel0(imm_switch_250_io_sel0),
    .io_sel1(imm_switch_250_io_sel1)
  );
  Switch imm_switch_251 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_251_io_y),
    .io_z(imm_switch_251_io_z),
    .io_in0(imm_switch_251_io_in0),
    .io_in1(imm_switch_251_io_in1),
    .io_sel0(imm_switch_251_io_sel0),
    .io_sel1(imm_switch_251_io_sel1)
  );
  Switch imm_switch_252 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_252_io_y),
    .io_z(imm_switch_252_io_z),
    .io_in0(imm_switch_252_io_in0),
    .io_in1(imm_switch_252_io_in1),
    .io_sel0(imm_switch_252_io_sel0),
    .io_sel1(imm_switch_252_io_sel1)
  );
  Switch imm_switch_253 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_253_io_y),
    .io_z(imm_switch_253_io_z),
    .io_in0(imm_switch_253_io_in0),
    .io_in1(imm_switch_253_io_in1),
    .io_sel0(imm_switch_253_io_sel0),
    .io_sel1(imm_switch_253_io_sel1)
  );
  Switch imm_switch_254 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_254_io_y),
    .io_z(imm_switch_254_io_z),
    .io_in0(imm_switch_254_io_in0),
    .io_in1(imm_switch_254_io_in1),
    .io_sel0(imm_switch_254_io_sel0),
    .io_sel1(imm_switch_254_io_sel1)
  );
  Switch imm_switch_255 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_255_io_y),
    .io_z(imm_switch_255_io_z),
    .io_in0(imm_switch_255_io_in0),
    .io_in1(imm_switch_255_io_in1),
    .io_sel0(imm_switch_255_io_sel0),
    .io_sel1(imm_switch_255_io_sel1)
  );
  Switch imm_switch_256 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_256_io_y),
    .io_z(imm_switch_256_io_z),
    .io_in0(imm_switch_256_io_in0),
    .io_in1(imm_switch_256_io_in1),
    .io_sel0(imm_switch_256_io_sel0),
    .io_sel1(imm_switch_256_io_sel1)
  );
  Switch imm_switch_257 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_257_io_y),
    .io_z(imm_switch_257_io_z),
    .io_in0(imm_switch_257_io_in0),
    .io_in1(imm_switch_257_io_in1),
    .io_sel0(imm_switch_257_io_sel0),
    .io_sel1(imm_switch_257_io_sel1)
  );
  Switch imm_switch_258 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_258_io_y),
    .io_z(imm_switch_258_io_z),
    .io_in0(imm_switch_258_io_in0),
    .io_in1(imm_switch_258_io_in1),
    .io_sel0(imm_switch_258_io_sel0),
    .io_sel1(imm_switch_258_io_sel1)
  );
  Switch imm_switch_259 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_259_io_y),
    .io_z(imm_switch_259_io_z),
    .io_in0(imm_switch_259_io_in0),
    .io_in1(imm_switch_259_io_in1),
    .io_sel0(imm_switch_259_io_sel0),
    .io_sel1(imm_switch_259_io_sel1)
  );
  Switch imm_switch_260 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_260_io_y),
    .io_z(imm_switch_260_io_z),
    .io_in0(imm_switch_260_io_in0),
    .io_in1(imm_switch_260_io_in1),
    .io_sel0(imm_switch_260_io_sel0),
    .io_sel1(imm_switch_260_io_sel1)
  );
  Switch imm_switch_261 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_261_io_y),
    .io_z(imm_switch_261_io_z),
    .io_in0(imm_switch_261_io_in0),
    .io_in1(imm_switch_261_io_in1),
    .io_sel0(imm_switch_261_io_sel0),
    .io_sel1(imm_switch_261_io_sel1)
  );
  Switch imm_switch_262 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_262_io_y),
    .io_z(imm_switch_262_io_z),
    .io_in0(imm_switch_262_io_in0),
    .io_in1(imm_switch_262_io_in1),
    .io_sel0(imm_switch_262_io_sel0),
    .io_sel1(imm_switch_262_io_sel1)
  );
  Switch imm_switch_263 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_263_io_y),
    .io_z(imm_switch_263_io_z),
    .io_in0(imm_switch_263_io_in0),
    .io_in1(imm_switch_263_io_in1),
    .io_sel0(imm_switch_263_io_sel0),
    .io_sel1(imm_switch_263_io_sel1)
  );
  Switch imm_switch_264 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_264_io_y),
    .io_z(imm_switch_264_io_z),
    .io_in0(imm_switch_264_io_in0),
    .io_in1(imm_switch_264_io_in1),
    .io_sel0(imm_switch_264_io_sel0),
    .io_sel1(imm_switch_264_io_sel1)
  );
  Switch imm_switch_265 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_265_io_y),
    .io_z(imm_switch_265_io_z),
    .io_in0(imm_switch_265_io_in0),
    .io_in1(imm_switch_265_io_in1),
    .io_sel0(imm_switch_265_io_sel0),
    .io_sel1(imm_switch_265_io_sel1)
  );
  Switch imm_switch_266 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_266_io_y),
    .io_z(imm_switch_266_io_z),
    .io_in0(imm_switch_266_io_in0),
    .io_in1(imm_switch_266_io_in1),
    .io_sel0(imm_switch_266_io_sel0),
    .io_sel1(imm_switch_266_io_sel1)
  );
  Switch imm_switch_267 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_267_io_y),
    .io_z(imm_switch_267_io_z),
    .io_in0(imm_switch_267_io_in0),
    .io_in1(imm_switch_267_io_in1),
    .io_sel0(imm_switch_267_io_sel0),
    .io_sel1(imm_switch_267_io_sel1)
  );
  Switch imm_switch_268 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_268_io_y),
    .io_z(imm_switch_268_io_z),
    .io_in0(imm_switch_268_io_in0),
    .io_in1(imm_switch_268_io_in1),
    .io_sel0(imm_switch_268_io_sel0),
    .io_sel1(imm_switch_268_io_sel1)
  );
  Switch imm_switch_269 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_269_io_y),
    .io_z(imm_switch_269_io_z),
    .io_in0(imm_switch_269_io_in0),
    .io_in1(imm_switch_269_io_in1),
    .io_sel0(imm_switch_269_io_sel0),
    .io_sel1(imm_switch_269_io_sel1)
  );
  Switch imm_switch_270 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_270_io_y),
    .io_z(imm_switch_270_io_z),
    .io_in0(imm_switch_270_io_in0),
    .io_in1(imm_switch_270_io_in1),
    .io_sel0(imm_switch_270_io_sel0),
    .io_sel1(imm_switch_270_io_sel1)
  );
  Switch imm_switch_271 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_271_io_y),
    .io_z(imm_switch_271_io_z),
    .io_in0(imm_switch_271_io_in0),
    .io_in1(imm_switch_271_io_in1),
    .io_sel0(imm_switch_271_io_sel0),
    .io_sel1(imm_switch_271_io_sel1)
  );
  Switch imm_switch_272 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_272_io_y),
    .io_z(imm_switch_272_io_z),
    .io_in0(imm_switch_272_io_in0),
    .io_in1(imm_switch_272_io_in1),
    .io_sel0(imm_switch_272_io_sel0),
    .io_sel1(imm_switch_272_io_sel1)
  );
  Switch imm_switch_273 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_273_io_y),
    .io_z(imm_switch_273_io_z),
    .io_in0(imm_switch_273_io_in0),
    .io_in1(imm_switch_273_io_in1),
    .io_sel0(imm_switch_273_io_sel0),
    .io_sel1(imm_switch_273_io_sel1)
  );
  Switch imm_switch_274 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_274_io_y),
    .io_z(imm_switch_274_io_z),
    .io_in0(imm_switch_274_io_in0),
    .io_in1(imm_switch_274_io_in1),
    .io_sel0(imm_switch_274_io_sel0),
    .io_sel1(imm_switch_274_io_sel1)
  );
  Switch imm_switch_275 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_275_io_y),
    .io_z(imm_switch_275_io_z),
    .io_in0(imm_switch_275_io_in0),
    .io_in1(imm_switch_275_io_in1),
    .io_sel0(imm_switch_275_io_sel0),
    .io_sel1(imm_switch_275_io_sel1)
  );
  Switch imm_switch_276 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_276_io_y),
    .io_z(imm_switch_276_io_z),
    .io_in0(imm_switch_276_io_in0),
    .io_in1(imm_switch_276_io_in1),
    .io_sel0(imm_switch_276_io_sel0),
    .io_sel1(imm_switch_276_io_sel1)
  );
  Switch imm_switch_277 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_277_io_y),
    .io_z(imm_switch_277_io_z),
    .io_in0(imm_switch_277_io_in0),
    .io_in1(imm_switch_277_io_in1),
    .io_sel0(imm_switch_277_io_sel0),
    .io_sel1(imm_switch_277_io_sel1)
  );
  Switch imm_switch_278 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_278_io_y),
    .io_z(imm_switch_278_io_z),
    .io_in0(imm_switch_278_io_in0),
    .io_in1(imm_switch_278_io_in1),
    .io_sel0(imm_switch_278_io_sel0),
    .io_sel1(imm_switch_278_io_sel1)
  );
  Switch imm_switch_279 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_279_io_y),
    .io_z(imm_switch_279_io_z),
    .io_in0(imm_switch_279_io_in0),
    .io_in1(imm_switch_279_io_in1),
    .io_sel0(imm_switch_279_io_sel0),
    .io_sel1(imm_switch_279_io_sel1)
  );
  Switch imm_switch_280 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_280_io_y),
    .io_z(imm_switch_280_io_z),
    .io_in0(imm_switch_280_io_in0),
    .io_in1(imm_switch_280_io_in1),
    .io_sel0(imm_switch_280_io_sel0),
    .io_sel1(imm_switch_280_io_sel1)
  );
  Switch imm_switch_281 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_281_io_y),
    .io_z(imm_switch_281_io_z),
    .io_in0(imm_switch_281_io_in0),
    .io_in1(imm_switch_281_io_in1),
    .io_sel0(imm_switch_281_io_sel0),
    .io_sel1(imm_switch_281_io_sel1)
  );
  Switch imm_switch_282 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_282_io_y),
    .io_z(imm_switch_282_io_z),
    .io_in0(imm_switch_282_io_in0),
    .io_in1(imm_switch_282_io_in1),
    .io_sel0(imm_switch_282_io_sel0),
    .io_sel1(imm_switch_282_io_sel1)
  );
  Switch imm_switch_283 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_283_io_y),
    .io_z(imm_switch_283_io_z),
    .io_in0(imm_switch_283_io_in0),
    .io_in1(imm_switch_283_io_in1),
    .io_sel0(imm_switch_283_io_sel0),
    .io_sel1(imm_switch_283_io_sel1)
  );
  Switch imm_switch_284 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_284_io_y),
    .io_z(imm_switch_284_io_z),
    .io_in0(imm_switch_284_io_in0),
    .io_in1(imm_switch_284_io_in1),
    .io_sel0(imm_switch_284_io_sel0),
    .io_sel1(imm_switch_284_io_sel1)
  );
  Switch imm_switch_285 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_285_io_y),
    .io_z(imm_switch_285_io_z),
    .io_in0(imm_switch_285_io_in0),
    .io_in1(imm_switch_285_io_in1),
    .io_sel0(imm_switch_285_io_sel0),
    .io_sel1(imm_switch_285_io_sel1)
  );
  Switch imm_switch_286 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_286_io_y),
    .io_z(imm_switch_286_io_z),
    .io_in0(imm_switch_286_io_in0),
    .io_in1(imm_switch_286_io_in1),
    .io_sel0(imm_switch_286_io_sel0),
    .io_sel1(imm_switch_286_io_sel1)
  );
  Switch imm_switch_287 ( // @[Benes.scala 108:30]
    .io_y(imm_switch_287_io_y),
    .io_z(imm_switch_287_io_z),
    .io_in0(imm_switch_287_io_in0),
    .io_in1(imm_switch_287_io_in1),
    .io_sel0(imm_switch_287_io_sel0),
    .io_sel1(imm_switch_287_io_sel1)
  );
  assign io_o_dist_bus_0 = reset ? 32'h0 : w_dist_bus_0; // @[Benes.scala 85:23]
  assign io_o_dist_bus_1 = reset ? 32'h0 : w_dist_bus_1; // @[Benes.scala 85:23]
  assign io_o_dist_bus_2 = reset ? 32'h0 : w_dist_bus_2; // @[Benes.scala 85:23]
  assign io_o_dist_bus_3 = reset ? 32'h0 : w_dist_bus_3; // @[Benes.scala 85:23]
  assign io_o_dist_bus_4 = reset ? 32'h0 : w_dist_bus_4; // @[Benes.scala 85:23]
  assign io_o_dist_bus_5 = reset ? 32'h0 : w_dist_bus_5; // @[Benes.scala 85:23]
  assign io_o_dist_bus_6 = reset ? 32'h0 : w_dist_bus_6; // @[Benes.scala 85:23]
  assign io_o_dist_bus_7 = reset ? 32'h0 : w_dist_bus_7; // @[Benes.scala 85:23]
  assign io_o_dist_bus_8 = reset ? 32'h0 : w_dist_bus_8; // @[Benes.scala 85:23]
  assign io_o_dist_bus_9 = reset ? 32'h0 : w_dist_bus_9; // @[Benes.scala 85:23]
  assign io_o_dist_bus_10 = reset ? 32'h0 : w_dist_bus_10; // @[Benes.scala 85:23]
  assign io_o_dist_bus_11 = reset ? 32'h0 : w_dist_bus_11; // @[Benes.scala 85:23]
  assign io_o_dist_bus_12 = reset ? 32'h0 : w_dist_bus_12; // @[Benes.scala 85:23]
  assign io_o_dist_bus_13 = reset ? 32'h0 : w_dist_bus_13; // @[Benes.scala 85:23]
  assign io_o_dist_bus_14 = reset ? 32'h0 : w_dist_bus_14; // @[Benes.scala 85:23]
  assign io_o_dist_bus_15 = reset ? 32'h0 : w_dist_bus_15; // @[Benes.scala 85:23]
  assign io_o_dist_bus_16 = reset ? 32'h0 : w_dist_bus_16; // @[Benes.scala 85:23]
  assign io_o_dist_bus_17 = reset ? 32'h0 : w_dist_bus_17; // @[Benes.scala 85:23]
  assign io_o_dist_bus_18 = reset ? 32'h0 : w_dist_bus_18; // @[Benes.scala 85:23]
  assign io_o_dist_bus_19 = reset ? 32'h0 : w_dist_bus_19; // @[Benes.scala 85:23]
  assign io_o_dist_bus_20 = reset ? 32'h0 : w_dist_bus_20; // @[Benes.scala 85:23]
  assign io_o_dist_bus_21 = reset ? 32'h0 : w_dist_bus_21; // @[Benes.scala 85:23]
  assign io_o_dist_bus_22 = reset ? 32'h0 : w_dist_bus_22; // @[Benes.scala 85:23]
  assign io_o_dist_bus_23 = reset ? 32'h0 : w_dist_bus_23; // @[Benes.scala 85:23]
  assign io_o_dist_bus_24 = reset ? 32'h0 : w_dist_bus_24; // @[Benes.scala 85:23]
  assign io_o_dist_bus_25 = reset ? 32'h0 : w_dist_bus_25; // @[Benes.scala 85:23]
  assign io_o_dist_bus_26 = reset ? 32'h0 : w_dist_bus_26; // @[Benes.scala 85:23]
  assign io_o_dist_bus_27 = reset ? 32'h0 : w_dist_bus_27; // @[Benes.scala 85:23]
  assign io_o_dist_bus_28 = reset ? 32'h0 : w_dist_bus_28; // @[Benes.scala 85:23]
  assign io_o_dist_bus_29 = reset ? 32'h0 : w_dist_bus_29; // @[Benes.scala 85:23]
  assign io_o_dist_bus_30 = reset ? 32'h0 : w_dist_bus_30; // @[Benes.scala 85:23]
  assign io_o_dist_bus_31 = reset ? 32'h0 : w_dist_bus_31; // @[Benes.scala 85:23]
  assign in_switch_io_in = r_data_bus_ff_0; // @[Benes.scala 90:21]
  assign in_switch_1_io_in = r_data_bus_ff_1; // @[Benes.scala 90:21]
  assign in_switch_2_io_in = r_data_bus_ff_2; // @[Benes.scala 90:21]
  assign in_switch_3_io_in = r_data_bus_ff_3; // @[Benes.scala 90:21]
  assign in_switch_4_io_in = r_data_bus_ff_4; // @[Benes.scala 90:21]
  assign in_switch_5_io_in = r_data_bus_ff_5; // @[Benes.scala 90:21]
  assign in_switch_6_io_in = r_data_bus_ff_6; // @[Benes.scala 90:21]
  assign in_switch_7_io_in = r_data_bus_ff_7; // @[Benes.scala 90:21]
  assign in_switch_8_io_in = r_data_bus_ff_8; // @[Benes.scala 90:21]
  assign in_switch_9_io_in = r_data_bus_ff_9; // @[Benes.scala 90:21]
  assign in_switch_10_io_in = r_data_bus_ff_10; // @[Benes.scala 90:21]
  assign in_switch_11_io_in = r_data_bus_ff_11; // @[Benes.scala 90:21]
  assign in_switch_12_io_in = r_data_bus_ff_12; // @[Benes.scala 90:21]
  assign in_switch_13_io_in = r_data_bus_ff_13; // @[Benes.scala 90:21]
  assign in_switch_14_io_in = r_data_bus_ff_14; // @[Benes.scala 90:21]
  assign in_switch_15_io_in = r_data_bus_ff_15; // @[Benes.scala 90:21]
  assign in_switch_16_io_in = r_data_bus_ff_16; // @[Benes.scala 90:21]
  assign in_switch_17_io_in = r_data_bus_ff_17; // @[Benes.scala 90:21]
  assign in_switch_18_io_in = r_data_bus_ff_18; // @[Benes.scala 90:21]
  assign in_switch_19_io_in = r_data_bus_ff_19; // @[Benes.scala 90:21]
  assign in_switch_20_io_in = r_data_bus_ff_20; // @[Benes.scala 90:21]
  assign in_switch_21_io_in = r_data_bus_ff_21; // @[Benes.scala 90:21]
  assign in_switch_22_io_in = r_data_bus_ff_22; // @[Benes.scala 90:21]
  assign in_switch_23_io_in = r_data_bus_ff_23; // @[Benes.scala 90:21]
  assign in_switch_24_io_in = r_data_bus_ff_24; // @[Benes.scala 90:21]
  assign in_switch_25_io_in = r_data_bus_ff_25; // @[Benes.scala 90:21]
  assign in_switch_26_io_in = r_data_bus_ff_26; // @[Benes.scala 90:21]
  assign in_switch_27_io_in = r_data_bus_ff_27; // @[Benes.scala 90:21]
  assign in_switch_28_io_in = r_data_bus_ff_28; // @[Benes.scala 90:21]
  assign in_switch_29_io_in = r_data_bus_ff_29; // @[Benes.scala 90:21]
  assign in_switch_30_io_in = r_data_bus_ff_30; // @[Benes.scala 90:21]
  assign in_switch_31_io_in = r_data_bus_ff_31; // @[Benes.scala 90:21]
  assign out_switch_io_in0 = w_internal_18; // @[Benes.scala 99:23]
  assign out_switch_io_in1 = w_internal_39; // @[Benes.scala 100:23]
  assign out_switch_io_sel = r_mux_bus_ff_576; // @[Benes.scala 101:23]
  assign out_switch_1_io_in0 = w_internal_38; // @[Benes.scala 99:23]
  assign out_switch_1_io_in1 = w_internal_19; // @[Benes.scala 100:23]
  assign out_switch_1_io_sel = r_mux_bus_ff_577; // @[Benes.scala 101:23]
  assign out_switch_2_io_in0 = w_internal_58; // @[Benes.scala 99:23]
  assign out_switch_2_io_in1 = w_internal_79; // @[Benes.scala 100:23]
  assign out_switch_2_io_sel = r_mux_bus_ff_578; // @[Benes.scala 101:23]
  assign out_switch_3_io_in0 = w_internal_78; // @[Benes.scala 99:23]
  assign out_switch_3_io_in1 = w_internal_59; // @[Benes.scala 100:23]
  assign out_switch_3_io_sel = r_mux_bus_ff_579; // @[Benes.scala 101:23]
  assign out_switch_4_io_in0 = w_internal_98; // @[Benes.scala 99:23]
  assign out_switch_4_io_in1 = w_internal_119; // @[Benes.scala 100:23]
  assign out_switch_4_io_sel = r_mux_bus_ff_580; // @[Benes.scala 101:23]
  assign out_switch_5_io_in0 = w_internal_118; // @[Benes.scala 99:23]
  assign out_switch_5_io_in1 = w_internal_99; // @[Benes.scala 100:23]
  assign out_switch_5_io_sel = r_mux_bus_ff_581; // @[Benes.scala 101:23]
  assign out_switch_6_io_in0 = w_internal_138; // @[Benes.scala 99:23]
  assign out_switch_6_io_in1 = w_internal_159; // @[Benes.scala 100:23]
  assign out_switch_6_io_sel = r_mux_bus_ff_582; // @[Benes.scala 101:23]
  assign out_switch_7_io_in0 = w_internal_158; // @[Benes.scala 99:23]
  assign out_switch_7_io_in1 = w_internal_139; // @[Benes.scala 100:23]
  assign out_switch_7_io_sel = r_mux_bus_ff_583; // @[Benes.scala 101:23]
  assign out_switch_8_io_in0 = w_internal_178; // @[Benes.scala 99:23]
  assign out_switch_8_io_in1 = w_internal_199; // @[Benes.scala 100:23]
  assign out_switch_8_io_sel = r_mux_bus_ff_584; // @[Benes.scala 101:23]
  assign out_switch_9_io_in0 = w_internal_198; // @[Benes.scala 99:23]
  assign out_switch_9_io_in1 = w_internal_179; // @[Benes.scala 100:23]
  assign out_switch_9_io_sel = r_mux_bus_ff_585; // @[Benes.scala 101:23]
  assign out_switch_10_io_in0 = w_internal_218; // @[Benes.scala 99:23]
  assign out_switch_10_io_in1 = w_internal_239; // @[Benes.scala 100:23]
  assign out_switch_10_io_sel = r_mux_bus_ff_586; // @[Benes.scala 101:23]
  assign out_switch_11_io_in0 = w_internal_238; // @[Benes.scala 99:23]
  assign out_switch_11_io_in1 = w_internal_219; // @[Benes.scala 100:23]
  assign out_switch_11_io_sel = r_mux_bus_ff_587; // @[Benes.scala 101:23]
  assign out_switch_12_io_in0 = w_internal_258; // @[Benes.scala 99:23]
  assign out_switch_12_io_in1 = w_internal_279; // @[Benes.scala 100:23]
  assign out_switch_12_io_sel = r_mux_bus_ff_588; // @[Benes.scala 101:23]
  assign out_switch_13_io_in0 = w_internal_278; // @[Benes.scala 99:23]
  assign out_switch_13_io_in1 = w_internal_259; // @[Benes.scala 100:23]
  assign out_switch_13_io_sel = r_mux_bus_ff_589; // @[Benes.scala 101:23]
  assign out_switch_14_io_in0 = w_internal_298; // @[Benes.scala 99:23]
  assign out_switch_14_io_in1 = w_internal_319; // @[Benes.scala 100:23]
  assign out_switch_14_io_sel = r_mux_bus_ff_590; // @[Benes.scala 101:23]
  assign out_switch_15_io_in0 = w_internal_318; // @[Benes.scala 99:23]
  assign out_switch_15_io_in1 = w_internal_299; // @[Benes.scala 100:23]
  assign out_switch_15_io_sel = r_mux_bus_ff_591; // @[Benes.scala 101:23]
  assign out_switch_16_io_in0 = w_internal_338; // @[Benes.scala 99:23]
  assign out_switch_16_io_in1 = w_internal_359; // @[Benes.scala 100:23]
  assign out_switch_16_io_sel = r_mux_bus_ff_592; // @[Benes.scala 101:23]
  assign out_switch_17_io_in0 = w_internal_358; // @[Benes.scala 99:23]
  assign out_switch_17_io_in1 = w_internal_339; // @[Benes.scala 100:23]
  assign out_switch_17_io_sel = r_mux_bus_ff_593; // @[Benes.scala 101:23]
  assign out_switch_18_io_in0 = w_internal_378; // @[Benes.scala 99:23]
  assign out_switch_18_io_in1 = w_internal_399; // @[Benes.scala 100:23]
  assign out_switch_18_io_sel = r_mux_bus_ff_594; // @[Benes.scala 101:23]
  assign out_switch_19_io_in0 = w_internal_398; // @[Benes.scala 99:23]
  assign out_switch_19_io_in1 = w_internal_379; // @[Benes.scala 100:23]
  assign out_switch_19_io_sel = r_mux_bus_ff_595; // @[Benes.scala 101:23]
  assign out_switch_20_io_in0 = w_internal_418; // @[Benes.scala 99:23]
  assign out_switch_20_io_in1 = w_internal_439; // @[Benes.scala 100:23]
  assign out_switch_20_io_sel = r_mux_bus_ff_596; // @[Benes.scala 101:23]
  assign out_switch_21_io_in0 = w_internal_438; // @[Benes.scala 99:23]
  assign out_switch_21_io_in1 = w_internal_419; // @[Benes.scala 100:23]
  assign out_switch_21_io_sel = r_mux_bus_ff_597; // @[Benes.scala 101:23]
  assign out_switch_22_io_in0 = w_internal_458; // @[Benes.scala 99:23]
  assign out_switch_22_io_in1 = w_internal_479; // @[Benes.scala 100:23]
  assign out_switch_22_io_sel = r_mux_bus_ff_598; // @[Benes.scala 101:23]
  assign out_switch_23_io_in0 = w_internal_478; // @[Benes.scala 99:23]
  assign out_switch_23_io_in1 = w_internal_459; // @[Benes.scala 100:23]
  assign out_switch_23_io_sel = r_mux_bus_ff_599; // @[Benes.scala 101:23]
  assign out_switch_24_io_in0 = w_internal_498; // @[Benes.scala 99:23]
  assign out_switch_24_io_in1 = w_internal_519; // @[Benes.scala 100:23]
  assign out_switch_24_io_sel = r_mux_bus_ff_600; // @[Benes.scala 101:23]
  assign out_switch_25_io_in0 = w_internal_518; // @[Benes.scala 99:23]
  assign out_switch_25_io_in1 = w_internal_499; // @[Benes.scala 100:23]
  assign out_switch_25_io_sel = r_mux_bus_ff_601; // @[Benes.scala 101:23]
  assign out_switch_26_io_in0 = w_internal_538; // @[Benes.scala 99:23]
  assign out_switch_26_io_in1 = w_internal_559; // @[Benes.scala 100:23]
  assign out_switch_26_io_sel = r_mux_bus_ff_602; // @[Benes.scala 101:23]
  assign out_switch_27_io_in0 = w_internal_558; // @[Benes.scala 99:23]
  assign out_switch_27_io_in1 = w_internal_539; // @[Benes.scala 100:23]
  assign out_switch_27_io_sel = r_mux_bus_ff_603; // @[Benes.scala 101:23]
  assign out_switch_28_io_in0 = w_internal_578; // @[Benes.scala 99:23]
  assign out_switch_28_io_in1 = w_internal_599; // @[Benes.scala 100:23]
  assign out_switch_28_io_sel = r_mux_bus_ff_604; // @[Benes.scala 101:23]
  assign out_switch_29_io_in0 = w_internal_598; // @[Benes.scala 99:23]
  assign out_switch_29_io_in1 = w_internal_579; // @[Benes.scala 100:23]
  assign out_switch_29_io_sel = r_mux_bus_ff_605; // @[Benes.scala 101:23]
  assign out_switch_30_io_in0 = w_internal_618; // @[Benes.scala 99:23]
  assign out_switch_30_io_in1 = w_internal_639; // @[Benes.scala 100:23]
  assign out_switch_30_io_sel = r_mux_bus_ff_606; // @[Benes.scala 101:23]
  assign out_switch_31_io_in0 = w_internal_638; // @[Benes.scala 99:23]
  assign out_switch_31_io_in1 = w_internal_619; // @[Benes.scala 100:23]
  assign out_switch_31_io_sel = r_mux_bus_ff_607; // @[Benes.scala 101:23]
  assign imm_switch_io_in0 = w_internal_0; // @[Benes.scala 109:25]
  assign imm_switch_io_in1 = w_internal_21; // @[Benes.scala 112:29]
  assign imm_switch_io_sel0 = r_mux_bus_ff_0; // @[Benes.scala 123:26]
  assign imm_switch_io_sel1 = r_mux_bus_ff_1; // @[Benes.scala 124:26]
  assign imm_switch_1_io_in0 = w_internal_2; // @[Benes.scala 109:25]
  assign imm_switch_1_io_in1 = w_internal_43; // @[Benes.scala 112:29]
  assign imm_switch_1_io_sel0 = r_mux_bus_ff_2; // @[Benes.scala 123:26]
  assign imm_switch_1_io_sel1 = r_mux_bus_ff_3; // @[Benes.scala 124:26]
  assign imm_switch_2_io_in0 = w_internal_4; // @[Benes.scala 109:25]
  assign imm_switch_2_io_in1 = w_internal_85; // @[Benes.scala 112:29]
  assign imm_switch_2_io_sel0 = r_mux_bus_ff_4; // @[Benes.scala 123:26]
  assign imm_switch_2_io_sel1 = r_mux_bus_ff_5; // @[Benes.scala 124:26]
  assign imm_switch_3_io_in0 = w_internal_6; // @[Benes.scala 109:25]
  assign imm_switch_3_io_in1 = w_internal_167; // @[Benes.scala 112:29]
  assign imm_switch_3_io_sel0 = r_mux_bus_ff_6; // @[Benes.scala 123:26]
  assign imm_switch_3_io_sel1 = r_mux_bus_ff_7; // @[Benes.scala 124:26]
  assign imm_switch_4_io_in0 = w_internal_8; // @[Benes.scala 109:25]
  assign imm_switch_4_io_in1 = w_internal_329; // @[Benes.scala 112:29]
  assign imm_switch_4_io_sel0 = r_mux_bus_ff_8; // @[Benes.scala 123:26]
  assign imm_switch_4_io_sel1 = r_mux_bus_ff_9; // @[Benes.scala 124:26]
  assign imm_switch_5_io_in0 = w_internal_10; // @[Benes.scala 109:25]
  assign imm_switch_5_io_in1 = w_internal_331; // @[Benes.scala 118:29]
  assign imm_switch_5_io_sel0 = r_mux_bus_ff_10; // @[Benes.scala 123:26]
  assign imm_switch_5_io_sel1 = r_mux_bus_ff_11; // @[Benes.scala 124:26]
  assign imm_switch_6_io_in0 = w_internal_12; // @[Benes.scala 109:25]
  assign imm_switch_6_io_in1 = w_internal_173; // @[Benes.scala 118:29]
  assign imm_switch_6_io_sel0 = r_mux_bus_ff_12; // @[Benes.scala 123:26]
  assign imm_switch_6_io_sel1 = r_mux_bus_ff_13; // @[Benes.scala 124:26]
  assign imm_switch_7_io_in0 = w_internal_14; // @[Benes.scala 109:25]
  assign imm_switch_7_io_in1 = w_internal_95; // @[Benes.scala 118:29]
  assign imm_switch_7_io_sel0 = r_mux_bus_ff_14; // @[Benes.scala 123:26]
  assign imm_switch_7_io_sel1 = r_mux_bus_ff_15; // @[Benes.scala 124:26]
  assign imm_switch_8_io_in0 = w_internal_16; // @[Benes.scala 109:25]
  assign imm_switch_8_io_in1 = w_internal_57; // @[Benes.scala 118:29]
  assign imm_switch_8_io_sel0 = r_mux_bus_ff_16; // @[Benes.scala 123:26]
  assign imm_switch_8_io_sel1 = r_mux_bus_ff_17; // @[Benes.scala 124:26]
  assign imm_switch_9_io_in0 = w_internal_20; // @[Benes.scala 109:25]
  assign imm_switch_9_io_in1 = w_internal_1; // @[Benes.scala 114:29]
  assign imm_switch_9_io_sel0 = r_mux_bus_ff_18; // @[Benes.scala 123:26]
  assign imm_switch_9_io_sel1 = r_mux_bus_ff_19; // @[Benes.scala 124:26]
  assign imm_switch_10_io_in0 = w_internal_22; // @[Benes.scala 109:25]
  assign imm_switch_10_io_in1 = w_internal_63; // @[Benes.scala 112:29]
  assign imm_switch_10_io_sel0 = r_mux_bus_ff_20; // @[Benes.scala 123:26]
  assign imm_switch_10_io_sel1 = r_mux_bus_ff_21; // @[Benes.scala 124:26]
  assign imm_switch_11_io_in0 = w_internal_24; // @[Benes.scala 109:25]
  assign imm_switch_11_io_in1 = w_internal_105; // @[Benes.scala 112:29]
  assign imm_switch_11_io_sel0 = r_mux_bus_ff_22; // @[Benes.scala 123:26]
  assign imm_switch_11_io_sel1 = r_mux_bus_ff_23; // @[Benes.scala 124:26]
  assign imm_switch_12_io_in0 = w_internal_26; // @[Benes.scala 109:25]
  assign imm_switch_12_io_in1 = w_internal_187; // @[Benes.scala 112:29]
  assign imm_switch_12_io_sel0 = r_mux_bus_ff_24; // @[Benes.scala 123:26]
  assign imm_switch_12_io_sel1 = r_mux_bus_ff_25; // @[Benes.scala 124:26]
  assign imm_switch_13_io_in0 = w_internal_28; // @[Benes.scala 109:25]
  assign imm_switch_13_io_in1 = w_internal_349; // @[Benes.scala 112:29]
  assign imm_switch_13_io_sel0 = r_mux_bus_ff_26; // @[Benes.scala 123:26]
  assign imm_switch_13_io_sel1 = r_mux_bus_ff_27; // @[Benes.scala 124:26]
  assign imm_switch_14_io_in0 = w_internal_30; // @[Benes.scala 109:25]
  assign imm_switch_14_io_in1 = w_internal_351; // @[Benes.scala 118:29]
  assign imm_switch_14_io_sel0 = r_mux_bus_ff_28; // @[Benes.scala 123:26]
  assign imm_switch_14_io_sel1 = r_mux_bus_ff_29; // @[Benes.scala 124:26]
  assign imm_switch_15_io_in0 = w_internal_32; // @[Benes.scala 109:25]
  assign imm_switch_15_io_in1 = w_internal_193; // @[Benes.scala 118:29]
  assign imm_switch_15_io_sel0 = r_mux_bus_ff_30; // @[Benes.scala 123:26]
  assign imm_switch_15_io_sel1 = r_mux_bus_ff_31; // @[Benes.scala 124:26]
  assign imm_switch_16_io_in0 = w_internal_34; // @[Benes.scala 109:25]
  assign imm_switch_16_io_in1 = w_internal_115; // @[Benes.scala 118:29]
  assign imm_switch_16_io_sel0 = r_mux_bus_ff_32; // @[Benes.scala 123:26]
  assign imm_switch_16_io_sel1 = r_mux_bus_ff_33; // @[Benes.scala 124:26]
  assign imm_switch_17_io_in0 = w_internal_36; // @[Benes.scala 109:25]
  assign imm_switch_17_io_in1 = w_internal_77; // @[Benes.scala 118:29]
  assign imm_switch_17_io_sel0 = r_mux_bus_ff_34; // @[Benes.scala 123:26]
  assign imm_switch_17_io_sel1 = r_mux_bus_ff_35; // @[Benes.scala 124:26]
  assign imm_switch_18_io_in0 = w_internal_40; // @[Benes.scala 109:25]
  assign imm_switch_18_io_in1 = w_internal_61; // @[Benes.scala 112:29]
  assign imm_switch_18_io_sel0 = r_mux_bus_ff_36; // @[Benes.scala 123:26]
  assign imm_switch_18_io_sel1 = r_mux_bus_ff_37; // @[Benes.scala 124:26]
  assign imm_switch_19_io_in0 = w_internal_42; // @[Benes.scala 109:25]
  assign imm_switch_19_io_in1 = w_internal_3; // @[Benes.scala 114:29]
  assign imm_switch_19_io_sel0 = r_mux_bus_ff_38; // @[Benes.scala 123:26]
  assign imm_switch_19_io_sel1 = r_mux_bus_ff_39; // @[Benes.scala 124:26]
  assign imm_switch_20_io_in0 = w_internal_44; // @[Benes.scala 109:25]
  assign imm_switch_20_io_in1 = w_internal_125; // @[Benes.scala 112:29]
  assign imm_switch_20_io_sel0 = r_mux_bus_ff_40; // @[Benes.scala 123:26]
  assign imm_switch_20_io_sel1 = r_mux_bus_ff_41; // @[Benes.scala 124:26]
  assign imm_switch_21_io_in0 = w_internal_46; // @[Benes.scala 109:25]
  assign imm_switch_21_io_in1 = w_internal_207; // @[Benes.scala 112:29]
  assign imm_switch_21_io_sel0 = r_mux_bus_ff_42; // @[Benes.scala 123:26]
  assign imm_switch_21_io_sel1 = r_mux_bus_ff_43; // @[Benes.scala 124:26]
  assign imm_switch_22_io_in0 = w_internal_48; // @[Benes.scala 109:25]
  assign imm_switch_22_io_in1 = w_internal_369; // @[Benes.scala 112:29]
  assign imm_switch_22_io_sel0 = r_mux_bus_ff_44; // @[Benes.scala 123:26]
  assign imm_switch_22_io_sel1 = r_mux_bus_ff_45; // @[Benes.scala 124:26]
  assign imm_switch_23_io_in0 = w_internal_50; // @[Benes.scala 109:25]
  assign imm_switch_23_io_in1 = w_internal_371; // @[Benes.scala 118:29]
  assign imm_switch_23_io_sel0 = r_mux_bus_ff_46; // @[Benes.scala 123:26]
  assign imm_switch_23_io_sel1 = r_mux_bus_ff_47; // @[Benes.scala 124:26]
  assign imm_switch_24_io_in0 = w_internal_52; // @[Benes.scala 109:25]
  assign imm_switch_24_io_in1 = w_internal_213; // @[Benes.scala 118:29]
  assign imm_switch_24_io_sel0 = r_mux_bus_ff_48; // @[Benes.scala 123:26]
  assign imm_switch_24_io_sel1 = r_mux_bus_ff_49; // @[Benes.scala 124:26]
  assign imm_switch_25_io_in0 = w_internal_54; // @[Benes.scala 109:25]
  assign imm_switch_25_io_in1 = w_internal_135; // @[Benes.scala 118:29]
  assign imm_switch_25_io_sel0 = r_mux_bus_ff_50; // @[Benes.scala 123:26]
  assign imm_switch_25_io_sel1 = r_mux_bus_ff_51; // @[Benes.scala 124:26]
  assign imm_switch_26_io_in0 = w_internal_56; // @[Benes.scala 109:25]
  assign imm_switch_26_io_in1 = w_internal_17; // @[Benes.scala 120:29]
  assign imm_switch_26_io_sel0 = r_mux_bus_ff_52; // @[Benes.scala 123:26]
  assign imm_switch_26_io_sel1 = r_mux_bus_ff_53; // @[Benes.scala 124:26]
  assign imm_switch_27_io_in0 = w_internal_60; // @[Benes.scala 109:25]
  assign imm_switch_27_io_in1 = w_internal_41; // @[Benes.scala 114:29]
  assign imm_switch_27_io_sel0 = r_mux_bus_ff_54; // @[Benes.scala 123:26]
  assign imm_switch_27_io_sel1 = r_mux_bus_ff_55; // @[Benes.scala 124:26]
  assign imm_switch_28_io_in0 = w_internal_62; // @[Benes.scala 109:25]
  assign imm_switch_28_io_in1 = w_internal_23; // @[Benes.scala 114:29]
  assign imm_switch_28_io_sel0 = r_mux_bus_ff_56; // @[Benes.scala 123:26]
  assign imm_switch_28_io_sel1 = r_mux_bus_ff_57; // @[Benes.scala 124:26]
  assign imm_switch_29_io_in0 = w_internal_64; // @[Benes.scala 109:25]
  assign imm_switch_29_io_in1 = w_internal_145; // @[Benes.scala 112:29]
  assign imm_switch_29_io_sel0 = r_mux_bus_ff_58; // @[Benes.scala 123:26]
  assign imm_switch_29_io_sel1 = r_mux_bus_ff_59; // @[Benes.scala 124:26]
  assign imm_switch_30_io_in0 = w_internal_66; // @[Benes.scala 109:25]
  assign imm_switch_30_io_in1 = w_internal_227; // @[Benes.scala 112:29]
  assign imm_switch_30_io_sel0 = r_mux_bus_ff_60; // @[Benes.scala 123:26]
  assign imm_switch_30_io_sel1 = r_mux_bus_ff_61; // @[Benes.scala 124:26]
  assign imm_switch_31_io_in0 = w_internal_68; // @[Benes.scala 109:25]
  assign imm_switch_31_io_in1 = w_internal_389; // @[Benes.scala 112:29]
  assign imm_switch_31_io_sel0 = r_mux_bus_ff_62; // @[Benes.scala 123:26]
  assign imm_switch_31_io_sel1 = r_mux_bus_ff_63; // @[Benes.scala 124:26]
  assign imm_switch_32_io_in0 = w_internal_70; // @[Benes.scala 109:25]
  assign imm_switch_32_io_in1 = w_internal_391; // @[Benes.scala 118:29]
  assign imm_switch_32_io_sel0 = r_mux_bus_ff_64; // @[Benes.scala 123:26]
  assign imm_switch_32_io_sel1 = r_mux_bus_ff_65; // @[Benes.scala 124:26]
  assign imm_switch_33_io_in0 = w_internal_72; // @[Benes.scala 109:25]
  assign imm_switch_33_io_in1 = w_internal_233; // @[Benes.scala 118:29]
  assign imm_switch_33_io_sel0 = r_mux_bus_ff_66; // @[Benes.scala 123:26]
  assign imm_switch_33_io_sel1 = r_mux_bus_ff_67; // @[Benes.scala 124:26]
  assign imm_switch_34_io_in0 = w_internal_74; // @[Benes.scala 109:25]
  assign imm_switch_34_io_in1 = w_internal_155; // @[Benes.scala 118:29]
  assign imm_switch_34_io_sel0 = r_mux_bus_ff_68; // @[Benes.scala 123:26]
  assign imm_switch_34_io_sel1 = r_mux_bus_ff_69; // @[Benes.scala 124:26]
  assign imm_switch_35_io_in0 = w_internal_76; // @[Benes.scala 109:25]
  assign imm_switch_35_io_in1 = w_internal_37; // @[Benes.scala 120:29]
  assign imm_switch_35_io_sel0 = r_mux_bus_ff_70; // @[Benes.scala 123:26]
  assign imm_switch_35_io_sel1 = r_mux_bus_ff_71; // @[Benes.scala 124:26]
  assign imm_switch_36_io_in0 = w_internal_80; // @[Benes.scala 109:25]
  assign imm_switch_36_io_in1 = w_internal_101; // @[Benes.scala 112:29]
  assign imm_switch_36_io_sel0 = r_mux_bus_ff_72; // @[Benes.scala 123:26]
  assign imm_switch_36_io_sel1 = r_mux_bus_ff_73; // @[Benes.scala 124:26]
  assign imm_switch_37_io_in0 = w_internal_82; // @[Benes.scala 109:25]
  assign imm_switch_37_io_in1 = w_internal_123; // @[Benes.scala 112:29]
  assign imm_switch_37_io_sel0 = r_mux_bus_ff_74; // @[Benes.scala 123:26]
  assign imm_switch_37_io_sel1 = r_mux_bus_ff_75; // @[Benes.scala 124:26]
  assign imm_switch_38_io_in0 = w_internal_84; // @[Benes.scala 109:25]
  assign imm_switch_38_io_in1 = w_internal_5; // @[Benes.scala 114:29]
  assign imm_switch_38_io_sel0 = r_mux_bus_ff_76; // @[Benes.scala 123:26]
  assign imm_switch_38_io_sel1 = r_mux_bus_ff_77; // @[Benes.scala 124:26]
  assign imm_switch_39_io_in0 = w_internal_86; // @[Benes.scala 109:25]
  assign imm_switch_39_io_in1 = w_internal_247; // @[Benes.scala 112:29]
  assign imm_switch_39_io_sel0 = r_mux_bus_ff_78; // @[Benes.scala 123:26]
  assign imm_switch_39_io_sel1 = r_mux_bus_ff_79; // @[Benes.scala 124:26]
  assign imm_switch_40_io_in0 = w_internal_88; // @[Benes.scala 109:25]
  assign imm_switch_40_io_in1 = w_internal_409; // @[Benes.scala 112:29]
  assign imm_switch_40_io_sel0 = r_mux_bus_ff_80; // @[Benes.scala 123:26]
  assign imm_switch_40_io_sel1 = r_mux_bus_ff_81; // @[Benes.scala 124:26]
  assign imm_switch_41_io_in0 = w_internal_90; // @[Benes.scala 109:25]
  assign imm_switch_41_io_in1 = w_internal_411; // @[Benes.scala 118:29]
  assign imm_switch_41_io_sel0 = r_mux_bus_ff_82; // @[Benes.scala 123:26]
  assign imm_switch_41_io_sel1 = r_mux_bus_ff_83; // @[Benes.scala 124:26]
  assign imm_switch_42_io_in0 = w_internal_92; // @[Benes.scala 109:25]
  assign imm_switch_42_io_in1 = w_internal_253; // @[Benes.scala 118:29]
  assign imm_switch_42_io_sel0 = r_mux_bus_ff_84; // @[Benes.scala 123:26]
  assign imm_switch_42_io_sel1 = r_mux_bus_ff_85; // @[Benes.scala 124:26]
  assign imm_switch_43_io_in0 = w_internal_94; // @[Benes.scala 109:25]
  assign imm_switch_43_io_in1 = w_internal_15; // @[Benes.scala 120:29]
  assign imm_switch_43_io_sel0 = r_mux_bus_ff_86; // @[Benes.scala 123:26]
  assign imm_switch_43_io_sel1 = r_mux_bus_ff_87; // @[Benes.scala 124:26]
  assign imm_switch_44_io_in0 = w_internal_96; // @[Benes.scala 109:25]
  assign imm_switch_44_io_in1 = w_internal_137; // @[Benes.scala 118:29]
  assign imm_switch_44_io_sel0 = r_mux_bus_ff_88; // @[Benes.scala 123:26]
  assign imm_switch_44_io_sel1 = r_mux_bus_ff_89; // @[Benes.scala 124:26]
  assign imm_switch_45_io_in0 = w_internal_100; // @[Benes.scala 109:25]
  assign imm_switch_45_io_in1 = w_internal_81; // @[Benes.scala 114:29]
  assign imm_switch_45_io_sel0 = r_mux_bus_ff_90; // @[Benes.scala 123:26]
  assign imm_switch_45_io_sel1 = r_mux_bus_ff_91; // @[Benes.scala 124:26]
  assign imm_switch_46_io_in0 = w_internal_102; // @[Benes.scala 109:25]
  assign imm_switch_46_io_in1 = w_internal_143; // @[Benes.scala 112:29]
  assign imm_switch_46_io_sel0 = r_mux_bus_ff_92; // @[Benes.scala 123:26]
  assign imm_switch_46_io_sel1 = r_mux_bus_ff_93; // @[Benes.scala 124:26]
  assign imm_switch_47_io_in0 = w_internal_104; // @[Benes.scala 109:25]
  assign imm_switch_47_io_in1 = w_internal_25; // @[Benes.scala 114:29]
  assign imm_switch_47_io_sel0 = r_mux_bus_ff_94; // @[Benes.scala 123:26]
  assign imm_switch_47_io_sel1 = r_mux_bus_ff_95; // @[Benes.scala 124:26]
  assign imm_switch_48_io_in0 = w_internal_106; // @[Benes.scala 109:25]
  assign imm_switch_48_io_in1 = w_internal_267; // @[Benes.scala 112:29]
  assign imm_switch_48_io_sel0 = r_mux_bus_ff_96; // @[Benes.scala 123:26]
  assign imm_switch_48_io_sel1 = r_mux_bus_ff_97; // @[Benes.scala 124:26]
  assign imm_switch_49_io_in0 = w_internal_108; // @[Benes.scala 109:25]
  assign imm_switch_49_io_in1 = w_internal_429; // @[Benes.scala 112:29]
  assign imm_switch_49_io_sel0 = r_mux_bus_ff_98; // @[Benes.scala 123:26]
  assign imm_switch_49_io_sel1 = r_mux_bus_ff_99; // @[Benes.scala 124:26]
  assign imm_switch_50_io_in0 = w_internal_110; // @[Benes.scala 109:25]
  assign imm_switch_50_io_in1 = w_internal_431; // @[Benes.scala 118:29]
  assign imm_switch_50_io_sel0 = r_mux_bus_ff_100; // @[Benes.scala 123:26]
  assign imm_switch_50_io_sel1 = r_mux_bus_ff_101; // @[Benes.scala 124:26]
  assign imm_switch_51_io_in0 = w_internal_112; // @[Benes.scala 109:25]
  assign imm_switch_51_io_in1 = w_internal_273; // @[Benes.scala 118:29]
  assign imm_switch_51_io_sel0 = r_mux_bus_ff_102; // @[Benes.scala 123:26]
  assign imm_switch_51_io_sel1 = r_mux_bus_ff_103; // @[Benes.scala 124:26]
  assign imm_switch_52_io_in0 = w_internal_114; // @[Benes.scala 109:25]
  assign imm_switch_52_io_in1 = w_internal_35; // @[Benes.scala 120:29]
  assign imm_switch_52_io_sel0 = r_mux_bus_ff_104; // @[Benes.scala 123:26]
  assign imm_switch_52_io_sel1 = r_mux_bus_ff_105; // @[Benes.scala 124:26]
  assign imm_switch_53_io_in0 = w_internal_116; // @[Benes.scala 109:25]
  assign imm_switch_53_io_in1 = w_internal_157; // @[Benes.scala 118:29]
  assign imm_switch_53_io_sel0 = r_mux_bus_ff_106; // @[Benes.scala 123:26]
  assign imm_switch_53_io_sel1 = r_mux_bus_ff_107; // @[Benes.scala 124:26]
  assign imm_switch_54_io_in0 = w_internal_120; // @[Benes.scala 109:25]
  assign imm_switch_54_io_in1 = w_internal_141; // @[Benes.scala 112:29]
  assign imm_switch_54_io_sel0 = r_mux_bus_ff_108; // @[Benes.scala 123:26]
  assign imm_switch_54_io_sel1 = r_mux_bus_ff_109; // @[Benes.scala 124:26]
  assign imm_switch_55_io_in0 = w_internal_122; // @[Benes.scala 109:25]
  assign imm_switch_55_io_in1 = w_internal_83; // @[Benes.scala 114:29]
  assign imm_switch_55_io_sel0 = r_mux_bus_ff_110; // @[Benes.scala 123:26]
  assign imm_switch_55_io_sel1 = r_mux_bus_ff_111; // @[Benes.scala 124:26]
  assign imm_switch_56_io_in0 = w_internal_124; // @[Benes.scala 109:25]
  assign imm_switch_56_io_in1 = w_internal_45; // @[Benes.scala 114:29]
  assign imm_switch_56_io_sel0 = r_mux_bus_ff_112; // @[Benes.scala 123:26]
  assign imm_switch_56_io_sel1 = r_mux_bus_ff_113; // @[Benes.scala 124:26]
  assign imm_switch_57_io_in0 = w_internal_126; // @[Benes.scala 109:25]
  assign imm_switch_57_io_in1 = w_internal_287; // @[Benes.scala 112:29]
  assign imm_switch_57_io_sel0 = r_mux_bus_ff_114; // @[Benes.scala 123:26]
  assign imm_switch_57_io_sel1 = r_mux_bus_ff_115; // @[Benes.scala 124:26]
  assign imm_switch_58_io_in0 = w_internal_128; // @[Benes.scala 109:25]
  assign imm_switch_58_io_in1 = w_internal_449; // @[Benes.scala 112:29]
  assign imm_switch_58_io_sel0 = r_mux_bus_ff_116; // @[Benes.scala 123:26]
  assign imm_switch_58_io_sel1 = r_mux_bus_ff_117; // @[Benes.scala 124:26]
  assign imm_switch_59_io_in0 = w_internal_130; // @[Benes.scala 109:25]
  assign imm_switch_59_io_in1 = w_internal_451; // @[Benes.scala 118:29]
  assign imm_switch_59_io_sel0 = r_mux_bus_ff_118; // @[Benes.scala 123:26]
  assign imm_switch_59_io_sel1 = r_mux_bus_ff_119; // @[Benes.scala 124:26]
  assign imm_switch_60_io_in0 = w_internal_132; // @[Benes.scala 109:25]
  assign imm_switch_60_io_in1 = w_internal_293; // @[Benes.scala 118:29]
  assign imm_switch_60_io_sel0 = r_mux_bus_ff_120; // @[Benes.scala 123:26]
  assign imm_switch_60_io_sel1 = r_mux_bus_ff_121; // @[Benes.scala 124:26]
  assign imm_switch_61_io_in0 = w_internal_134; // @[Benes.scala 109:25]
  assign imm_switch_61_io_in1 = w_internal_55; // @[Benes.scala 120:29]
  assign imm_switch_61_io_sel0 = r_mux_bus_ff_122; // @[Benes.scala 123:26]
  assign imm_switch_61_io_sel1 = r_mux_bus_ff_123; // @[Benes.scala 124:26]
  assign imm_switch_62_io_in0 = w_internal_136; // @[Benes.scala 109:25]
  assign imm_switch_62_io_in1 = w_internal_97; // @[Benes.scala 120:29]
  assign imm_switch_62_io_sel0 = r_mux_bus_ff_124; // @[Benes.scala 123:26]
  assign imm_switch_62_io_sel1 = r_mux_bus_ff_125; // @[Benes.scala 124:26]
  assign imm_switch_63_io_in0 = w_internal_140; // @[Benes.scala 109:25]
  assign imm_switch_63_io_in1 = w_internal_121; // @[Benes.scala 114:29]
  assign imm_switch_63_io_sel0 = r_mux_bus_ff_126; // @[Benes.scala 123:26]
  assign imm_switch_63_io_sel1 = r_mux_bus_ff_127; // @[Benes.scala 124:26]
  assign imm_switch_64_io_in0 = w_internal_142; // @[Benes.scala 109:25]
  assign imm_switch_64_io_in1 = w_internal_103; // @[Benes.scala 114:29]
  assign imm_switch_64_io_sel0 = r_mux_bus_ff_128; // @[Benes.scala 123:26]
  assign imm_switch_64_io_sel1 = r_mux_bus_ff_129; // @[Benes.scala 124:26]
  assign imm_switch_65_io_in0 = w_internal_144; // @[Benes.scala 109:25]
  assign imm_switch_65_io_in1 = w_internal_65; // @[Benes.scala 114:29]
  assign imm_switch_65_io_sel0 = r_mux_bus_ff_130; // @[Benes.scala 123:26]
  assign imm_switch_65_io_sel1 = r_mux_bus_ff_131; // @[Benes.scala 124:26]
  assign imm_switch_66_io_in0 = w_internal_146; // @[Benes.scala 109:25]
  assign imm_switch_66_io_in1 = w_internal_307; // @[Benes.scala 112:29]
  assign imm_switch_66_io_sel0 = r_mux_bus_ff_132; // @[Benes.scala 123:26]
  assign imm_switch_66_io_sel1 = r_mux_bus_ff_133; // @[Benes.scala 124:26]
  assign imm_switch_67_io_in0 = w_internal_148; // @[Benes.scala 109:25]
  assign imm_switch_67_io_in1 = w_internal_469; // @[Benes.scala 112:29]
  assign imm_switch_67_io_sel0 = r_mux_bus_ff_134; // @[Benes.scala 123:26]
  assign imm_switch_67_io_sel1 = r_mux_bus_ff_135; // @[Benes.scala 124:26]
  assign imm_switch_68_io_in0 = w_internal_150; // @[Benes.scala 109:25]
  assign imm_switch_68_io_in1 = w_internal_471; // @[Benes.scala 118:29]
  assign imm_switch_68_io_sel0 = r_mux_bus_ff_136; // @[Benes.scala 123:26]
  assign imm_switch_68_io_sel1 = r_mux_bus_ff_137; // @[Benes.scala 124:26]
  assign imm_switch_69_io_in0 = w_internal_152; // @[Benes.scala 109:25]
  assign imm_switch_69_io_in1 = w_internal_313; // @[Benes.scala 118:29]
  assign imm_switch_69_io_sel0 = r_mux_bus_ff_138; // @[Benes.scala 123:26]
  assign imm_switch_69_io_sel1 = r_mux_bus_ff_139; // @[Benes.scala 124:26]
  assign imm_switch_70_io_in0 = w_internal_154; // @[Benes.scala 109:25]
  assign imm_switch_70_io_in1 = w_internal_75; // @[Benes.scala 120:29]
  assign imm_switch_70_io_sel0 = r_mux_bus_ff_140; // @[Benes.scala 123:26]
  assign imm_switch_70_io_sel1 = r_mux_bus_ff_141; // @[Benes.scala 124:26]
  assign imm_switch_71_io_in0 = w_internal_156; // @[Benes.scala 109:25]
  assign imm_switch_71_io_in1 = w_internal_117; // @[Benes.scala 120:29]
  assign imm_switch_71_io_sel0 = r_mux_bus_ff_142; // @[Benes.scala 123:26]
  assign imm_switch_71_io_sel1 = r_mux_bus_ff_143; // @[Benes.scala 124:26]
  assign imm_switch_72_io_in0 = w_internal_160; // @[Benes.scala 109:25]
  assign imm_switch_72_io_in1 = w_internal_181; // @[Benes.scala 112:29]
  assign imm_switch_72_io_sel0 = r_mux_bus_ff_144; // @[Benes.scala 123:26]
  assign imm_switch_72_io_sel1 = r_mux_bus_ff_145; // @[Benes.scala 124:26]
  assign imm_switch_73_io_in0 = w_internal_162; // @[Benes.scala 109:25]
  assign imm_switch_73_io_in1 = w_internal_203; // @[Benes.scala 112:29]
  assign imm_switch_73_io_sel0 = r_mux_bus_ff_146; // @[Benes.scala 123:26]
  assign imm_switch_73_io_sel1 = r_mux_bus_ff_147; // @[Benes.scala 124:26]
  assign imm_switch_74_io_in0 = w_internal_164; // @[Benes.scala 109:25]
  assign imm_switch_74_io_in1 = w_internal_245; // @[Benes.scala 112:29]
  assign imm_switch_74_io_sel0 = r_mux_bus_ff_148; // @[Benes.scala 123:26]
  assign imm_switch_74_io_sel1 = r_mux_bus_ff_149; // @[Benes.scala 124:26]
  assign imm_switch_75_io_in0 = w_internal_166; // @[Benes.scala 109:25]
  assign imm_switch_75_io_in1 = w_internal_7; // @[Benes.scala 114:29]
  assign imm_switch_75_io_sel0 = r_mux_bus_ff_150; // @[Benes.scala 123:26]
  assign imm_switch_75_io_sel1 = r_mux_bus_ff_151; // @[Benes.scala 124:26]
  assign imm_switch_76_io_in0 = w_internal_168; // @[Benes.scala 109:25]
  assign imm_switch_76_io_in1 = w_internal_489; // @[Benes.scala 112:29]
  assign imm_switch_76_io_sel0 = r_mux_bus_ff_152; // @[Benes.scala 123:26]
  assign imm_switch_76_io_sel1 = r_mux_bus_ff_153; // @[Benes.scala 124:26]
  assign imm_switch_77_io_in0 = w_internal_170; // @[Benes.scala 109:25]
  assign imm_switch_77_io_in1 = w_internal_491; // @[Benes.scala 118:29]
  assign imm_switch_77_io_sel0 = r_mux_bus_ff_154; // @[Benes.scala 123:26]
  assign imm_switch_77_io_sel1 = r_mux_bus_ff_155; // @[Benes.scala 124:26]
  assign imm_switch_78_io_in0 = w_internal_172; // @[Benes.scala 109:25]
  assign imm_switch_78_io_in1 = w_internal_13; // @[Benes.scala 120:29]
  assign imm_switch_78_io_sel0 = r_mux_bus_ff_156; // @[Benes.scala 123:26]
  assign imm_switch_78_io_sel1 = r_mux_bus_ff_157; // @[Benes.scala 124:26]
  assign imm_switch_79_io_in0 = w_internal_174; // @[Benes.scala 109:25]
  assign imm_switch_79_io_in1 = w_internal_255; // @[Benes.scala 118:29]
  assign imm_switch_79_io_sel0 = r_mux_bus_ff_158; // @[Benes.scala 123:26]
  assign imm_switch_79_io_sel1 = r_mux_bus_ff_159; // @[Benes.scala 124:26]
  assign imm_switch_80_io_in0 = w_internal_176; // @[Benes.scala 109:25]
  assign imm_switch_80_io_in1 = w_internal_217; // @[Benes.scala 118:29]
  assign imm_switch_80_io_sel0 = r_mux_bus_ff_160; // @[Benes.scala 123:26]
  assign imm_switch_80_io_sel1 = r_mux_bus_ff_161; // @[Benes.scala 124:26]
  assign imm_switch_81_io_in0 = w_internal_180; // @[Benes.scala 109:25]
  assign imm_switch_81_io_in1 = w_internal_161; // @[Benes.scala 114:29]
  assign imm_switch_81_io_sel0 = r_mux_bus_ff_162; // @[Benes.scala 123:26]
  assign imm_switch_81_io_sel1 = r_mux_bus_ff_163; // @[Benes.scala 124:26]
  assign imm_switch_82_io_in0 = w_internal_182; // @[Benes.scala 109:25]
  assign imm_switch_82_io_in1 = w_internal_223; // @[Benes.scala 112:29]
  assign imm_switch_82_io_sel0 = r_mux_bus_ff_164; // @[Benes.scala 123:26]
  assign imm_switch_82_io_sel1 = r_mux_bus_ff_165; // @[Benes.scala 124:26]
  assign imm_switch_83_io_in0 = w_internal_184; // @[Benes.scala 109:25]
  assign imm_switch_83_io_in1 = w_internal_265; // @[Benes.scala 112:29]
  assign imm_switch_83_io_sel0 = r_mux_bus_ff_166; // @[Benes.scala 123:26]
  assign imm_switch_83_io_sel1 = r_mux_bus_ff_167; // @[Benes.scala 124:26]
  assign imm_switch_84_io_in0 = w_internal_186; // @[Benes.scala 109:25]
  assign imm_switch_84_io_in1 = w_internal_27; // @[Benes.scala 114:29]
  assign imm_switch_84_io_sel0 = r_mux_bus_ff_168; // @[Benes.scala 123:26]
  assign imm_switch_84_io_sel1 = r_mux_bus_ff_169; // @[Benes.scala 124:26]
  assign imm_switch_85_io_in0 = w_internal_188; // @[Benes.scala 109:25]
  assign imm_switch_85_io_in1 = w_internal_509; // @[Benes.scala 112:29]
  assign imm_switch_85_io_sel0 = r_mux_bus_ff_170; // @[Benes.scala 123:26]
  assign imm_switch_85_io_sel1 = r_mux_bus_ff_171; // @[Benes.scala 124:26]
  assign imm_switch_86_io_in0 = w_internal_190; // @[Benes.scala 109:25]
  assign imm_switch_86_io_in1 = w_internal_511; // @[Benes.scala 118:29]
  assign imm_switch_86_io_sel0 = r_mux_bus_ff_172; // @[Benes.scala 123:26]
  assign imm_switch_86_io_sel1 = r_mux_bus_ff_173; // @[Benes.scala 124:26]
  assign imm_switch_87_io_in0 = w_internal_192; // @[Benes.scala 109:25]
  assign imm_switch_87_io_in1 = w_internal_33; // @[Benes.scala 120:29]
  assign imm_switch_87_io_sel0 = r_mux_bus_ff_174; // @[Benes.scala 123:26]
  assign imm_switch_87_io_sel1 = r_mux_bus_ff_175; // @[Benes.scala 124:26]
  assign imm_switch_88_io_in0 = w_internal_194; // @[Benes.scala 109:25]
  assign imm_switch_88_io_in1 = w_internal_275; // @[Benes.scala 118:29]
  assign imm_switch_88_io_sel0 = r_mux_bus_ff_176; // @[Benes.scala 123:26]
  assign imm_switch_88_io_sel1 = r_mux_bus_ff_177; // @[Benes.scala 124:26]
  assign imm_switch_89_io_in0 = w_internal_196; // @[Benes.scala 109:25]
  assign imm_switch_89_io_in1 = w_internal_237; // @[Benes.scala 118:29]
  assign imm_switch_89_io_sel0 = r_mux_bus_ff_178; // @[Benes.scala 123:26]
  assign imm_switch_89_io_sel1 = r_mux_bus_ff_179; // @[Benes.scala 124:26]
  assign imm_switch_90_io_in0 = w_internal_200; // @[Benes.scala 109:25]
  assign imm_switch_90_io_in1 = w_internal_221; // @[Benes.scala 112:29]
  assign imm_switch_90_io_sel0 = r_mux_bus_ff_180; // @[Benes.scala 123:26]
  assign imm_switch_90_io_sel1 = r_mux_bus_ff_181; // @[Benes.scala 124:26]
  assign imm_switch_91_io_in0 = w_internal_202; // @[Benes.scala 109:25]
  assign imm_switch_91_io_in1 = w_internal_163; // @[Benes.scala 114:29]
  assign imm_switch_91_io_sel0 = r_mux_bus_ff_182; // @[Benes.scala 123:26]
  assign imm_switch_91_io_sel1 = r_mux_bus_ff_183; // @[Benes.scala 124:26]
  assign imm_switch_92_io_in0 = w_internal_204; // @[Benes.scala 109:25]
  assign imm_switch_92_io_in1 = w_internal_285; // @[Benes.scala 112:29]
  assign imm_switch_92_io_sel0 = r_mux_bus_ff_184; // @[Benes.scala 123:26]
  assign imm_switch_92_io_sel1 = r_mux_bus_ff_185; // @[Benes.scala 124:26]
  assign imm_switch_93_io_in0 = w_internal_206; // @[Benes.scala 109:25]
  assign imm_switch_93_io_in1 = w_internal_47; // @[Benes.scala 114:29]
  assign imm_switch_93_io_sel0 = r_mux_bus_ff_186; // @[Benes.scala 123:26]
  assign imm_switch_93_io_sel1 = r_mux_bus_ff_187; // @[Benes.scala 124:26]
  assign imm_switch_94_io_in0 = w_internal_208; // @[Benes.scala 109:25]
  assign imm_switch_94_io_in1 = w_internal_529; // @[Benes.scala 112:29]
  assign imm_switch_94_io_sel0 = r_mux_bus_ff_188; // @[Benes.scala 123:26]
  assign imm_switch_94_io_sel1 = r_mux_bus_ff_189; // @[Benes.scala 124:26]
  assign imm_switch_95_io_in0 = w_internal_210; // @[Benes.scala 109:25]
  assign imm_switch_95_io_in1 = w_internal_531; // @[Benes.scala 118:29]
  assign imm_switch_95_io_sel0 = r_mux_bus_ff_190; // @[Benes.scala 123:26]
  assign imm_switch_95_io_sel1 = r_mux_bus_ff_191; // @[Benes.scala 124:26]
  assign imm_switch_96_io_in0 = w_internal_212; // @[Benes.scala 109:25]
  assign imm_switch_96_io_in1 = w_internal_53; // @[Benes.scala 120:29]
  assign imm_switch_96_io_sel0 = r_mux_bus_ff_192; // @[Benes.scala 123:26]
  assign imm_switch_96_io_sel1 = r_mux_bus_ff_193; // @[Benes.scala 124:26]
  assign imm_switch_97_io_in0 = w_internal_214; // @[Benes.scala 109:25]
  assign imm_switch_97_io_in1 = w_internal_295; // @[Benes.scala 118:29]
  assign imm_switch_97_io_sel0 = r_mux_bus_ff_194; // @[Benes.scala 123:26]
  assign imm_switch_97_io_sel1 = r_mux_bus_ff_195; // @[Benes.scala 124:26]
  assign imm_switch_98_io_in0 = w_internal_216; // @[Benes.scala 109:25]
  assign imm_switch_98_io_in1 = w_internal_177; // @[Benes.scala 120:29]
  assign imm_switch_98_io_sel0 = r_mux_bus_ff_196; // @[Benes.scala 123:26]
  assign imm_switch_98_io_sel1 = r_mux_bus_ff_197; // @[Benes.scala 124:26]
  assign imm_switch_99_io_in0 = w_internal_220; // @[Benes.scala 109:25]
  assign imm_switch_99_io_in1 = w_internal_201; // @[Benes.scala 114:29]
  assign imm_switch_99_io_sel0 = r_mux_bus_ff_198; // @[Benes.scala 123:26]
  assign imm_switch_99_io_sel1 = r_mux_bus_ff_199; // @[Benes.scala 124:26]
  assign imm_switch_100_io_in0 = w_internal_222; // @[Benes.scala 109:25]
  assign imm_switch_100_io_in1 = w_internal_183; // @[Benes.scala 114:29]
  assign imm_switch_100_io_sel0 = r_mux_bus_ff_200; // @[Benes.scala 123:26]
  assign imm_switch_100_io_sel1 = r_mux_bus_ff_201; // @[Benes.scala 124:26]
  assign imm_switch_101_io_in0 = w_internal_224; // @[Benes.scala 109:25]
  assign imm_switch_101_io_in1 = w_internal_305; // @[Benes.scala 112:29]
  assign imm_switch_101_io_sel0 = r_mux_bus_ff_202; // @[Benes.scala 123:26]
  assign imm_switch_101_io_sel1 = r_mux_bus_ff_203; // @[Benes.scala 124:26]
  assign imm_switch_102_io_in0 = w_internal_226; // @[Benes.scala 109:25]
  assign imm_switch_102_io_in1 = w_internal_67; // @[Benes.scala 114:29]
  assign imm_switch_102_io_sel0 = r_mux_bus_ff_204; // @[Benes.scala 123:26]
  assign imm_switch_102_io_sel1 = r_mux_bus_ff_205; // @[Benes.scala 124:26]
  assign imm_switch_103_io_in0 = w_internal_228; // @[Benes.scala 109:25]
  assign imm_switch_103_io_in1 = w_internal_549; // @[Benes.scala 112:29]
  assign imm_switch_103_io_sel0 = r_mux_bus_ff_206; // @[Benes.scala 123:26]
  assign imm_switch_103_io_sel1 = r_mux_bus_ff_207; // @[Benes.scala 124:26]
  assign imm_switch_104_io_in0 = w_internal_230; // @[Benes.scala 109:25]
  assign imm_switch_104_io_in1 = w_internal_551; // @[Benes.scala 118:29]
  assign imm_switch_104_io_sel0 = r_mux_bus_ff_208; // @[Benes.scala 123:26]
  assign imm_switch_104_io_sel1 = r_mux_bus_ff_209; // @[Benes.scala 124:26]
  assign imm_switch_105_io_in0 = w_internal_232; // @[Benes.scala 109:25]
  assign imm_switch_105_io_in1 = w_internal_73; // @[Benes.scala 120:29]
  assign imm_switch_105_io_sel0 = r_mux_bus_ff_210; // @[Benes.scala 123:26]
  assign imm_switch_105_io_sel1 = r_mux_bus_ff_211; // @[Benes.scala 124:26]
  assign imm_switch_106_io_in0 = w_internal_234; // @[Benes.scala 109:25]
  assign imm_switch_106_io_in1 = w_internal_315; // @[Benes.scala 118:29]
  assign imm_switch_106_io_sel0 = r_mux_bus_ff_212; // @[Benes.scala 123:26]
  assign imm_switch_106_io_sel1 = r_mux_bus_ff_213; // @[Benes.scala 124:26]
  assign imm_switch_107_io_in0 = w_internal_236; // @[Benes.scala 109:25]
  assign imm_switch_107_io_in1 = w_internal_197; // @[Benes.scala 120:29]
  assign imm_switch_107_io_sel0 = r_mux_bus_ff_214; // @[Benes.scala 123:26]
  assign imm_switch_107_io_sel1 = r_mux_bus_ff_215; // @[Benes.scala 124:26]
  assign imm_switch_108_io_in0 = w_internal_240; // @[Benes.scala 109:25]
  assign imm_switch_108_io_in1 = w_internal_261; // @[Benes.scala 112:29]
  assign imm_switch_108_io_sel0 = r_mux_bus_ff_216; // @[Benes.scala 123:26]
  assign imm_switch_108_io_sel1 = r_mux_bus_ff_217; // @[Benes.scala 124:26]
  assign imm_switch_109_io_in0 = w_internal_242; // @[Benes.scala 109:25]
  assign imm_switch_109_io_in1 = w_internal_283; // @[Benes.scala 112:29]
  assign imm_switch_109_io_sel0 = r_mux_bus_ff_218; // @[Benes.scala 123:26]
  assign imm_switch_109_io_sel1 = r_mux_bus_ff_219; // @[Benes.scala 124:26]
  assign imm_switch_110_io_in0 = w_internal_244; // @[Benes.scala 109:25]
  assign imm_switch_110_io_in1 = w_internal_165; // @[Benes.scala 114:29]
  assign imm_switch_110_io_sel0 = r_mux_bus_ff_220; // @[Benes.scala 123:26]
  assign imm_switch_110_io_sel1 = r_mux_bus_ff_221; // @[Benes.scala 124:26]
  assign imm_switch_111_io_in0 = w_internal_246; // @[Benes.scala 109:25]
  assign imm_switch_111_io_in1 = w_internal_87; // @[Benes.scala 114:29]
  assign imm_switch_111_io_sel0 = r_mux_bus_ff_222; // @[Benes.scala 123:26]
  assign imm_switch_111_io_sel1 = r_mux_bus_ff_223; // @[Benes.scala 124:26]
  assign imm_switch_112_io_in0 = w_internal_248; // @[Benes.scala 109:25]
  assign imm_switch_112_io_in1 = w_internal_569; // @[Benes.scala 112:29]
  assign imm_switch_112_io_sel0 = r_mux_bus_ff_224; // @[Benes.scala 123:26]
  assign imm_switch_112_io_sel1 = r_mux_bus_ff_225; // @[Benes.scala 124:26]
  assign imm_switch_113_io_in0 = w_internal_250; // @[Benes.scala 109:25]
  assign imm_switch_113_io_in1 = w_internal_571; // @[Benes.scala 118:29]
  assign imm_switch_113_io_sel0 = r_mux_bus_ff_226; // @[Benes.scala 123:26]
  assign imm_switch_113_io_sel1 = r_mux_bus_ff_227; // @[Benes.scala 124:26]
  assign imm_switch_114_io_in0 = w_internal_252; // @[Benes.scala 109:25]
  assign imm_switch_114_io_in1 = w_internal_93; // @[Benes.scala 120:29]
  assign imm_switch_114_io_sel0 = r_mux_bus_ff_228; // @[Benes.scala 123:26]
  assign imm_switch_114_io_sel1 = r_mux_bus_ff_229; // @[Benes.scala 124:26]
  assign imm_switch_115_io_in0 = w_internal_254; // @[Benes.scala 109:25]
  assign imm_switch_115_io_in1 = w_internal_175; // @[Benes.scala 120:29]
  assign imm_switch_115_io_sel0 = r_mux_bus_ff_230; // @[Benes.scala 123:26]
  assign imm_switch_115_io_sel1 = r_mux_bus_ff_231; // @[Benes.scala 124:26]
  assign imm_switch_116_io_in0 = w_internal_256; // @[Benes.scala 109:25]
  assign imm_switch_116_io_in1 = w_internal_297; // @[Benes.scala 118:29]
  assign imm_switch_116_io_sel0 = r_mux_bus_ff_232; // @[Benes.scala 123:26]
  assign imm_switch_116_io_sel1 = r_mux_bus_ff_233; // @[Benes.scala 124:26]
  assign imm_switch_117_io_in0 = w_internal_260; // @[Benes.scala 109:25]
  assign imm_switch_117_io_in1 = w_internal_241; // @[Benes.scala 114:29]
  assign imm_switch_117_io_sel0 = r_mux_bus_ff_234; // @[Benes.scala 123:26]
  assign imm_switch_117_io_sel1 = r_mux_bus_ff_235; // @[Benes.scala 124:26]
  assign imm_switch_118_io_in0 = w_internal_262; // @[Benes.scala 109:25]
  assign imm_switch_118_io_in1 = w_internal_303; // @[Benes.scala 112:29]
  assign imm_switch_118_io_sel0 = r_mux_bus_ff_236; // @[Benes.scala 123:26]
  assign imm_switch_118_io_sel1 = r_mux_bus_ff_237; // @[Benes.scala 124:26]
  assign imm_switch_119_io_in0 = w_internal_264; // @[Benes.scala 109:25]
  assign imm_switch_119_io_in1 = w_internal_185; // @[Benes.scala 114:29]
  assign imm_switch_119_io_sel0 = r_mux_bus_ff_238; // @[Benes.scala 123:26]
  assign imm_switch_119_io_sel1 = r_mux_bus_ff_239; // @[Benes.scala 124:26]
  assign imm_switch_120_io_in0 = w_internal_266; // @[Benes.scala 109:25]
  assign imm_switch_120_io_in1 = w_internal_107; // @[Benes.scala 114:29]
  assign imm_switch_120_io_sel0 = r_mux_bus_ff_240; // @[Benes.scala 123:26]
  assign imm_switch_120_io_sel1 = r_mux_bus_ff_241; // @[Benes.scala 124:26]
  assign imm_switch_121_io_in0 = w_internal_268; // @[Benes.scala 109:25]
  assign imm_switch_121_io_in1 = w_internal_589; // @[Benes.scala 112:29]
  assign imm_switch_121_io_sel0 = r_mux_bus_ff_242; // @[Benes.scala 123:26]
  assign imm_switch_121_io_sel1 = r_mux_bus_ff_243; // @[Benes.scala 124:26]
  assign imm_switch_122_io_in0 = w_internal_270; // @[Benes.scala 109:25]
  assign imm_switch_122_io_in1 = w_internal_591; // @[Benes.scala 118:29]
  assign imm_switch_122_io_sel0 = r_mux_bus_ff_244; // @[Benes.scala 123:26]
  assign imm_switch_122_io_sel1 = r_mux_bus_ff_245; // @[Benes.scala 124:26]
  assign imm_switch_123_io_in0 = w_internal_272; // @[Benes.scala 109:25]
  assign imm_switch_123_io_in1 = w_internal_113; // @[Benes.scala 120:29]
  assign imm_switch_123_io_sel0 = r_mux_bus_ff_246; // @[Benes.scala 123:26]
  assign imm_switch_123_io_sel1 = r_mux_bus_ff_247; // @[Benes.scala 124:26]
  assign imm_switch_124_io_in0 = w_internal_274; // @[Benes.scala 109:25]
  assign imm_switch_124_io_in1 = w_internal_195; // @[Benes.scala 120:29]
  assign imm_switch_124_io_sel0 = r_mux_bus_ff_248; // @[Benes.scala 123:26]
  assign imm_switch_124_io_sel1 = r_mux_bus_ff_249; // @[Benes.scala 124:26]
  assign imm_switch_125_io_in0 = w_internal_276; // @[Benes.scala 109:25]
  assign imm_switch_125_io_in1 = w_internal_317; // @[Benes.scala 118:29]
  assign imm_switch_125_io_sel0 = r_mux_bus_ff_250; // @[Benes.scala 123:26]
  assign imm_switch_125_io_sel1 = r_mux_bus_ff_251; // @[Benes.scala 124:26]
  assign imm_switch_126_io_in0 = w_internal_280; // @[Benes.scala 109:25]
  assign imm_switch_126_io_in1 = w_internal_301; // @[Benes.scala 112:29]
  assign imm_switch_126_io_sel0 = r_mux_bus_ff_252; // @[Benes.scala 123:26]
  assign imm_switch_126_io_sel1 = r_mux_bus_ff_253; // @[Benes.scala 124:26]
  assign imm_switch_127_io_in0 = w_internal_282; // @[Benes.scala 109:25]
  assign imm_switch_127_io_in1 = w_internal_243; // @[Benes.scala 114:29]
  assign imm_switch_127_io_sel0 = r_mux_bus_ff_254; // @[Benes.scala 123:26]
  assign imm_switch_127_io_sel1 = r_mux_bus_ff_255; // @[Benes.scala 124:26]
  assign imm_switch_128_io_in0 = w_internal_284; // @[Benes.scala 109:25]
  assign imm_switch_128_io_in1 = w_internal_205; // @[Benes.scala 114:29]
  assign imm_switch_128_io_sel0 = r_mux_bus_ff_256; // @[Benes.scala 123:26]
  assign imm_switch_128_io_sel1 = r_mux_bus_ff_257; // @[Benes.scala 124:26]
  assign imm_switch_129_io_in0 = w_internal_286; // @[Benes.scala 109:25]
  assign imm_switch_129_io_in1 = w_internal_127; // @[Benes.scala 114:29]
  assign imm_switch_129_io_sel0 = r_mux_bus_ff_258; // @[Benes.scala 123:26]
  assign imm_switch_129_io_sel1 = r_mux_bus_ff_259; // @[Benes.scala 124:26]
  assign imm_switch_130_io_in0 = w_internal_288; // @[Benes.scala 109:25]
  assign imm_switch_130_io_in1 = w_internal_609; // @[Benes.scala 112:29]
  assign imm_switch_130_io_sel0 = r_mux_bus_ff_260; // @[Benes.scala 123:26]
  assign imm_switch_130_io_sel1 = r_mux_bus_ff_261; // @[Benes.scala 124:26]
  assign imm_switch_131_io_in0 = w_internal_290; // @[Benes.scala 109:25]
  assign imm_switch_131_io_in1 = w_internal_611; // @[Benes.scala 118:29]
  assign imm_switch_131_io_sel0 = r_mux_bus_ff_262; // @[Benes.scala 123:26]
  assign imm_switch_131_io_sel1 = r_mux_bus_ff_263; // @[Benes.scala 124:26]
  assign imm_switch_132_io_in0 = w_internal_292; // @[Benes.scala 109:25]
  assign imm_switch_132_io_in1 = w_internal_133; // @[Benes.scala 120:29]
  assign imm_switch_132_io_sel0 = r_mux_bus_ff_264; // @[Benes.scala 123:26]
  assign imm_switch_132_io_sel1 = r_mux_bus_ff_265; // @[Benes.scala 124:26]
  assign imm_switch_133_io_in0 = w_internal_294; // @[Benes.scala 109:25]
  assign imm_switch_133_io_in1 = w_internal_215; // @[Benes.scala 120:29]
  assign imm_switch_133_io_sel0 = r_mux_bus_ff_266; // @[Benes.scala 123:26]
  assign imm_switch_133_io_sel1 = r_mux_bus_ff_267; // @[Benes.scala 124:26]
  assign imm_switch_134_io_in0 = w_internal_296; // @[Benes.scala 109:25]
  assign imm_switch_134_io_in1 = w_internal_257; // @[Benes.scala 120:29]
  assign imm_switch_134_io_sel0 = r_mux_bus_ff_268; // @[Benes.scala 123:26]
  assign imm_switch_134_io_sel1 = r_mux_bus_ff_269; // @[Benes.scala 124:26]
  assign imm_switch_135_io_in0 = w_internal_300; // @[Benes.scala 109:25]
  assign imm_switch_135_io_in1 = w_internal_281; // @[Benes.scala 114:29]
  assign imm_switch_135_io_sel0 = r_mux_bus_ff_270; // @[Benes.scala 123:26]
  assign imm_switch_135_io_sel1 = r_mux_bus_ff_271; // @[Benes.scala 124:26]
  assign imm_switch_136_io_in0 = w_internal_302; // @[Benes.scala 109:25]
  assign imm_switch_136_io_in1 = w_internal_263; // @[Benes.scala 114:29]
  assign imm_switch_136_io_sel0 = r_mux_bus_ff_272; // @[Benes.scala 123:26]
  assign imm_switch_136_io_sel1 = r_mux_bus_ff_273; // @[Benes.scala 124:26]
  assign imm_switch_137_io_in0 = w_internal_304; // @[Benes.scala 109:25]
  assign imm_switch_137_io_in1 = w_internal_225; // @[Benes.scala 114:29]
  assign imm_switch_137_io_sel0 = r_mux_bus_ff_274; // @[Benes.scala 123:26]
  assign imm_switch_137_io_sel1 = r_mux_bus_ff_275; // @[Benes.scala 124:26]
  assign imm_switch_138_io_in0 = w_internal_306; // @[Benes.scala 109:25]
  assign imm_switch_138_io_in1 = w_internal_147; // @[Benes.scala 114:29]
  assign imm_switch_138_io_sel0 = r_mux_bus_ff_276; // @[Benes.scala 123:26]
  assign imm_switch_138_io_sel1 = r_mux_bus_ff_277; // @[Benes.scala 124:26]
  assign imm_switch_139_io_in0 = w_internal_308; // @[Benes.scala 109:25]
  assign imm_switch_139_io_in1 = w_internal_629; // @[Benes.scala 112:29]
  assign imm_switch_139_io_sel0 = r_mux_bus_ff_278; // @[Benes.scala 123:26]
  assign imm_switch_139_io_sel1 = r_mux_bus_ff_279; // @[Benes.scala 124:26]
  assign imm_switch_140_io_in0 = w_internal_310; // @[Benes.scala 109:25]
  assign imm_switch_140_io_in1 = w_internal_631; // @[Benes.scala 118:29]
  assign imm_switch_140_io_sel0 = r_mux_bus_ff_280; // @[Benes.scala 123:26]
  assign imm_switch_140_io_sel1 = r_mux_bus_ff_281; // @[Benes.scala 124:26]
  assign imm_switch_141_io_in0 = w_internal_312; // @[Benes.scala 109:25]
  assign imm_switch_141_io_in1 = w_internal_153; // @[Benes.scala 120:29]
  assign imm_switch_141_io_sel0 = r_mux_bus_ff_282; // @[Benes.scala 123:26]
  assign imm_switch_141_io_sel1 = r_mux_bus_ff_283; // @[Benes.scala 124:26]
  assign imm_switch_142_io_in0 = w_internal_314; // @[Benes.scala 109:25]
  assign imm_switch_142_io_in1 = w_internal_235; // @[Benes.scala 120:29]
  assign imm_switch_142_io_sel0 = r_mux_bus_ff_284; // @[Benes.scala 123:26]
  assign imm_switch_142_io_sel1 = r_mux_bus_ff_285; // @[Benes.scala 124:26]
  assign imm_switch_143_io_in0 = w_internal_316; // @[Benes.scala 109:25]
  assign imm_switch_143_io_in1 = w_internal_277; // @[Benes.scala 120:29]
  assign imm_switch_143_io_sel0 = r_mux_bus_ff_286; // @[Benes.scala 123:26]
  assign imm_switch_143_io_sel1 = r_mux_bus_ff_287; // @[Benes.scala 124:26]
  assign imm_switch_144_io_in0 = w_internal_320; // @[Benes.scala 109:25]
  assign imm_switch_144_io_in1 = w_internal_341; // @[Benes.scala 112:29]
  assign imm_switch_144_io_sel0 = r_mux_bus_ff_288; // @[Benes.scala 123:26]
  assign imm_switch_144_io_sel1 = r_mux_bus_ff_289; // @[Benes.scala 124:26]
  assign imm_switch_145_io_in0 = w_internal_322; // @[Benes.scala 109:25]
  assign imm_switch_145_io_in1 = w_internal_363; // @[Benes.scala 112:29]
  assign imm_switch_145_io_sel0 = r_mux_bus_ff_290; // @[Benes.scala 123:26]
  assign imm_switch_145_io_sel1 = r_mux_bus_ff_291; // @[Benes.scala 124:26]
  assign imm_switch_146_io_in0 = w_internal_324; // @[Benes.scala 109:25]
  assign imm_switch_146_io_in1 = w_internal_405; // @[Benes.scala 112:29]
  assign imm_switch_146_io_sel0 = r_mux_bus_ff_292; // @[Benes.scala 123:26]
  assign imm_switch_146_io_sel1 = r_mux_bus_ff_293; // @[Benes.scala 124:26]
  assign imm_switch_147_io_in0 = w_internal_326; // @[Benes.scala 109:25]
  assign imm_switch_147_io_in1 = w_internal_487; // @[Benes.scala 112:29]
  assign imm_switch_147_io_sel0 = r_mux_bus_ff_294; // @[Benes.scala 123:26]
  assign imm_switch_147_io_sel1 = r_mux_bus_ff_295; // @[Benes.scala 124:26]
  assign imm_switch_148_io_in0 = w_internal_328; // @[Benes.scala 109:25]
  assign imm_switch_148_io_in1 = w_internal_9; // @[Benes.scala 114:29]
  assign imm_switch_148_io_sel0 = r_mux_bus_ff_296; // @[Benes.scala 123:26]
  assign imm_switch_148_io_sel1 = r_mux_bus_ff_297; // @[Benes.scala 124:26]
  assign imm_switch_149_io_in0 = w_internal_330; // @[Benes.scala 109:25]
  assign imm_switch_149_io_in1 = w_internal_11; // @[Benes.scala 120:29]
  assign imm_switch_149_io_sel0 = r_mux_bus_ff_298; // @[Benes.scala 123:26]
  assign imm_switch_149_io_sel1 = r_mux_bus_ff_299; // @[Benes.scala 124:26]
  assign imm_switch_150_io_in0 = w_internal_332; // @[Benes.scala 109:25]
  assign imm_switch_150_io_in1 = w_internal_493; // @[Benes.scala 118:29]
  assign imm_switch_150_io_sel0 = r_mux_bus_ff_300; // @[Benes.scala 123:26]
  assign imm_switch_150_io_sel1 = r_mux_bus_ff_301; // @[Benes.scala 124:26]
  assign imm_switch_151_io_in0 = w_internal_334; // @[Benes.scala 109:25]
  assign imm_switch_151_io_in1 = w_internal_415; // @[Benes.scala 118:29]
  assign imm_switch_151_io_sel0 = r_mux_bus_ff_302; // @[Benes.scala 123:26]
  assign imm_switch_151_io_sel1 = r_mux_bus_ff_303; // @[Benes.scala 124:26]
  assign imm_switch_152_io_in0 = w_internal_336; // @[Benes.scala 109:25]
  assign imm_switch_152_io_in1 = w_internal_377; // @[Benes.scala 118:29]
  assign imm_switch_152_io_sel0 = r_mux_bus_ff_304; // @[Benes.scala 123:26]
  assign imm_switch_152_io_sel1 = r_mux_bus_ff_305; // @[Benes.scala 124:26]
  assign imm_switch_153_io_in0 = w_internal_340; // @[Benes.scala 109:25]
  assign imm_switch_153_io_in1 = w_internal_321; // @[Benes.scala 114:29]
  assign imm_switch_153_io_sel0 = r_mux_bus_ff_306; // @[Benes.scala 123:26]
  assign imm_switch_153_io_sel1 = r_mux_bus_ff_307; // @[Benes.scala 124:26]
  assign imm_switch_154_io_in0 = w_internal_342; // @[Benes.scala 109:25]
  assign imm_switch_154_io_in1 = w_internal_383; // @[Benes.scala 112:29]
  assign imm_switch_154_io_sel0 = r_mux_bus_ff_308; // @[Benes.scala 123:26]
  assign imm_switch_154_io_sel1 = r_mux_bus_ff_309; // @[Benes.scala 124:26]
  assign imm_switch_155_io_in0 = w_internal_344; // @[Benes.scala 109:25]
  assign imm_switch_155_io_in1 = w_internal_425; // @[Benes.scala 112:29]
  assign imm_switch_155_io_sel0 = r_mux_bus_ff_310; // @[Benes.scala 123:26]
  assign imm_switch_155_io_sel1 = r_mux_bus_ff_311; // @[Benes.scala 124:26]
  assign imm_switch_156_io_in0 = w_internal_346; // @[Benes.scala 109:25]
  assign imm_switch_156_io_in1 = w_internal_507; // @[Benes.scala 112:29]
  assign imm_switch_156_io_sel0 = r_mux_bus_ff_312; // @[Benes.scala 123:26]
  assign imm_switch_156_io_sel1 = r_mux_bus_ff_313; // @[Benes.scala 124:26]
  assign imm_switch_157_io_in0 = w_internal_348; // @[Benes.scala 109:25]
  assign imm_switch_157_io_in1 = w_internal_29; // @[Benes.scala 114:29]
  assign imm_switch_157_io_sel0 = r_mux_bus_ff_314; // @[Benes.scala 123:26]
  assign imm_switch_157_io_sel1 = r_mux_bus_ff_315; // @[Benes.scala 124:26]
  assign imm_switch_158_io_in0 = w_internal_350; // @[Benes.scala 109:25]
  assign imm_switch_158_io_in1 = w_internal_31; // @[Benes.scala 120:29]
  assign imm_switch_158_io_sel0 = r_mux_bus_ff_316; // @[Benes.scala 123:26]
  assign imm_switch_158_io_sel1 = r_mux_bus_ff_317; // @[Benes.scala 124:26]
  assign imm_switch_159_io_in0 = w_internal_352; // @[Benes.scala 109:25]
  assign imm_switch_159_io_in1 = w_internal_513; // @[Benes.scala 118:29]
  assign imm_switch_159_io_sel0 = r_mux_bus_ff_318; // @[Benes.scala 123:26]
  assign imm_switch_159_io_sel1 = r_mux_bus_ff_319; // @[Benes.scala 124:26]
  assign imm_switch_160_io_in0 = w_internal_354; // @[Benes.scala 109:25]
  assign imm_switch_160_io_in1 = w_internal_435; // @[Benes.scala 118:29]
  assign imm_switch_160_io_sel0 = r_mux_bus_ff_320; // @[Benes.scala 123:26]
  assign imm_switch_160_io_sel1 = r_mux_bus_ff_321; // @[Benes.scala 124:26]
  assign imm_switch_161_io_in0 = w_internal_356; // @[Benes.scala 109:25]
  assign imm_switch_161_io_in1 = w_internal_397; // @[Benes.scala 118:29]
  assign imm_switch_161_io_sel0 = r_mux_bus_ff_322; // @[Benes.scala 123:26]
  assign imm_switch_161_io_sel1 = r_mux_bus_ff_323; // @[Benes.scala 124:26]
  assign imm_switch_162_io_in0 = w_internal_360; // @[Benes.scala 109:25]
  assign imm_switch_162_io_in1 = w_internal_381; // @[Benes.scala 112:29]
  assign imm_switch_162_io_sel0 = r_mux_bus_ff_324; // @[Benes.scala 123:26]
  assign imm_switch_162_io_sel1 = r_mux_bus_ff_325; // @[Benes.scala 124:26]
  assign imm_switch_163_io_in0 = w_internal_362; // @[Benes.scala 109:25]
  assign imm_switch_163_io_in1 = w_internal_323; // @[Benes.scala 114:29]
  assign imm_switch_163_io_sel0 = r_mux_bus_ff_326; // @[Benes.scala 123:26]
  assign imm_switch_163_io_sel1 = r_mux_bus_ff_327; // @[Benes.scala 124:26]
  assign imm_switch_164_io_in0 = w_internal_364; // @[Benes.scala 109:25]
  assign imm_switch_164_io_in1 = w_internal_445; // @[Benes.scala 112:29]
  assign imm_switch_164_io_sel0 = r_mux_bus_ff_328; // @[Benes.scala 123:26]
  assign imm_switch_164_io_sel1 = r_mux_bus_ff_329; // @[Benes.scala 124:26]
  assign imm_switch_165_io_in0 = w_internal_366; // @[Benes.scala 109:25]
  assign imm_switch_165_io_in1 = w_internal_527; // @[Benes.scala 112:29]
  assign imm_switch_165_io_sel0 = r_mux_bus_ff_330; // @[Benes.scala 123:26]
  assign imm_switch_165_io_sel1 = r_mux_bus_ff_331; // @[Benes.scala 124:26]
  assign imm_switch_166_io_in0 = w_internal_368; // @[Benes.scala 109:25]
  assign imm_switch_166_io_in1 = w_internal_49; // @[Benes.scala 114:29]
  assign imm_switch_166_io_sel0 = r_mux_bus_ff_332; // @[Benes.scala 123:26]
  assign imm_switch_166_io_sel1 = r_mux_bus_ff_333; // @[Benes.scala 124:26]
  assign imm_switch_167_io_in0 = w_internal_370; // @[Benes.scala 109:25]
  assign imm_switch_167_io_in1 = w_internal_51; // @[Benes.scala 120:29]
  assign imm_switch_167_io_sel0 = r_mux_bus_ff_334; // @[Benes.scala 123:26]
  assign imm_switch_167_io_sel1 = r_mux_bus_ff_335; // @[Benes.scala 124:26]
  assign imm_switch_168_io_in0 = w_internal_372; // @[Benes.scala 109:25]
  assign imm_switch_168_io_in1 = w_internal_533; // @[Benes.scala 118:29]
  assign imm_switch_168_io_sel0 = r_mux_bus_ff_336; // @[Benes.scala 123:26]
  assign imm_switch_168_io_sel1 = r_mux_bus_ff_337; // @[Benes.scala 124:26]
  assign imm_switch_169_io_in0 = w_internal_374; // @[Benes.scala 109:25]
  assign imm_switch_169_io_in1 = w_internal_455; // @[Benes.scala 118:29]
  assign imm_switch_169_io_sel0 = r_mux_bus_ff_338; // @[Benes.scala 123:26]
  assign imm_switch_169_io_sel1 = r_mux_bus_ff_339; // @[Benes.scala 124:26]
  assign imm_switch_170_io_in0 = w_internal_376; // @[Benes.scala 109:25]
  assign imm_switch_170_io_in1 = w_internal_337; // @[Benes.scala 120:29]
  assign imm_switch_170_io_sel0 = r_mux_bus_ff_340; // @[Benes.scala 123:26]
  assign imm_switch_170_io_sel1 = r_mux_bus_ff_341; // @[Benes.scala 124:26]
  assign imm_switch_171_io_in0 = w_internal_380; // @[Benes.scala 109:25]
  assign imm_switch_171_io_in1 = w_internal_361; // @[Benes.scala 114:29]
  assign imm_switch_171_io_sel0 = r_mux_bus_ff_342; // @[Benes.scala 123:26]
  assign imm_switch_171_io_sel1 = r_mux_bus_ff_343; // @[Benes.scala 124:26]
  assign imm_switch_172_io_in0 = w_internal_382; // @[Benes.scala 109:25]
  assign imm_switch_172_io_in1 = w_internal_343; // @[Benes.scala 114:29]
  assign imm_switch_172_io_sel0 = r_mux_bus_ff_344; // @[Benes.scala 123:26]
  assign imm_switch_172_io_sel1 = r_mux_bus_ff_345; // @[Benes.scala 124:26]
  assign imm_switch_173_io_in0 = w_internal_384; // @[Benes.scala 109:25]
  assign imm_switch_173_io_in1 = w_internal_465; // @[Benes.scala 112:29]
  assign imm_switch_173_io_sel0 = r_mux_bus_ff_346; // @[Benes.scala 123:26]
  assign imm_switch_173_io_sel1 = r_mux_bus_ff_347; // @[Benes.scala 124:26]
  assign imm_switch_174_io_in0 = w_internal_386; // @[Benes.scala 109:25]
  assign imm_switch_174_io_in1 = w_internal_547; // @[Benes.scala 112:29]
  assign imm_switch_174_io_sel0 = r_mux_bus_ff_348; // @[Benes.scala 123:26]
  assign imm_switch_174_io_sel1 = r_mux_bus_ff_349; // @[Benes.scala 124:26]
  assign imm_switch_175_io_in0 = w_internal_388; // @[Benes.scala 109:25]
  assign imm_switch_175_io_in1 = w_internal_69; // @[Benes.scala 114:29]
  assign imm_switch_175_io_sel0 = r_mux_bus_ff_350; // @[Benes.scala 123:26]
  assign imm_switch_175_io_sel1 = r_mux_bus_ff_351; // @[Benes.scala 124:26]
  assign imm_switch_176_io_in0 = w_internal_390; // @[Benes.scala 109:25]
  assign imm_switch_176_io_in1 = w_internal_71; // @[Benes.scala 120:29]
  assign imm_switch_176_io_sel0 = r_mux_bus_ff_352; // @[Benes.scala 123:26]
  assign imm_switch_176_io_sel1 = r_mux_bus_ff_353; // @[Benes.scala 124:26]
  assign imm_switch_177_io_in0 = w_internal_392; // @[Benes.scala 109:25]
  assign imm_switch_177_io_in1 = w_internal_553; // @[Benes.scala 118:29]
  assign imm_switch_177_io_sel0 = r_mux_bus_ff_354; // @[Benes.scala 123:26]
  assign imm_switch_177_io_sel1 = r_mux_bus_ff_355; // @[Benes.scala 124:26]
  assign imm_switch_178_io_in0 = w_internal_394; // @[Benes.scala 109:25]
  assign imm_switch_178_io_in1 = w_internal_475; // @[Benes.scala 118:29]
  assign imm_switch_178_io_sel0 = r_mux_bus_ff_356; // @[Benes.scala 123:26]
  assign imm_switch_178_io_sel1 = r_mux_bus_ff_357; // @[Benes.scala 124:26]
  assign imm_switch_179_io_in0 = w_internal_396; // @[Benes.scala 109:25]
  assign imm_switch_179_io_in1 = w_internal_357; // @[Benes.scala 120:29]
  assign imm_switch_179_io_sel0 = r_mux_bus_ff_358; // @[Benes.scala 123:26]
  assign imm_switch_179_io_sel1 = r_mux_bus_ff_359; // @[Benes.scala 124:26]
  assign imm_switch_180_io_in0 = w_internal_400; // @[Benes.scala 109:25]
  assign imm_switch_180_io_in1 = w_internal_421; // @[Benes.scala 112:29]
  assign imm_switch_180_io_sel0 = r_mux_bus_ff_360; // @[Benes.scala 123:26]
  assign imm_switch_180_io_sel1 = r_mux_bus_ff_361; // @[Benes.scala 124:26]
  assign imm_switch_181_io_in0 = w_internal_402; // @[Benes.scala 109:25]
  assign imm_switch_181_io_in1 = w_internal_443; // @[Benes.scala 112:29]
  assign imm_switch_181_io_sel0 = r_mux_bus_ff_362; // @[Benes.scala 123:26]
  assign imm_switch_181_io_sel1 = r_mux_bus_ff_363; // @[Benes.scala 124:26]
  assign imm_switch_182_io_in0 = w_internal_404; // @[Benes.scala 109:25]
  assign imm_switch_182_io_in1 = w_internal_325; // @[Benes.scala 114:29]
  assign imm_switch_182_io_sel0 = r_mux_bus_ff_364; // @[Benes.scala 123:26]
  assign imm_switch_182_io_sel1 = r_mux_bus_ff_365; // @[Benes.scala 124:26]
  assign imm_switch_183_io_in0 = w_internal_406; // @[Benes.scala 109:25]
  assign imm_switch_183_io_in1 = w_internal_567; // @[Benes.scala 112:29]
  assign imm_switch_183_io_sel0 = r_mux_bus_ff_366; // @[Benes.scala 123:26]
  assign imm_switch_183_io_sel1 = r_mux_bus_ff_367; // @[Benes.scala 124:26]
  assign imm_switch_184_io_in0 = w_internal_408; // @[Benes.scala 109:25]
  assign imm_switch_184_io_in1 = w_internal_89; // @[Benes.scala 114:29]
  assign imm_switch_184_io_sel0 = r_mux_bus_ff_368; // @[Benes.scala 123:26]
  assign imm_switch_184_io_sel1 = r_mux_bus_ff_369; // @[Benes.scala 124:26]
  assign imm_switch_185_io_in0 = w_internal_410; // @[Benes.scala 109:25]
  assign imm_switch_185_io_in1 = w_internal_91; // @[Benes.scala 120:29]
  assign imm_switch_185_io_sel0 = r_mux_bus_ff_370; // @[Benes.scala 123:26]
  assign imm_switch_185_io_sel1 = r_mux_bus_ff_371; // @[Benes.scala 124:26]
  assign imm_switch_186_io_in0 = w_internal_412; // @[Benes.scala 109:25]
  assign imm_switch_186_io_in1 = w_internal_573; // @[Benes.scala 118:29]
  assign imm_switch_186_io_sel0 = r_mux_bus_ff_372; // @[Benes.scala 123:26]
  assign imm_switch_186_io_sel1 = r_mux_bus_ff_373; // @[Benes.scala 124:26]
  assign imm_switch_187_io_in0 = w_internal_414; // @[Benes.scala 109:25]
  assign imm_switch_187_io_in1 = w_internal_335; // @[Benes.scala 120:29]
  assign imm_switch_187_io_sel0 = r_mux_bus_ff_374; // @[Benes.scala 123:26]
  assign imm_switch_187_io_sel1 = r_mux_bus_ff_375; // @[Benes.scala 124:26]
  assign imm_switch_188_io_in0 = w_internal_416; // @[Benes.scala 109:25]
  assign imm_switch_188_io_in1 = w_internal_457; // @[Benes.scala 118:29]
  assign imm_switch_188_io_sel0 = r_mux_bus_ff_376; // @[Benes.scala 123:26]
  assign imm_switch_188_io_sel1 = r_mux_bus_ff_377; // @[Benes.scala 124:26]
  assign imm_switch_189_io_in0 = w_internal_420; // @[Benes.scala 109:25]
  assign imm_switch_189_io_in1 = w_internal_401; // @[Benes.scala 114:29]
  assign imm_switch_189_io_sel0 = r_mux_bus_ff_378; // @[Benes.scala 123:26]
  assign imm_switch_189_io_sel1 = r_mux_bus_ff_379; // @[Benes.scala 124:26]
  assign imm_switch_190_io_in0 = w_internal_422; // @[Benes.scala 109:25]
  assign imm_switch_190_io_in1 = w_internal_463; // @[Benes.scala 112:29]
  assign imm_switch_190_io_sel0 = r_mux_bus_ff_380; // @[Benes.scala 123:26]
  assign imm_switch_190_io_sel1 = r_mux_bus_ff_381; // @[Benes.scala 124:26]
  assign imm_switch_191_io_in0 = w_internal_424; // @[Benes.scala 109:25]
  assign imm_switch_191_io_in1 = w_internal_345; // @[Benes.scala 114:29]
  assign imm_switch_191_io_sel0 = r_mux_bus_ff_382; // @[Benes.scala 123:26]
  assign imm_switch_191_io_sel1 = r_mux_bus_ff_383; // @[Benes.scala 124:26]
  assign imm_switch_192_io_in0 = w_internal_426; // @[Benes.scala 109:25]
  assign imm_switch_192_io_in1 = w_internal_587; // @[Benes.scala 112:29]
  assign imm_switch_192_io_sel0 = r_mux_bus_ff_384; // @[Benes.scala 123:26]
  assign imm_switch_192_io_sel1 = r_mux_bus_ff_385; // @[Benes.scala 124:26]
  assign imm_switch_193_io_in0 = w_internal_428; // @[Benes.scala 109:25]
  assign imm_switch_193_io_in1 = w_internal_109; // @[Benes.scala 114:29]
  assign imm_switch_193_io_sel0 = r_mux_bus_ff_386; // @[Benes.scala 123:26]
  assign imm_switch_193_io_sel1 = r_mux_bus_ff_387; // @[Benes.scala 124:26]
  assign imm_switch_194_io_in0 = w_internal_430; // @[Benes.scala 109:25]
  assign imm_switch_194_io_in1 = w_internal_111; // @[Benes.scala 120:29]
  assign imm_switch_194_io_sel0 = r_mux_bus_ff_388; // @[Benes.scala 123:26]
  assign imm_switch_194_io_sel1 = r_mux_bus_ff_389; // @[Benes.scala 124:26]
  assign imm_switch_195_io_in0 = w_internal_432; // @[Benes.scala 109:25]
  assign imm_switch_195_io_in1 = w_internal_593; // @[Benes.scala 118:29]
  assign imm_switch_195_io_sel0 = r_mux_bus_ff_390; // @[Benes.scala 123:26]
  assign imm_switch_195_io_sel1 = r_mux_bus_ff_391; // @[Benes.scala 124:26]
  assign imm_switch_196_io_in0 = w_internal_434; // @[Benes.scala 109:25]
  assign imm_switch_196_io_in1 = w_internal_355; // @[Benes.scala 120:29]
  assign imm_switch_196_io_sel0 = r_mux_bus_ff_392; // @[Benes.scala 123:26]
  assign imm_switch_196_io_sel1 = r_mux_bus_ff_393; // @[Benes.scala 124:26]
  assign imm_switch_197_io_in0 = w_internal_436; // @[Benes.scala 109:25]
  assign imm_switch_197_io_in1 = w_internal_477; // @[Benes.scala 118:29]
  assign imm_switch_197_io_sel0 = r_mux_bus_ff_394; // @[Benes.scala 123:26]
  assign imm_switch_197_io_sel1 = r_mux_bus_ff_395; // @[Benes.scala 124:26]
  assign imm_switch_198_io_in0 = w_internal_440; // @[Benes.scala 109:25]
  assign imm_switch_198_io_in1 = w_internal_461; // @[Benes.scala 112:29]
  assign imm_switch_198_io_sel0 = r_mux_bus_ff_396; // @[Benes.scala 123:26]
  assign imm_switch_198_io_sel1 = r_mux_bus_ff_397; // @[Benes.scala 124:26]
  assign imm_switch_199_io_in0 = w_internal_442; // @[Benes.scala 109:25]
  assign imm_switch_199_io_in1 = w_internal_403; // @[Benes.scala 114:29]
  assign imm_switch_199_io_sel0 = r_mux_bus_ff_398; // @[Benes.scala 123:26]
  assign imm_switch_199_io_sel1 = r_mux_bus_ff_399; // @[Benes.scala 124:26]
  assign imm_switch_200_io_in0 = w_internal_444; // @[Benes.scala 109:25]
  assign imm_switch_200_io_in1 = w_internal_365; // @[Benes.scala 114:29]
  assign imm_switch_200_io_sel0 = r_mux_bus_ff_400; // @[Benes.scala 123:26]
  assign imm_switch_200_io_sel1 = r_mux_bus_ff_401; // @[Benes.scala 124:26]
  assign imm_switch_201_io_in0 = w_internal_446; // @[Benes.scala 109:25]
  assign imm_switch_201_io_in1 = w_internal_607; // @[Benes.scala 112:29]
  assign imm_switch_201_io_sel0 = r_mux_bus_ff_402; // @[Benes.scala 123:26]
  assign imm_switch_201_io_sel1 = r_mux_bus_ff_403; // @[Benes.scala 124:26]
  assign imm_switch_202_io_in0 = w_internal_448; // @[Benes.scala 109:25]
  assign imm_switch_202_io_in1 = w_internal_129; // @[Benes.scala 114:29]
  assign imm_switch_202_io_sel0 = r_mux_bus_ff_404; // @[Benes.scala 123:26]
  assign imm_switch_202_io_sel1 = r_mux_bus_ff_405; // @[Benes.scala 124:26]
  assign imm_switch_203_io_in0 = w_internal_450; // @[Benes.scala 109:25]
  assign imm_switch_203_io_in1 = w_internal_131; // @[Benes.scala 120:29]
  assign imm_switch_203_io_sel0 = r_mux_bus_ff_406; // @[Benes.scala 123:26]
  assign imm_switch_203_io_sel1 = r_mux_bus_ff_407; // @[Benes.scala 124:26]
  assign imm_switch_204_io_in0 = w_internal_452; // @[Benes.scala 109:25]
  assign imm_switch_204_io_in1 = w_internal_613; // @[Benes.scala 118:29]
  assign imm_switch_204_io_sel0 = r_mux_bus_ff_408; // @[Benes.scala 123:26]
  assign imm_switch_204_io_sel1 = r_mux_bus_ff_409; // @[Benes.scala 124:26]
  assign imm_switch_205_io_in0 = w_internal_454; // @[Benes.scala 109:25]
  assign imm_switch_205_io_in1 = w_internal_375; // @[Benes.scala 120:29]
  assign imm_switch_205_io_sel0 = r_mux_bus_ff_410; // @[Benes.scala 123:26]
  assign imm_switch_205_io_sel1 = r_mux_bus_ff_411; // @[Benes.scala 124:26]
  assign imm_switch_206_io_in0 = w_internal_456; // @[Benes.scala 109:25]
  assign imm_switch_206_io_in1 = w_internal_417; // @[Benes.scala 120:29]
  assign imm_switch_206_io_sel0 = r_mux_bus_ff_412; // @[Benes.scala 123:26]
  assign imm_switch_206_io_sel1 = r_mux_bus_ff_413; // @[Benes.scala 124:26]
  assign imm_switch_207_io_in0 = w_internal_460; // @[Benes.scala 109:25]
  assign imm_switch_207_io_in1 = w_internal_441; // @[Benes.scala 114:29]
  assign imm_switch_207_io_sel0 = r_mux_bus_ff_414; // @[Benes.scala 123:26]
  assign imm_switch_207_io_sel1 = r_mux_bus_ff_415; // @[Benes.scala 124:26]
  assign imm_switch_208_io_in0 = w_internal_462; // @[Benes.scala 109:25]
  assign imm_switch_208_io_in1 = w_internal_423; // @[Benes.scala 114:29]
  assign imm_switch_208_io_sel0 = r_mux_bus_ff_416; // @[Benes.scala 123:26]
  assign imm_switch_208_io_sel1 = r_mux_bus_ff_417; // @[Benes.scala 124:26]
  assign imm_switch_209_io_in0 = w_internal_464; // @[Benes.scala 109:25]
  assign imm_switch_209_io_in1 = w_internal_385; // @[Benes.scala 114:29]
  assign imm_switch_209_io_sel0 = r_mux_bus_ff_418; // @[Benes.scala 123:26]
  assign imm_switch_209_io_sel1 = r_mux_bus_ff_419; // @[Benes.scala 124:26]
  assign imm_switch_210_io_in0 = w_internal_466; // @[Benes.scala 109:25]
  assign imm_switch_210_io_in1 = w_internal_627; // @[Benes.scala 112:29]
  assign imm_switch_210_io_sel0 = r_mux_bus_ff_420; // @[Benes.scala 123:26]
  assign imm_switch_210_io_sel1 = r_mux_bus_ff_421; // @[Benes.scala 124:26]
  assign imm_switch_211_io_in0 = w_internal_468; // @[Benes.scala 109:25]
  assign imm_switch_211_io_in1 = w_internal_149; // @[Benes.scala 114:29]
  assign imm_switch_211_io_sel0 = r_mux_bus_ff_422; // @[Benes.scala 123:26]
  assign imm_switch_211_io_sel1 = r_mux_bus_ff_423; // @[Benes.scala 124:26]
  assign imm_switch_212_io_in0 = w_internal_470; // @[Benes.scala 109:25]
  assign imm_switch_212_io_in1 = w_internal_151; // @[Benes.scala 120:29]
  assign imm_switch_212_io_sel0 = r_mux_bus_ff_424; // @[Benes.scala 123:26]
  assign imm_switch_212_io_sel1 = r_mux_bus_ff_425; // @[Benes.scala 124:26]
  assign imm_switch_213_io_in0 = w_internal_472; // @[Benes.scala 109:25]
  assign imm_switch_213_io_in1 = w_internal_633; // @[Benes.scala 118:29]
  assign imm_switch_213_io_sel0 = r_mux_bus_ff_426; // @[Benes.scala 123:26]
  assign imm_switch_213_io_sel1 = r_mux_bus_ff_427; // @[Benes.scala 124:26]
  assign imm_switch_214_io_in0 = w_internal_474; // @[Benes.scala 109:25]
  assign imm_switch_214_io_in1 = w_internal_395; // @[Benes.scala 120:29]
  assign imm_switch_214_io_sel0 = r_mux_bus_ff_428; // @[Benes.scala 123:26]
  assign imm_switch_214_io_sel1 = r_mux_bus_ff_429; // @[Benes.scala 124:26]
  assign imm_switch_215_io_in0 = w_internal_476; // @[Benes.scala 109:25]
  assign imm_switch_215_io_in1 = w_internal_437; // @[Benes.scala 120:29]
  assign imm_switch_215_io_sel0 = r_mux_bus_ff_430; // @[Benes.scala 123:26]
  assign imm_switch_215_io_sel1 = r_mux_bus_ff_431; // @[Benes.scala 124:26]
  assign imm_switch_216_io_in0 = w_internal_480; // @[Benes.scala 109:25]
  assign imm_switch_216_io_in1 = w_internal_501; // @[Benes.scala 112:29]
  assign imm_switch_216_io_sel0 = r_mux_bus_ff_432; // @[Benes.scala 123:26]
  assign imm_switch_216_io_sel1 = r_mux_bus_ff_433; // @[Benes.scala 124:26]
  assign imm_switch_217_io_in0 = w_internal_482; // @[Benes.scala 109:25]
  assign imm_switch_217_io_in1 = w_internal_523; // @[Benes.scala 112:29]
  assign imm_switch_217_io_sel0 = r_mux_bus_ff_434; // @[Benes.scala 123:26]
  assign imm_switch_217_io_sel1 = r_mux_bus_ff_435; // @[Benes.scala 124:26]
  assign imm_switch_218_io_in0 = w_internal_484; // @[Benes.scala 109:25]
  assign imm_switch_218_io_in1 = w_internal_565; // @[Benes.scala 112:29]
  assign imm_switch_218_io_sel0 = r_mux_bus_ff_436; // @[Benes.scala 123:26]
  assign imm_switch_218_io_sel1 = r_mux_bus_ff_437; // @[Benes.scala 124:26]
  assign imm_switch_219_io_in0 = w_internal_486; // @[Benes.scala 109:25]
  assign imm_switch_219_io_in1 = w_internal_327; // @[Benes.scala 114:29]
  assign imm_switch_219_io_sel0 = r_mux_bus_ff_438; // @[Benes.scala 123:26]
  assign imm_switch_219_io_sel1 = r_mux_bus_ff_439; // @[Benes.scala 124:26]
  assign imm_switch_220_io_in0 = w_internal_488; // @[Benes.scala 109:25]
  assign imm_switch_220_io_in1 = w_internal_169; // @[Benes.scala 114:29]
  assign imm_switch_220_io_sel0 = r_mux_bus_ff_440; // @[Benes.scala 123:26]
  assign imm_switch_220_io_sel1 = r_mux_bus_ff_441; // @[Benes.scala 124:26]
  assign imm_switch_221_io_in0 = w_internal_490; // @[Benes.scala 109:25]
  assign imm_switch_221_io_in1 = w_internal_171; // @[Benes.scala 120:29]
  assign imm_switch_221_io_sel0 = r_mux_bus_ff_442; // @[Benes.scala 123:26]
  assign imm_switch_221_io_sel1 = r_mux_bus_ff_443; // @[Benes.scala 124:26]
  assign imm_switch_222_io_in0 = w_internal_492; // @[Benes.scala 109:25]
  assign imm_switch_222_io_in1 = w_internal_333; // @[Benes.scala 120:29]
  assign imm_switch_222_io_sel0 = r_mux_bus_ff_444; // @[Benes.scala 123:26]
  assign imm_switch_222_io_sel1 = r_mux_bus_ff_445; // @[Benes.scala 124:26]
  assign imm_switch_223_io_in0 = w_internal_494; // @[Benes.scala 109:25]
  assign imm_switch_223_io_in1 = w_internal_575; // @[Benes.scala 118:29]
  assign imm_switch_223_io_sel0 = r_mux_bus_ff_446; // @[Benes.scala 123:26]
  assign imm_switch_223_io_sel1 = r_mux_bus_ff_447; // @[Benes.scala 124:26]
  assign imm_switch_224_io_in0 = w_internal_496; // @[Benes.scala 109:25]
  assign imm_switch_224_io_in1 = w_internal_537; // @[Benes.scala 118:29]
  assign imm_switch_224_io_sel0 = r_mux_bus_ff_448; // @[Benes.scala 123:26]
  assign imm_switch_224_io_sel1 = r_mux_bus_ff_449; // @[Benes.scala 124:26]
  assign imm_switch_225_io_in0 = w_internal_500; // @[Benes.scala 109:25]
  assign imm_switch_225_io_in1 = w_internal_481; // @[Benes.scala 114:29]
  assign imm_switch_225_io_sel0 = r_mux_bus_ff_450; // @[Benes.scala 123:26]
  assign imm_switch_225_io_sel1 = r_mux_bus_ff_451; // @[Benes.scala 124:26]
  assign imm_switch_226_io_in0 = w_internal_502; // @[Benes.scala 109:25]
  assign imm_switch_226_io_in1 = w_internal_543; // @[Benes.scala 112:29]
  assign imm_switch_226_io_sel0 = r_mux_bus_ff_452; // @[Benes.scala 123:26]
  assign imm_switch_226_io_sel1 = r_mux_bus_ff_453; // @[Benes.scala 124:26]
  assign imm_switch_227_io_in0 = w_internal_504; // @[Benes.scala 109:25]
  assign imm_switch_227_io_in1 = w_internal_585; // @[Benes.scala 112:29]
  assign imm_switch_227_io_sel0 = r_mux_bus_ff_454; // @[Benes.scala 123:26]
  assign imm_switch_227_io_sel1 = r_mux_bus_ff_455; // @[Benes.scala 124:26]
  assign imm_switch_228_io_in0 = w_internal_506; // @[Benes.scala 109:25]
  assign imm_switch_228_io_in1 = w_internal_347; // @[Benes.scala 114:29]
  assign imm_switch_228_io_sel0 = r_mux_bus_ff_456; // @[Benes.scala 123:26]
  assign imm_switch_228_io_sel1 = r_mux_bus_ff_457; // @[Benes.scala 124:26]
  assign imm_switch_229_io_in0 = w_internal_508; // @[Benes.scala 109:25]
  assign imm_switch_229_io_in1 = w_internal_189; // @[Benes.scala 114:29]
  assign imm_switch_229_io_sel0 = r_mux_bus_ff_458; // @[Benes.scala 123:26]
  assign imm_switch_229_io_sel1 = r_mux_bus_ff_459; // @[Benes.scala 124:26]
  assign imm_switch_230_io_in0 = w_internal_510; // @[Benes.scala 109:25]
  assign imm_switch_230_io_in1 = w_internal_191; // @[Benes.scala 120:29]
  assign imm_switch_230_io_sel0 = r_mux_bus_ff_460; // @[Benes.scala 123:26]
  assign imm_switch_230_io_sel1 = r_mux_bus_ff_461; // @[Benes.scala 124:26]
  assign imm_switch_231_io_in0 = w_internal_512; // @[Benes.scala 109:25]
  assign imm_switch_231_io_in1 = w_internal_353; // @[Benes.scala 120:29]
  assign imm_switch_231_io_sel0 = r_mux_bus_ff_462; // @[Benes.scala 123:26]
  assign imm_switch_231_io_sel1 = r_mux_bus_ff_463; // @[Benes.scala 124:26]
  assign imm_switch_232_io_in0 = w_internal_514; // @[Benes.scala 109:25]
  assign imm_switch_232_io_in1 = w_internal_595; // @[Benes.scala 118:29]
  assign imm_switch_232_io_sel0 = r_mux_bus_ff_464; // @[Benes.scala 123:26]
  assign imm_switch_232_io_sel1 = r_mux_bus_ff_465; // @[Benes.scala 124:26]
  assign imm_switch_233_io_in0 = w_internal_516; // @[Benes.scala 109:25]
  assign imm_switch_233_io_in1 = w_internal_557; // @[Benes.scala 118:29]
  assign imm_switch_233_io_sel0 = r_mux_bus_ff_466; // @[Benes.scala 123:26]
  assign imm_switch_233_io_sel1 = r_mux_bus_ff_467; // @[Benes.scala 124:26]
  assign imm_switch_234_io_in0 = w_internal_520; // @[Benes.scala 109:25]
  assign imm_switch_234_io_in1 = w_internal_541; // @[Benes.scala 112:29]
  assign imm_switch_234_io_sel0 = r_mux_bus_ff_468; // @[Benes.scala 123:26]
  assign imm_switch_234_io_sel1 = r_mux_bus_ff_469; // @[Benes.scala 124:26]
  assign imm_switch_235_io_in0 = w_internal_522; // @[Benes.scala 109:25]
  assign imm_switch_235_io_in1 = w_internal_483; // @[Benes.scala 114:29]
  assign imm_switch_235_io_sel0 = r_mux_bus_ff_470; // @[Benes.scala 123:26]
  assign imm_switch_235_io_sel1 = r_mux_bus_ff_471; // @[Benes.scala 124:26]
  assign imm_switch_236_io_in0 = w_internal_524; // @[Benes.scala 109:25]
  assign imm_switch_236_io_in1 = w_internal_605; // @[Benes.scala 112:29]
  assign imm_switch_236_io_sel0 = r_mux_bus_ff_472; // @[Benes.scala 123:26]
  assign imm_switch_236_io_sel1 = r_mux_bus_ff_473; // @[Benes.scala 124:26]
  assign imm_switch_237_io_in0 = w_internal_526; // @[Benes.scala 109:25]
  assign imm_switch_237_io_in1 = w_internal_367; // @[Benes.scala 114:29]
  assign imm_switch_237_io_sel0 = r_mux_bus_ff_474; // @[Benes.scala 123:26]
  assign imm_switch_237_io_sel1 = r_mux_bus_ff_475; // @[Benes.scala 124:26]
  assign imm_switch_238_io_in0 = w_internal_528; // @[Benes.scala 109:25]
  assign imm_switch_238_io_in1 = w_internal_209; // @[Benes.scala 114:29]
  assign imm_switch_238_io_sel0 = r_mux_bus_ff_476; // @[Benes.scala 123:26]
  assign imm_switch_238_io_sel1 = r_mux_bus_ff_477; // @[Benes.scala 124:26]
  assign imm_switch_239_io_in0 = w_internal_530; // @[Benes.scala 109:25]
  assign imm_switch_239_io_in1 = w_internal_211; // @[Benes.scala 120:29]
  assign imm_switch_239_io_sel0 = r_mux_bus_ff_478; // @[Benes.scala 123:26]
  assign imm_switch_239_io_sel1 = r_mux_bus_ff_479; // @[Benes.scala 124:26]
  assign imm_switch_240_io_in0 = w_internal_532; // @[Benes.scala 109:25]
  assign imm_switch_240_io_in1 = w_internal_373; // @[Benes.scala 120:29]
  assign imm_switch_240_io_sel0 = r_mux_bus_ff_480; // @[Benes.scala 123:26]
  assign imm_switch_240_io_sel1 = r_mux_bus_ff_481; // @[Benes.scala 124:26]
  assign imm_switch_241_io_in0 = w_internal_534; // @[Benes.scala 109:25]
  assign imm_switch_241_io_in1 = w_internal_615; // @[Benes.scala 118:29]
  assign imm_switch_241_io_sel0 = r_mux_bus_ff_482; // @[Benes.scala 123:26]
  assign imm_switch_241_io_sel1 = r_mux_bus_ff_483; // @[Benes.scala 124:26]
  assign imm_switch_242_io_in0 = w_internal_536; // @[Benes.scala 109:25]
  assign imm_switch_242_io_in1 = w_internal_497; // @[Benes.scala 120:29]
  assign imm_switch_242_io_sel0 = r_mux_bus_ff_484; // @[Benes.scala 123:26]
  assign imm_switch_242_io_sel1 = r_mux_bus_ff_485; // @[Benes.scala 124:26]
  assign imm_switch_243_io_in0 = w_internal_540; // @[Benes.scala 109:25]
  assign imm_switch_243_io_in1 = w_internal_521; // @[Benes.scala 114:29]
  assign imm_switch_243_io_sel0 = r_mux_bus_ff_486; // @[Benes.scala 123:26]
  assign imm_switch_243_io_sel1 = r_mux_bus_ff_487; // @[Benes.scala 124:26]
  assign imm_switch_244_io_in0 = w_internal_542; // @[Benes.scala 109:25]
  assign imm_switch_244_io_in1 = w_internal_503; // @[Benes.scala 114:29]
  assign imm_switch_244_io_sel0 = r_mux_bus_ff_488; // @[Benes.scala 123:26]
  assign imm_switch_244_io_sel1 = r_mux_bus_ff_489; // @[Benes.scala 124:26]
  assign imm_switch_245_io_in0 = w_internal_544; // @[Benes.scala 109:25]
  assign imm_switch_245_io_in1 = w_internal_625; // @[Benes.scala 112:29]
  assign imm_switch_245_io_sel0 = r_mux_bus_ff_490; // @[Benes.scala 123:26]
  assign imm_switch_245_io_sel1 = r_mux_bus_ff_491; // @[Benes.scala 124:26]
  assign imm_switch_246_io_in0 = w_internal_546; // @[Benes.scala 109:25]
  assign imm_switch_246_io_in1 = w_internal_387; // @[Benes.scala 114:29]
  assign imm_switch_246_io_sel0 = r_mux_bus_ff_492; // @[Benes.scala 123:26]
  assign imm_switch_246_io_sel1 = r_mux_bus_ff_493; // @[Benes.scala 124:26]
  assign imm_switch_247_io_in0 = w_internal_548; // @[Benes.scala 109:25]
  assign imm_switch_247_io_in1 = w_internal_229; // @[Benes.scala 114:29]
  assign imm_switch_247_io_sel0 = r_mux_bus_ff_494; // @[Benes.scala 123:26]
  assign imm_switch_247_io_sel1 = r_mux_bus_ff_495; // @[Benes.scala 124:26]
  assign imm_switch_248_io_in0 = w_internal_550; // @[Benes.scala 109:25]
  assign imm_switch_248_io_in1 = w_internal_231; // @[Benes.scala 120:29]
  assign imm_switch_248_io_sel0 = r_mux_bus_ff_496; // @[Benes.scala 123:26]
  assign imm_switch_248_io_sel1 = r_mux_bus_ff_497; // @[Benes.scala 124:26]
  assign imm_switch_249_io_in0 = w_internal_552; // @[Benes.scala 109:25]
  assign imm_switch_249_io_in1 = w_internal_393; // @[Benes.scala 120:29]
  assign imm_switch_249_io_sel0 = r_mux_bus_ff_498; // @[Benes.scala 123:26]
  assign imm_switch_249_io_sel1 = r_mux_bus_ff_499; // @[Benes.scala 124:26]
  assign imm_switch_250_io_in0 = w_internal_554; // @[Benes.scala 109:25]
  assign imm_switch_250_io_in1 = w_internal_635; // @[Benes.scala 118:29]
  assign imm_switch_250_io_sel0 = r_mux_bus_ff_500; // @[Benes.scala 123:26]
  assign imm_switch_250_io_sel1 = r_mux_bus_ff_501; // @[Benes.scala 124:26]
  assign imm_switch_251_io_in0 = w_internal_556; // @[Benes.scala 109:25]
  assign imm_switch_251_io_in1 = w_internal_517; // @[Benes.scala 120:29]
  assign imm_switch_251_io_sel0 = r_mux_bus_ff_502; // @[Benes.scala 123:26]
  assign imm_switch_251_io_sel1 = r_mux_bus_ff_503; // @[Benes.scala 124:26]
  assign imm_switch_252_io_in0 = w_internal_560; // @[Benes.scala 109:25]
  assign imm_switch_252_io_in1 = w_internal_581; // @[Benes.scala 112:29]
  assign imm_switch_252_io_sel0 = r_mux_bus_ff_504; // @[Benes.scala 123:26]
  assign imm_switch_252_io_sel1 = r_mux_bus_ff_505; // @[Benes.scala 124:26]
  assign imm_switch_253_io_in0 = w_internal_562; // @[Benes.scala 109:25]
  assign imm_switch_253_io_in1 = w_internal_603; // @[Benes.scala 112:29]
  assign imm_switch_253_io_sel0 = r_mux_bus_ff_506; // @[Benes.scala 123:26]
  assign imm_switch_253_io_sel1 = r_mux_bus_ff_507; // @[Benes.scala 124:26]
  assign imm_switch_254_io_in0 = w_internal_564; // @[Benes.scala 109:25]
  assign imm_switch_254_io_in1 = w_internal_485; // @[Benes.scala 114:29]
  assign imm_switch_254_io_sel0 = r_mux_bus_ff_508; // @[Benes.scala 123:26]
  assign imm_switch_254_io_sel1 = r_mux_bus_ff_509; // @[Benes.scala 124:26]
  assign imm_switch_255_io_in0 = w_internal_566; // @[Benes.scala 109:25]
  assign imm_switch_255_io_in1 = w_internal_407; // @[Benes.scala 114:29]
  assign imm_switch_255_io_sel0 = r_mux_bus_ff_510; // @[Benes.scala 123:26]
  assign imm_switch_255_io_sel1 = r_mux_bus_ff_511; // @[Benes.scala 124:26]
  assign imm_switch_256_io_in0 = w_internal_568; // @[Benes.scala 109:25]
  assign imm_switch_256_io_in1 = w_internal_249; // @[Benes.scala 114:29]
  assign imm_switch_256_io_sel0 = r_mux_bus_ff_512; // @[Benes.scala 123:26]
  assign imm_switch_256_io_sel1 = r_mux_bus_ff_513; // @[Benes.scala 124:26]
  assign imm_switch_257_io_in0 = w_internal_570; // @[Benes.scala 109:25]
  assign imm_switch_257_io_in1 = w_internal_251; // @[Benes.scala 120:29]
  assign imm_switch_257_io_sel0 = r_mux_bus_ff_514; // @[Benes.scala 123:26]
  assign imm_switch_257_io_sel1 = r_mux_bus_ff_515; // @[Benes.scala 124:26]
  assign imm_switch_258_io_in0 = w_internal_572; // @[Benes.scala 109:25]
  assign imm_switch_258_io_in1 = w_internal_413; // @[Benes.scala 120:29]
  assign imm_switch_258_io_sel0 = r_mux_bus_ff_516; // @[Benes.scala 123:26]
  assign imm_switch_258_io_sel1 = r_mux_bus_ff_517; // @[Benes.scala 124:26]
  assign imm_switch_259_io_in0 = w_internal_574; // @[Benes.scala 109:25]
  assign imm_switch_259_io_in1 = w_internal_495; // @[Benes.scala 120:29]
  assign imm_switch_259_io_sel0 = r_mux_bus_ff_518; // @[Benes.scala 123:26]
  assign imm_switch_259_io_sel1 = r_mux_bus_ff_519; // @[Benes.scala 124:26]
  assign imm_switch_260_io_in0 = w_internal_576; // @[Benes.scala 109:25]
  assign imm_switch_260_io_in1 = w_internal_617; // @[Benes.scala 118:29]
  assign imm_switch_260_io_sel0 = r_mux_bus_ff_520; // @[Benes.scala 123:26]
  assign imm_switch_260_io_sel1 = r_mux_bus_ff_521; // @[Benes.scala 124:26]
  assign imm_switch_261_io_in0 = w_internal_580; // @[Benes.scala 109:25]
  assign imm_switch_261_io_in1 = w_internal_561; // @[Benes.scala 114:29]
  assign imm_switch_261_io_sel0 = r_mux_bus_ff_522; // @[Benes.scala 123:26]
  assign imm_switch_261_io_sel1 = r_mux_bus_ff_523; // @[Benes.scala 124:26]
  assign imm_switch_262_io_in0 = w_internal_582; // @[Benes.scala 109:25]
  assign imm_switch_262_io_in1 = w_internal_623; // @[Benes.scala 112:29]
  assign imm_switch_262_io_sel0 = r_mux_bus_ff_524; // @[Benes.scala 123:26]
  assign imm_switch_262_io_sel1 = r_mux_bus_ff_525; // @[Benes.scala 124:26]
  assign imm_switch_263_io_in0 = w_internal_584; // @[Benes.scala 109:25]
  assign imm_switch_263_io_in1 = w_internal_505; // @[Benes.scala 114:29]
  assign imm_switch_263_io_sel0 = r_mux_bus_ff_526; // @[Benes.scala 123:26]
  assign imm_switch_263_io_sel1 = r_mux_bus_ff_527; // @[Benes.scala 124:26]
  assign imm_switch_264_io_in0 = w_internal_586; // @[Benes.scala 109:25]
  assign imm_switch_264_io_in1 = w_internal_427; // @[Benes.scala 114:29]
  assign imm_switch_264_io_sel0 = r_mux_bus_ff_528; // @[Benes.scala 123:26]
  assign imm_switch_264_io_sel1 = r_mux_bus_ff_529; // @[Benes.scala 124:26]
  assign imm_switch_265_io_in0 = w_internal_588; // @[Benes.scala 109:25]
  assign imm_switch_265_io_in1 = w_internal_269; // @[Benes.scala 114:29]
  assign imm_switch_265_io_sel0 = r_mux_bus_ff_530; // @[Benes.scala 123:26]
  assign imm_switch_265_io_sel1 = r_mux_bus_ff_531; // @[Benes.scala 124:26]
  assign imm_switch_266_io_in0 = w_internal_590; // @[Benes.scala 109:25]
  assign imm_switch_266_io_in1 = w_internal_271; // @[Benes.scala 120:29]
  assign imm_switch_266_io_sel0 = r_mux_bus_ff_532; // @[Benes.scala 123:26]
  assign imm_switch_266_io_sel1 = r_mux_bus_ff_533; // @[Benes.scala 124:26]
  assign imm_switch_267_io_in0 = w_internal_592; // @[Benes.scala 109:25]
  assign imm_switch_267_io_in1 = w_internal_433; // @[Benes.scala 120:29]
  assign imm_switch_267_io_sel0 = r_mux_bus_ff_534; // @[Benes.scala 123:26]
  assign imm_switch_267_io_sel1 = r_mux_bus_ff_535; // @[Benes.scala 124:26]
  assign imm_switch_268_io_in0 = w_internal_594; // @[Benes.scala 109:25]
  assign imm_switch_268_io_in1 = w_internal_515; // @[Benes.scala 120:29]
  assign imm_switch_268_io_sel0 = r_mux_bus_ff_536; // @[Benes.scala 123:26]
  assign imm_switch_268_io_sel1 = r_mux_bus_ff_537; // @[Benes.scala 124:26]
  assign imm_switch_269_io_in0 = w_internal_596; // @[Benes.scala 109:25]
  assign imm_switch_269_io_in1 = w_internal_637; // @[Benes.scala 118:29]
  assign imm_switch_269_io_sel0 = r_mux_bus_ff_538; // @[Benes.scala 123:26]
  assign imm_switch_269_io_sel1 = r_mux_bus_ff_539; // @[Benes.scala 124:26]
  assign imm_switch_270_io_in0 = w_internal_600; // @[Benes.scala 109:25]
  assign imm_switch_270_io_in1 = w_internal_621; // @[Benes.scala 112:29]
  assign imm_switch_270_io_sel0 = r_mux_bus_ff_540; // @[Benes.scala 123:26]
  assign imm_switch_270_io_sel1 = r_mux_bus_ff_541; // @[Benes.scala 124:26]
  assign imm_switch_271_io_in0 = w_internal_602; // @[Benes.scala 109:25]
  assign imm_switch_271_io_in1 = w_internal_563; // @[Benes.scala 114:29]
  assign imm_switch_271_io_sel0 = r_mux_bus_ff_542; // @[Benes.scala 123:26]
  assign imm_switch_271_io_sel1 = r_mux_bus_ff_543; // @[Benes.scala 124:26]
  assign imm_switch_272_io_in0 = w_internal_604; // @[Benes.scala 109:25]
  assign imm_switch_272_io_in1 = w_internal_525; // @[Benes.scala 114:29]
  assign imm_switch_272_io_sel0 = r_mux_bus_ff_544; // @[Benes.scala 123:26]
  assign imm_switch_272_io_sel1 = r_mux_bus_ff_545; // @[Benes.scala 124:26]
  assign imm_switch_273_io_in0 = w_internal_606; // @[Benes.scala 109:25]
  assign imm_switch_273_io_in1 = w_internal_447; // @[Benes.scala 114:29]
  assign imm_switch_273_io_sel0 = r_mux_bus_ff_546; // @[Benes.scala 123:26]
  assign imm_switch_273_io_sel1 = r_mux_bus_ff_547; // @[Benes.scala 124:26]
  assign imm_switch_274_io_in0 = w_internal_608; // @[Benes.scala 109:25]
  assign imm_switch_274_io_in1 = w_internal_289; // @[Benes.scala 114:29]
  assign imm_switch_274_io_sel0 = r_mux_bus_ff_548; // @[Benes.scala 123:26]
  assign imm_switch_274_io_sel1 = r_mux_bus_ff_549; // @[Benes.scala 124:26]
  assign imm_switch_275_io_in0 = w_internal_610; // @[Benes.scala 109:25]
  assign imm_switch_275_io_in1 = w_internal_291; // @[Benes.scala 120:29]
  assign imm_switch_275_io_sel0 = r_mux_bus_ff_550; // @[Benes.scala 123:26]
  assign imm_switch_275_io_sel1 = r_mux_bus_ff_551; // @[Benes.scala 124:26]
  assign imm_switch_276_io_in0 = w_internal_612; // @[Benes.scala 109:25]
  assign imm_switch_276_io_in1 = w_internal_453; // @[Benes.scala 120:29]
  assign imm_switch_276_io_sel0 = r_mux_bus_ff_552; // @[Benes.scala 123:26]
  assign imm_switch_276_io_sel1 = r_mux_bus_ff_553; // @[Benes.scala 124:26]
  assign imm_switch_277_io_in0 = w_internal_614; // @[Benes.scala 109:25]
  assign imm_switch_277_io_in1 = w_internal_535; // @[Benes.scala 120:29]
  assign imm_switch_277_io_sel0 = r_mux_bus_ff_554; // @[Benes.scala 123:26]
  assign imm_switch_277_io_sel1 = r_mux_bus_ff_555; // @[Benes.scala 124:26]
  assign imm_switch_278_io_in0 = w_internal_616; // @[Benes.scala 109:25]
  assign imm_switch_278_io_in1 = w_internal_577; // @[Benes.scala 120:29]
  assign imm_switch_278_io_sel0 = r_mux_bus_ff_556; // @[Benes.scala 123:26]
  assign imm_switch_278_io_sel1 = r_mux_bus_ff_557; // @[Benes.scala 124:26]
  assign imm_switch_279_io_in0 = w_internal_620; // @[Benes.scala 109:25]
  assign imm_switch_279_io_in1 = w_internal_601; // @[Benes.scala 114:29]
  assign imm_switch_279_io_sel0 = r_mux_bus_ff_558; // @[Benes.scala 123:26]
  assign imm_switch_279_io_sel1 = r_mux_bus_ff_559; // @[Benes.scala 124:26]
  assign imm_switch_280_io_in0 = w_internal_622; // @[Benes.scala 109:25]
  assign imm_switch_280_io_in1 = w_internal_583; // @[Benes.scala 114:29]
  assign imm_switch_280_io_sel0 = r_mux_bus_ff_560; // @[Benes.scala 123:26]
  assign imm_switch_280_io_sel1 = r_mux_bus_ff_561; // @[Benes.scala 124:26]
  assign imm_switch_281_io_in0 = w_internal_624; // @[Benes.scala 109:25]
  assign imm_switch_281_io_in1 = w_internal_545; // @[Benes.scala 114:29]
  assign imm_switch_281_io_sel0 = r_mux_bus_ff_562; // @[Benes.scala 123:26]
  assign imm_switch_281_io_sel1 = r_mux_bus_ff_563; // @[Benes.scala 124:26]
  assign imm_switch_282_io_in0 = w_internal_626; // @[Benes.scala 109:25]
  assign imm_switch_282_io_in1 = w_internal_467; // @[Benes.scala 114:29]
  assign imm_switch_282_io_sel0 = r_mux_bus_ff_564; // @[Benes.scala 123:26]
  assign imm_switch_282_io_sel1 = r_mux_bus_ff_565; // @[Benes.scala 124:26]
  assign imm_switch_283_io_in0 = w_internal_628; // @[Benes.scala 109:25]
  assign imm_switch_283_io_in1 = w_internal_309; // @[Benes.scala 114:29]
  assign imm_switch_283_io_sel0 = r_mux_bus_ff_566; // @[Benes.scala 123:26]
  assign imm_switch_283_io_sel1 = r_mux_bus_ff_567; // @[Benes.scala 124:26]
  assign imm_switch_284_io_in0 = w_internal_630; // @[Benes.scala 109:25]
  assign imm_switch_284_io_in1 = w_internal_311; // @[Benes.scala 120:29]
  assign imm_switch_284_io_sel0 = r_mux_bus_ff_568; // @[Benes.scala 123:26]
  assign imm_switch_284_io_sel1 = r_mux_bus_ff_569; // @[Benes.scala 124:26]
  assign imm_switch_285_io_in0 = w_internal_632; // @[Benes.scala 109:25]
  assign imm_switch_285_io_in1 = w_internal_473; // @[Benes.scala 120:29]
  assign imm_switch_285_io_sel0 = r_mux_bus_ff_570; // @[Benes.scala 123:26]
  assign imm_switch_285_io_sel1 = r_mux_bus_ff_571; // @[Benes.scala 124:26]
  assign imm_switch_286_io_in0 = w_internal_634; // @[Benes.scala 109:25]
  assign imm_switch_286_io_in1 = w_internal_555; // @[Benes.scala 120:29]
  assign imm_switch_286_io_sel0 = r_mux_bus_ff_572; // @[Benes.scala 123:26]
  assign imm_switch_286_io_sel1 = r_mux_bus_ff_573; // @[Benes.scala 124:26]
  assign imm_switch_287_io_in0 = w_internal_636; // @[Benes.scala 109:25]
  assign imm_switch_287_io_in1 = w_internal_597; // @[Benes.scala 120:29]
  assign imm_switch_287_io_sel0 = r_mux_bus_ff_574; // @[Benes.scala 123:26]
  assign imm_switch_287_io_sel1 = r_mux_bus_ff_575; // @[Benes.scala 124:26]
  always @(posedge clock) begin
    if (reset) begin // @[Benes.scala 76:32]
      r_data_bus_ff_0 <= 32'h0; // @[Benes.scala 76:32]
    end else if (reset) begin // @[Benes.scala 83:23]
      r_data_bus_ff_0 <= 32'h0;
    end else begin
      r_data_bus_ff_0 <= io_i_data_bus_0;
    end
    if (reset) begin // @[Benes.scala 76:32]
      r_data_bus_ff_1 <= 32'h0; // @[Benes.scala 76:32]
    end else if (reset) begin // @[Benes.scala 83:23]
      r_data_bus_ff_1 <= 32'h0;
    end else begin
      r_data_bus_ff_1 <= io_i_data_bus_1;
    end
    if (reset) begin // @[Benes.scala 76:32]
      r_data_bus_ff_2 <= 32'h0; // @[Benes.scala 76:32]
    end else if (reset) begin // @[Benes.scala 83:23]
      r_data_bus_ff_2 <= 32'h0;
    end else begin
      r_data_bus_ff_2 <= io_i_data_bus_2;
    end
    if (reset) begin // @[Benes.scala 76:32]
      r_data_bus_ff_3 <= 32'h0; // @[Benes.scala 76:32]
    end else if (reset) begin // @[Benes.scala 83:23]
      r_data_bus_ff_3 <= 32'h0;
    end else begin
      r_data_bus_ff_3 <= io_i_data_bus_3;
    end
    if (reset) begin // @[Benes.scala 76:32]
      r_data_bus_ff_4 <= 32'h0; // @[Benes.scala 76:32]
    end else if (reset) begin // @[Benes.scala 83:23]
      r_data_bus_ff_4 <= 32'h0;
    end else begin
      r_data_bus_ff_4 <= io_i_data_bus_4;
    end
    if (reset) begin // @[Benes.scala 76:32]
      r_data_bus_ff_5 <= 32'h0; // @[Benes.scala 76:32]
    end else if (reset) begin // @[Benes.scala 83:23]
      r_data_bus_ff_5 <= 32'h0;
    end else begin
      r_data_bus_ff_5 <= io_i_data_bus_5;
    end
    if (reset) begin // @[Benes.scala 76:32]
      r_data_bus_ff_6 <= 32'h0; // @[Benes.scala 76:32]
    end else if (reset) begin // @[Benes.scala 83:23]
      r_data_bus_ff_6 <= 32'h0;
    end else begin
      r_data_bus_ff_6 <= io_i_data_bus_6;
    end
    if (reset) begin // @[Benes.scala 76:32]
      r_data_bus_ff_7 <= 32'h0; // @[Benes.scala 76:32]
    end else if (reset) begin // @[Benes.scala 83:23]
      r_data_bus_ff_7 <= 32'h0;
    end else begin
      r_data_bus_ff_7 <= io_i_data_bus_7;
    end
    if (reset) begin // @[Benes.scala 76:32]
      r_data_bus_ff_8 <= 32'h0; // @[Benes.scala 76:32]
    end else if (reset) begin // @[Benes.scala 83:23]
      r_data_bus_ff_8 <= 32'h0;
    end else begin
      r_data_bus_ff_8 <= io_i_data_bus_8;
    end
    if (reset) begin // @[Benes.scala 76:32]
      r_data_bus_ff_9 <= 32'h0; // @[Benes.scala 76:32]
    end else if (reset) begin // @[Benes.scala 83:23]
      r_data_bus_ff_9 <= 32'h0;
    end else begin
      r_data_bus_ff_9 <= io_i_data_bus_9;
    end
    if (reset) begin // @[Benes.scala 76:32]
      r_data_bus_ff_10 <= 32'h0; // @[Benes.scala 76:32]
    end else if (reset) begin // @[Benes.scala 83:23]
      r_data_bus_ff_10 <= 32'h0;
    end else begin
      r_data_bus_ff_10 <= io_i_data_bus_10;
    end
    if (reset) begin // @[Benes.scala 76:32]
      r_data_bus_ff_11 <= 32'h0; // @[Benes.scala 76:32]
    end else if (reset) begin // @[Benes.scala 83:23]
      r_data_bus_ff_11 <= 32'h0;
    end else begin
      r_data_bus_ff_11 <= io_i_data_bus_11;
    end
    if (reset) begin // @[Benes.scala 76:32]
      r_data_bus_ff_12 <= 32'h0; // @[Benes.scala 76:32]
    end else if (reset) begin // @[Benes.scala 83:23]
      r_data_bus_ff_12 <= 32'h0;
    end else begin
      r_data_bus_ff_12 <= io_i_data_bus_12;
    end
    if (reset) begin // @[Benes.scala 76:32]
      r_data_bus_ff_13 <= 32'h0; // @[Benes.scala 76:32]
    end else if (reset) begin // @[Benes.scala 83:23]
      r_data_bus_ff_13 <= 32'h0;
    end else begin
      r_data_bus_ff_13 <= io_i_data_bus_13;
    end
    if (reset) begin // @[Benes.scala 76:32]
      r_data_bus_ff_14 <= 32'h0; // @[Benes.scala 76:32]
    end else if (reset) begin // @[Benes.scala 83:23]
      r_data_bus_ff_14 <= 32'h0;
    end else begin
      r_data_bus_ff_14 <= io_i_data_bus_14;
    end
    if (reset) begin // @[Benes.scala 76:32]
      r_data_bus_ff_15 <= 32'h0; // @[Benes.scala 76:32]
    end else if (reset) begin // @[Benes.scala 83:23]
      r_data_bus_ff_15 <= 32'h0;
    end else begin
      r_data_bus_ff_15 <= io_i_data_bus_15;
    end
    if (reset) begin // @[Benes.scala 76:32]
      r_data_bus_ff_16 <= 32'h0; // @[Benes.scala 76:32]
    end else if (reset) begin // @[Benes.scala 83:23]
      r_data_bus_ff_16 <= 32'h0;
    end else begin
      r_data_bus_ff_16 <= io_i_data_bus_16;
    end
    if (reset) begin // @[Benes.scala 76:32]
      r_data_bus_ff_17 <= 32'h0; // @[Benes.scala 76:32]
    end else if (reset) begin // @[Benes.scala 83:23]
      r_data_bus_ff_17 <= 32'h0;
    end else begin
      r_data_bus_ff_17 <= io_i_data_bus_17;
    end
    if (reset) begin // @[Benes.scala 76:32]
      r_data_bus_ff_18 <= 32'h0; // @[Benes.scala 76:32]
    end else if (reset) begin // @[Benes.scala 83:23]
      r_data_bus_ff_18 <= 32'h0;
    end else begin
      r_data_bus_ff_18 <= io_i_data_bus_18;
    end
    if (reset) begin // @[Benes.scala 76:32]
      r_data_bus_ff_19 <= 32'h0; // @[Benes.scala 76:32]
    end else if (reset) begin // @[Benes.scala 83:23]
      r_data_bus_ff_19 <= 32'h0;
    end else begin
      r_data_bus_ff_19 <= io_i_data_bus_19;
    end
    if (reset) begin // @[Benes.scala 76:32]
      r_data_bus_ff_20 <= 32'h0; // @[Benes.scala 76:32]
    end else if (reset) begin // @[Benes.scala 83:23]
      r_data_bus_ff_20 <= 32'h0;
    end else begin
      r_data_bus_ff_20 <= io_i_data_bus_20;
    end
    if (reset) begin // @[Benes.scala 76:32]
      r_data_bus_ff_21 <= 32'h0; // @[Benes.scala 76:32]
    end else if (reset) begin // @[Benes.scala 83:23]
      r_data_bus_ff_21 <= 32'h0;
    end else begin
      r_data_bus_ff_21 <= io_i_data_bus_21;
    end
    if (reset) begin // @[Benes.scala 76:32]
      r_data_bus_ff_22 <= 32'h0; // @[Benes.scala 76:32]
    end else if (reset) begin // @[Benes.scala 83:23]
      r_data_bus_ff_22 <= 32'h0;
    end else begin
      r_data_bus_ff_22 <= io_i_data_bus_22;
    end
    if (reset) begin // @[Benes.scala 76:32]
      r_data_bus_ff_23 <= 32'h0; // @[Benes.scala 76:32]
    end else if (reset) begin // @[Benes.scala 83:23]
      r_data_bus_ff_23 <= 32'h0;
    end else begin
      r_data_bus_ff_23 <= io_i_data_bus_23;
    end
    if (reset) begin // @[Benes.scala 76:32]
      r_data_bus_ff_24 <= 32'h0; // @[Benes.scala 76:32]
    end else if (reset) begin // @[Benes.scala 83:23]
      r_data_bus_ff_24 <= 32'h0;
    end else begin
      r_data_bus_ff_24 <= io_i_data_bus_24;
    end
    if (reset) begin // @[Benes.scala 76:32]
      r_data_bus_ff_25 <= 32'h0; // @[Benes.scala 76:32]
    end else if (reset) begin // @[Benes.scala 83:23]
      r_data_bus_ff_25 <= 32'h0;
    end else begin
      r_data_bus_ff_25 <= io_i_data_bus_25;
    end
    if (reset) begin // @[Benes.scala 76:32]
      r_data_bus_ff_26 <= 32'h0; // @[Benes.scala 76:32]
    end else if (reset) begin // @[Benes.scala 83:23]
      r_data_bus_ff_26 <= 32'h0;
    end else begin
      r_data_bus_ff_26 <= io_i_data_bus_26;
    end
    if (reset) begin // @[Benes.scala 76:32]
      r_data_bus_ff_27 <= 32'h0; // @[Benes.scala 76:32]
    end else if (reset) begin // @[Benes.scala 83:23]
      r_data_bus_ff_27 <= 32'h0;
    end else begin
      r_data_bus_ff_27 <= io_i_data_bus_27;
    end
    if (reset) begin // @[Benes.scala 76:32]
      r_data_bus_ff_28 <= 32'h0; // @[Benes.scala 76:32]
    end else if (reset) begin // @[Benes.scala 83:23]
      r_data_bus_ff_28 <= 32'h0;
    end else begin
      r_data_bus_ff_28 <= io_i_data_bus_28;
    end
    if (reset) begin // @[Benes.scala 76:32]
      r_data_bus_ff_29 <= 32'h0; // @[Benes.scala 76:32]
    end else if (reset) begin // @[Benes.scala 83:23]
      r_data_bus_ff_29 <= 32'h0;
    end else begin
      r_data_bus_ff_29 <= io_i_data_bus_29;
    end
    if (reset) begin // @[Benes.scala 76:32]
      r_data_bus_ff_30 <= 32'h0; // @[Benes.scala 76:32]
    end else if (reset) begin // @[Benes.scala 83:23]
      r_data_bus_ff_30 <= 32'h0;
    end else begin
      r_data_bus_ff_30 <= io_i_data_bus_30;
    end
    if (reset) begin // @[Benes.scala 76:32]
      r_data_bus_ff_31 <= 32'h0; // @[Benes.scala 76:32]
    end else if (reset) begin // @[Benes.scala 83:23]
      r_data_bus_ff_31 <= 32'h0;
    end else begin
      r_data_bus_ff_31 <= io_i_data_bus_31;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_0 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_0 <= 1'h0;
    end else begin
      r_mux_bus_ff_0 <= io_i_mux_bus_0;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_1 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_1 <= 1'h0;
    end else begin
      r_mux_bus_ff_1 <= io_i_mux_bus_1;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_2 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_2 <= 1'h0;
    end else begin
      r_mux_bus_ff_2 <= io_i_mux_bus_2;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_3 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_3 <= 1'h0;
    end else begin
      r_mux_bus_ff_3 <= io_i_mux_bus_3;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_4 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_4 <= 1'h0;
    end else begin
      r_mux_bus_ff_4 <= io_i_mux_bus_4;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_5 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_5 <= 1'h0;
    end else begin
      r_mux_bus_ff_5 <= io_i_mux_bus_5;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_6 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_6 <= 1'h0;
    end else begin
      r_mux_bus_ff_6 <= io_i_mux_bus_6;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_7 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_7 <= 1'h0;
    end else begin
      r_mux_bus_ff_7 <= io_i_mux_bus_7;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_8 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_8 <= 1'h0;
    end else begin
      r_mux_bus_ff_8 <= io_i_mux_bus_8;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_9 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_9 <= 1'h0;
    end else begin
      r_mux_bus_ff_9 <= io_i_mux_bus_9;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_10 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_10 <= 1'h0;
    end else begin
      r_mux_bus_ff_10 <= io_i_mux_bus_10;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_11 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_11 <= 1'h0;
    end else begin
      r_mux_bus_ff_11 <= io_i_mux_bus_11;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_12 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_12 <= 1'h0;
    end else begin
      r_mux_bus_ff_12 <= io_i_mux_bus_12;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_13 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_13 <= 1'h0;
    end else begin
      r_mux_bus_ff_13 <= io_i_mux_bus_13;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_14 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_14 <= 1'h0;
    end else begin
      r_mux_bus_ff_14 <= io_i_mux_bus_14;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_15 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_15 <= 1'h0;
    end else begin
      r_mux_bus_ff_15 <= io_i_mux_bus_15;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_16 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_16 <= 1'h0;
    end else begin
      r_mux_bus_ff_16 <= io_i_mux_bus_16;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_17 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_17 <= 1'h0;
    end else begin
      r_mux_bus_ff_17 <= io_i_mux_bus_17;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_18 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_18 <= 1'h0;
    end else begin
      r_mux_bus_ff_18 <= io_i_mux_bus_18;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_19 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_19 <= 1'h0;
    end else begin
      r_mux_bus_ff_19 <= io_i_mux_bus_19;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_20 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_20 <= 1'h0;
    end else begin
      r_mux_bus_ff_20 <= io_i_mux_bus_20;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_21 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_21 <= 1'h0;
    end else begin
      r_mux_bus_ff_21 <= io_i_mux_bus_21;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_22 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_22 <= 1'h0;
    end else begin
      r_mux_bus_ff_22 <= io_i_mux_bus_22;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_23 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_23 <= 1'h0;
    end else begin
      r_mux_bus_ff_23 <= io_i_mux_bus_23;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_24 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_24 <= 1'h0;
    end else begin
      r_mux_bus_ff_24 <= io_i_mux_bus_24;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_25 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_25 <= 1'h0;
    end else begin
      r_mux_bus_ff_25 <= io_i_mux_bus_25;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_26 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_26 <= 1'h0;
    end else begin
      r_mux_bus_ff_26 <= io_i_mux_bus_26;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_27 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_27 <= 1'h0;
    end else begin
      r_mux_bus_ff_27 <= io_i_mux_bus_27;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_28 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_28 <= 1'h0;
    end else begin
      r_mux_bus_ff_28 <= io_i_mux_bus_28;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_29 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_29 <= 1'h0;
    end else begin
      r_mux_bus_ff_29 <= io_i_mux_bus_29;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_30 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_30 <= 1'h0;
    end else begin
      r_mux_bus_ff_30 <= io_i_mux_bus_30;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_31 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_31 <= 1'h0;
    end else begin
      r_mux_bus_ff_31 <= io_i_mux_bus_31;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_32 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_32 <= 1'h0;
    end else begin
      r_mux_bus_ff_32 <= io_i_mux_bus_32;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_33 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_33 <= 1'h0;
    end else begin
      r_mux_bus_ff_33 <= io_i_mux_bus_33;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_34 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_34 <= 1'h0;
    end else begin
      r_mux_bus_ff_34 <= io_i_mux_bus_34;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_35 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_35 <= 1'h0;
    end else begin
      r_mux_bus_ff_35 <= io_i_mux_bus_35;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_36 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_36 <= 1'h0;
    end else begin
      r_mux_bus_ff_36 <= io_i_mux_bus_36;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_37 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_37 <= 1'h0;
    end else begin
      r_mux_bus_ff_37 <= io_i_mux_bus_37;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_38 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_38 <= 1'h0;
    end else begin
      r_mux_bus_ff_38 <= io_i_mux_bus_38;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_39 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_39 <= 1'h0;
    end else begin
      r_mux_bus_ff_39 <= io_i_mux_bus_39;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_40 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_40 <= 1'h0;
    end else begin
      r_mux_bus_ff_40 <= io_i_mux_bus_40;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_41 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_41 <= 1'h0;
    end else begin
      r_mux_bus_ff_41 <= io_i_mux_bus_41;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_42 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_42 <= 1'h0;
    end else begin
      r_mux_bus_ff_42 <= io_i_mux_bus_42;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_43 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_43 <= 1'h0;
    end else begin
      r_mux_bus_ff_43 <= io_i_mux_bus_43;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_44 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_44 <= 1'h0;
    end else begin
      r_mux_bus_ff_44 <= io_i_mux_bus_44;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_45 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_45 <= 1'h0;
    end else begin
      r_mux_bus_ff_45 <= io_i_mux_bus_45;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_46 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_46 <= 1'h0;
    end else begin
      r_mux_bus_ff_46 <= io_i_mux_bus_46;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_47 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_47 <= 1'h0;
    end else begin
      r_mux_bus_ff_47 <= io_i_mux_bus_47;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_48 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_48 <= 1'h0;
    end else begin
      r_mux_bus_ff_48 <= io_i_mux_bus_48;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_49 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_49 <= 1'h0;
    end else begin
      r_mux_bus_ff_49 <= io_i_mux_bus_49;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_50 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_50 <= 1'h0;
    end else begin
      r_mux_bus_ff_50 <= io_i_mux_bus_50;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_51 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_51 <= 1'h0;
    end else begin
      r_mux_bus_ff_51 <= io_i_mux_bus_51;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_52 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_52 <= 1'h0;
    end else begin
      r_mux_bus_ff_52 <= io_i_mux_bus_52;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_53 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_53 <= 1'h0;
    end else begin
      r_mux_bus_ff_53 <= io_i_mux_bus_53;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_54 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_54 <= 1'h0;
    end else begin
      r_mux_bus_ff_54 <= io_i_mux_bus_54;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_55 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_55 <= 1'h0;
    end else begin
      r_mux_bus_ff_55 <= io_i_mux_bus_55;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_56 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_56 <= 1'h0;
    end else begin
      r_mux_bus_ff_56 <= io_i_mux_bus_56;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_57 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_57 <= 1'h0;
    end else begin
      r_mux_bus_ff_57 <= io_i_mux_bus_57;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_58 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_58 <= 1'h0;
    end else begin
      r_mux_bus_ff_58 <= io_i_mux_bus_58;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_59 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_59 <= 1'h0;
    end else begin
      r_mux_bus_ff_59 <= io_i_mux_bus_59;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_60 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_60 <= 1'h0;
    end else begin
      r_mux_bus_ff_60 <= io_i_mux_bus_60;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_61 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_61 <= 1'h0;
    end else begin
      r_mux_bus_ff_61 <= io_i_mux_bus_61;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_62 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_62 <= 1'h0;
    end else begin
      r_mux_bus_ff_62 <= io_i_mux_bus_62;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_63 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_63 <= 1'h0;
    end else begin
      r_mux_bus_ff_63 <= io_i_mux_bus_63;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_64 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_64 <= 1'h0;
    end else begin
      r_mux_bus_ff_64 <= io_i_mux_bus_64;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_65 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_65 <= 1'h0;
    end else begin
      r_mux_bus_ff_65 <= io_i_mux_bus_65;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_66 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_66 <= 1'h0;
    end else begin
      r_mux_bus_ff_66 <= io_i_mux_bus_66;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_67 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_67 <= 1'h0;
    end else begin
      r_mux_bus_ff_67 <= io_i_mux_bus_67;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_68 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_68 <= 1'h0;
    end else begin
      r_mux_bus_ff_68 <= io_i_mux_bus_68;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_69 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_69 <= 1'h0;
    end else begin
      r_mux_bus_ff_69 <= io_i_mux_bus_69;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_70 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_70 <= 1'h0;
    end else begin
      r_mux_bus_ff_70 <= io_i_mux_bus_70;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_71 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_71 <= 1'h0;
    end else begin
      r_mux_bus_ff_71 <= io_i_mux_bus_71;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_72 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_72 <= 1'h0;
    end else begin
      r_mux_bus_ff_72 <= io_i_mux_bus_72;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_73 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_73 <= 1'h0;
    end else begin
      r_mux_bus_ff_73 <= io_i_mux_bus_73;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_74 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_74 <= 1'h0;
    end else begin
      r_mux_bus_ff_74 <= io_i_mux_bus_74;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_75 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_75 <= 1'h0;
    end else begin
      r_mux_bus_ff_75 <= io_i_mux_bus_75;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_76 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_76 <= 1'h0;
    end else begin
      r_mux_bus_ff_76 <= io_i_mux_bus_76;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_77 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_77 <= 1'h0;
    end else begin
      r_mux_bus_ff_77 <= io_i_mux_bus_77;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_78 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_78 <= 1'h0;
    end else begin
      r_mux_bus_ff_78 <= io_i_mux_bus_78;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_79 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_79 <= 1'h0;
    end else begin
      r_mux_bus_ff_79 <= io_i_mux_bus_79;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_80 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_80 <= 1'h0;
    end else begin
      r_mux_bus_ff_80 <= io_i_mux_bus_80;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_81 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_81 <= 1'h0;
    end else begin
      r_mux_bus_ff_81 <= io_i_mux_bus_81;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_82 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_82 <= 1'h0;
    end else begin
      r_mux_bus_ff_82 <= io_i_mux_bus_82;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_83 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_83 <= 1'h0;
    end else begin
      r_mux_bus_ff_83 <= io_i_mux_bus_83;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_84 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_84 <= 1'h0;
    end else begin
      r_mux_bus_ff_84 <= io_i_mux_bus_84;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_85 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_85 <= 1'h0;
    end else begin
      r_mux_bus_ff_85 <= io_i_mux_bus_85;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_86 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_86 <= 1'h0;
    end else begin
      r_mux_bus_ff_86 <= io_i_mux_bus_86;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_87 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_87 <= 1'h0;
    end else begin
      r_mux_bus_ff_87 <= io_i_mux_bus_87;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_88 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_88 <= 1'h0;
    end else begin
      r_mux_bus_ff_88 <= io_i_mux_bus_88;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_89 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_89 <= 1'h0;
    end else begin
      r_mux_bus_ff_89 <= io_i_mux_bus_89;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_90 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_90 <= 1'h0;
    end else begin
      r_mux_bus_ff_90 <= io_i_mux_bus_90;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_91 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_91 <= 1'h0;
    end else begin
      r_mux_bus_ff_91 <= io_i_mux_bus_91;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_92 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_92 <= 1'h0;
    end else begin
      r_mux_bus_ff_92 <= io_i_mux_bus_92;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_93 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_93 <= 1'h0;
    end else begin
      r_mux_bus_ff_93 <= io_i_mux_bus_93;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_94 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_94 <= 1'h0;
    end else begin
      r_mux_bus_ff_94 <= io_i_mux_bus_94;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_95 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_95 <= 1'h0;
    end else begin
      r_mux_bus_ff_95 <= io_i_mux_bus_95;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_96 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_96 <= 1'h0;
    end else begin
      r_mux_bus_ff_96 <= io_i_mux_bus_96;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_97 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_97 <= 1'h0;
    end else begin
      r_mux_bus_ff_97 <= io_i_mux_bus_97;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_98 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_98 <= 1'h0;
    end else begin
      r_mux_bus_ff_98 <= io_i_mux_bus_98;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_99 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_99 <= 1'h0;
    end else begin
      r_mux_bus_ff_99 <= io_i_mux_bus_99;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_100 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_100 <= 1'h0;
    end else begin
      r_mux_bus_ff_100 <= io_i_mux_bus_100;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_101 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_101 <= 1'h0;
    end else begin
      r_mux_bus_ff_101 <= io_i_mux_bus_101;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_102 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_102 <= 1'h0;
    end else begin
      r_mux_bus_ff_102 <= io_i_mux_bus_102;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_103 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_103 <= 1'h0;
    end else begin
      r_mux_bus_ff_103 <= io_i_mux_bus_103;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_104 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_104 <= 1'h0;
    end else begin
      r_mux_bus_ff_104 <= io_i_mux_bus_104;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_105 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_105 <= 1'h0;
    end else begin
      r_mux_bus_ff_105 <= io_i_mux_bus_105;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_106 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_106 <= 1'h0;
    end else begin
      r_mux_bus_ff_106 <= io_i_mux_bus_106;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_107 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_107 <= 1'h0;
    end else begin
      r_mux_bus_ff_107 <= io_i_mux_bus_107;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_108 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_108 <= 1'h0;
    end else begin
      r_mux_bus_ff_108 <= io_i_mux_bus_108;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_109 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_109 <= 1'h0;
    end else begin
      r_mux_bus_ff_109 <= io_i_mux_bus_109;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_110 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_110 <= 1'h0;
    end else begin
      r_mux_bus_ff_110 <= io_i_mux_bus_110;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_111 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_111 <= 1'h0;
    end else begin
      r_mux_bus_ff_111 <= io_i_mux_bus_111;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_112 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_112 <= 1'h0;
    end else begin
      r_mux_bus_ff_112 <= io_i_mux_bus_112;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_113 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_113 <= 1'h0;
    end else begin
      r_mux_bus_ff_113 <= io_i_mux_bus_113;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_114 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_114 <= 1'h0;
    end else begin
      r_mux_bus_ff_114 <= io_i_mux_bus_114;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_115 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_115 <= 1'h0;
    end else begin
      r_mux_bus_ff_115 <= io_i_mux_bus_115;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_116 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_116 <= 1'h0;
    end else begin
      r_mux_bus_ff_116 <= io_i_mux_bus_116;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_117 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_117 <= 1'h0;
    end else begin
      r_mux_bus_ff_117 <= io_i_mux_bus_117;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_118 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_118 <= 1'h0;
    end else begin
      r_mux_bus_ff_118 <= io_i_mux_bus_118;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_119 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_119 <= 1'h0;
    end else begin
      r_mux_bus_ff_119 <= io_i_mux_bus_119;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_120 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_120 <= 1'h0;
    end else begin
      r_mux_bus_ff_120 <= io_i_mux_bus_120;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_121 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_121 <= 1'h0;
    end else begin
      r_mux_bus_ff_121 <= io_i_mux_bus_121;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_122 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_122 <= 1'h0;
    end else begin
      r_mux_bus_ff_122 <= io_i_mux_bus_122;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_123 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_123 <= 1'h0;
    end else begin
      r_mux_bus_ff_123 <= io_i_mux_bus_123;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_124 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_124 <= 1'h0;
    end else begin
      r_mux_bus_ff_124 <= io_i_mux_bus_124;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_125 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_125 <= 1'h0;
    end else begin
      r_mux_bus_ff_125 <= io_i_mux_bus_125;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_126 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_126 <= 1'h0;
    end else begin
      r_mux_bus_ff_126 <= io_i_mux_bus_126;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_127 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_127 <= 1'h0;
    end else begin
      r_mux_bus_ff_127 <= io_i_mux_bus_127;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_128 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_128 <= 1'h0;
    end else begin
      r_mux_bus_ff_128 <= io_i_mux_bus_128;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_129 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_129 <= 1'h0;
    end else begin
      r_mux_bus_ff_129 <= io_i_mux_bus_129;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_130 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_130 <= 1'h0;
    end else begin
      r_mux_bus_ff_130 <= io_i_mux_bus_130;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_131 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_131 <= 1'h0;
    end else begin
      r_mux_bus_ff_131 <= io_i_mux_bus_131;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_132 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_132 <= 1'h0;
    end else begin
      r_mux_bus_ff_132 <= io_i_mux_bus_132;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_133 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_133 <= 1'h0;
    end else begin
      r_mux_bus_ff_133 <= io_i_mux_bus_133;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_134 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_134 <= 1'h0;
    end else begin
      r_mux_bus_ff_134 <= io_i_mux_bus_134;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_135 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_135 <= 1'h0;
    end else begin
      r_mux_bus_ff_135 <= io_i_mux_bus_135;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_136 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_136 <= 1'h0;
    end else begin
      r_mux_bus_ff_136 <= io_i_mux_bus_136;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_137 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_137 <= 1'h0;
    end else begin
      r_mux_bus_ff_137 <= io_i_mux_bus_137;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_138 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_138 <= 1'h0;
    end else begin
      r_mux_bus_ff_138 <= io_i_mux_bus_138;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_139 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_139 <= 1'h0;
    end else begin
      r_mux_bus_ff_139 <= io_i_mux_bus_139;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_140 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_140 <= 1'h0;
    end else begin
      r_mux_bus_ff_140 <= io_i_mux_bus_140;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_141 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_141 <= 1'h0;
    end else begin
      r_mux_bus_ff_141 <= io_i_mux_bus_141;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_142 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_142 <= 1'h0;
    end else begin
      r_mux_bus_ff_142 <= io_i_mux_bus_142;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_143 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_143 <= 1'h0;
    end else begin
      r_mux_bus_ff_143 <= io_i_mux_bus_143;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_144 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_144 <= 1'h0;
    end else begin
      r_mux_bus_ff_144 <= io_i_mux_bus_144;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_145 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_145 <= 1'h0;
    end else begin
      r_mux_bus_ff_145 <= io_i_mux_bus_145;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_146 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_146 <= 1'h0;
    end else begin
      r_mux_bus_ff_146 <= io_i_mux_bus_146;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_147 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_147 <= 1'h0;
    end else begin
      r_mux_bus_ff_147 <= io_i_mux_bus_147;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_148 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_148 <= 1'h0;
    end else begin
      r_mux_bus_ff_148 <= io_i_mux_bus_148;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_149 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_149 <= 1'h0;
    end else begin
      r_mux_bus_ff_149 <= io_i_mux_bus_149;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_150 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_150 <= 1'h0;
    end else begin
      r_mux_bus_ff_150 <= io_i_mux_bus_150;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_151 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_151 <= 1'h0;
    end else begin
      r_mux_bus_ff_151 <= io_i_mux_bus_151;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_152 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_152 <= 1'h0;
    end else begin
      r_mux_bus_ff_152 <= io_i_mux_bus_152;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_153 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_153 <= 1'h0;
    end else begin
      r_mux_bus_ff_153 <= io_i_mux_bus_153;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_154 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_154 <= 1'h0;
    end else begin
      r_mux_bus_ff_154 <= io_i_mux_bus_154;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_155 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_155 <= 1'h0;
    end else begin
      r_mux_bus_ff_155 <= io_i_mux_bus_155;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_156 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_156 <= 1'h0;
    end else begin
      r_mux_bus_ff_156 <= io_i_mux_bus_156;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_157 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_157 <= 1'h0;
    end else begin
      r_mux_bus_ff_157 <= io_i_mux_bus_157;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_158 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_158 <= 1'h0;
    end else begin
      r_mux_bus_ff_158 <= io_i_mux_bus_158;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_159 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_159 <= 1'h0;
    end else begin
      r_mux_bus_ff_159 <= io_i_mux_bus_159;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_160 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_160 <= 1'h0;
    end else begin
      r_mux_bus_ff_160 <= io_i_mux_bus_160;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_161 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_161 <= 1'h0;
    end else begin
      r_mux_bus_ff_161 <= io_i_mux_bus_161;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_162 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_162 <= 1'h0;
    end else begin
      r_mux_bus_ff_162 <= io_i_mux_bus_162;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_163 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_163 <= 1'h0;
    end else begin
      r_mux_bus_ff_163 <= io_i_mux_bus_163;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_164 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_164 <= 1'h0;
    end else begin
      r_mux_bus_ff_164 <= io_i_mux_bus_164;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_165 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_165 <= 1'h0;
    end else begin
      r_mux_bus_ff_165 <= io_i_mux_bus_165;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_166 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_166 <= 1'h0;
    end else begin
      r_mux_bus_ff_166 <= io_i_mux_bus_166;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_167 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_167 <= 1'h0;
    end else begin
      r_mux_bus_ff_167 <= io_i_mux_bus_167;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_168 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_168 <= 1'h0;
    end else begin
      r_mux_bus_ff_168 <= io_i_mux_bus_168;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_169 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_169 <= 1'h0;
    end else begin
      r_mux_bus_ff_169 <= io_i_mux_bus_169;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_170 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_170 <= 1'h0;
    end else begin
      r_mux_bus_ff_170 <= io_i_mux_bus_170;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_171 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_171 <= 1'h0;
    end else begin
      r_mux_bus_ff_171 <= io_i_mux_bus_171;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_172 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_172 <= 1'h0;
    end else begin
      r_mux_bus_ff_172 <= io_i_mux_bus_172;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_173 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_173 <= 1'h0;
    end else begin
      r_mux_bus_ff_173 <= io_i_mux_bus_173;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_174 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_174 <= 1'h0;
    end else begin
      r_mux_bus_ff_174 <= io_i_mux_bus_174;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_175 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_175 <= 1'h0;
    end else begin
      r_mux_bus_ff_175 <= io_i_mux_bus_175;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_176 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_176 <= 1'h0;
    end else begin
      r_mux_bus_ff_176 <= io_i_mux_bus_176;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_177 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_177 <= 1'h0;
    end else begin
      r_mux_bus_ff_177 <= io_i_mux_bus_177;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_178 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_178 <= 1'h0;
    end else begin
      r_mux_bus_ff_178 <= io_i_mux_bus_178;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_179 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_179 <= 1'h0;
    end else begin
      r_mux_bus_ff_179 <= io_i_mux_bus_179;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_180 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_180 <= 1'h0;
    end else begin
      r_mux_bus_ff_180 <= io_i_mux_bus_180;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_181 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_181 <= 1'h0;
    end else begin
      r_mux_bus_ff_181 <= io_i_mux_bus_181;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_182 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_182 <= 1'h0;
    end else begin
      r_mux_bus_ff_182 <= io_i_mux_bus_182;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_183 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_183 <= 1'h0;
    end else begin
      r_mux_bus_ff_183 <= io_i_mux_bus_183;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_184 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_184 <= 1'h0;
    end else begin
      r_mux_bus_ff_184 <= io_i_mux_bus_184;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_185 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_185 <= 1'h0;
    end else begin
      r_mux_bus_ff_185 <= io_i_mux_bus_185;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_186 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_186 <= 1'h0;
    end else begin
      r_mux_bus_ff_186 <= io_i_mux_bus_186;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_187 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_187 <= 1'h0;
    end else begin
      r_mux_bus_ff_187 <= io_i_mux_bus_187;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_188 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_188 <= 1'h0;
    end else begin
      r_mux_bus_ff_188 <= io_i_mux_bus_188;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_189 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_189 <= 1'h0;
    end else begin
      r_mux_bus_ff_189 <= io_i_mux_bus_189;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_190 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_190 <= 1'h0;
    end else begin
      r_mux_bus_ff_190 <= io_i_mux_bus_190;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_191 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_191 <= 1'h0;
    end else begin
      r_mux_bus_ff_191 <= io_i_mux_bus_191;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_192 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_192 <= 1'h0;
    end else begin
      r_mux_bus_ff_192 <= io_i_mux_bus_192;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_193 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_193 <= 1'h0;
    end else begin
      r_mux_bus_ff_193 <= io_i_mux_bus_193;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_194 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_194 <= 1'h0;
    end else begin
      r_mux_bus_ff_194 <= io_i_mux_bus_194;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_195 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_195 <= 1'h0;
    end else begin
      r_mux_bus_ff_195 <= io_i_mux_bus_195;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_196 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_196 <= 1'h0;
    end else begin
      r_mux_bus_ff_196 <= io_i_mux_bus_196;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_197 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_197 <= 1'h0;
    end else begin
      r_mux_bus_ff_197 <= io_i_mux_bus_197;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_198 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_198 <= 1'h0;
    end else begin
      r_mux_bus_ff_198 <= io_i_mux_bus_198;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_199 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_199 <= 1'h0;
    end else begin
      r_mux_bus_ff_199 <= io_i_mux_bus_199;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_200 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_200 <= 1'h0;
    end else begin
      r_mux_bus_ff_200 <= io_i_mux_bus_200;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_201 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_201 <= 1'h0;
    end else begin
      r_mux_bus_ff_201 <= io_i_mux_bus_201;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_202 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_202 <= 1'h0;
    end else begin
      r_mux_bus_ff_202 <= io_i_mux_bus_202;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_203 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_203 <= 1'h0;
    end else begin
      r_mux_bus_ff_203 <= io_i_mux_bus_203;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_204 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_204 <= 1'h0;
    end else begin
      r_mux_bus_ff_204 <= io_i_mux_bus_204;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_205 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_205 <= 1'h0;
    end else begin
      r_mux_bus_ff_205 <= io_i_mux_bus_205;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_206 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_206 <= 1'h0;
    end else begin
      r_mux_bus_ff_206 <= io_i_mux_bus_206;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_207 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_207 <= 1'h0;
    end else begin
      r_mux_bus_ff_207 <= io_i_mux_bus_207;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_208 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_208 <= 1'h0;
    end else begin
      r_mux_bus_ff_208 <= io_i_mux_bus_208;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_209 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_209 <= 1'h0;
    end else begin
      r_mux_bus_ff_209 <= io_i_mux_bus_209;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_210 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_210 <= 1'h0;
    end else begin
      r_mux_bus_ff_210 <= io_i_mux_bus_210;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_211 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_211 <= 1'h0;
    end else begin
      r_mux_bus_ff_211 <= io_i_mux_bus_211;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_212 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_212 <= 1'h0;
    end else begin
      r_mux_bus_ff_212 <= io_i_mux_bus_212;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_213 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_213 <= 1'h0;
    end else begin
      r_mux_bus_ff_213 <= io_i_mux_bus_213;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_214 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_214 <= 1'h0;
    end else begin
      r_mux_bus_ff_214 <= io_i_mux_bus_214;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_215 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_215 <= 1'h0;
    end else begin
      r_mux_bus_ff_215 <= io_i_mux_bus_215;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_216 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_216 <= 1'h0;
    end else begin
      r_mux_bus_ff_216 <= io_i_mux_bus_216;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_217 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_217 <= 1'h0;
    end else begin
      r_mux_bus_ff_217 <= io_i_mux_bus_217;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_218 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_218 <= 1'h0;
    end else begin
      r_mux_bus_ff_218 <= io_i_mux_bus_218;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_219 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_219 <= 1'h0;
    end else begin
      r_mux_bus_ff_219 <= io_i_mux_bus_219;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_220 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_220 <= 1'h0;
    end else begin
      r_mux_bus_ff_220 <= io_i_mux_bus_220;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_221 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_221 <= 1'h0;
    end else begin
      r_mux_bus_ff_221 <= io_i_mux_bus_221;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_222 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_222 <= 1'h0;
    end else begin
      r_mux_bus_ff_222 <= io_i_mux_bus_222;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_223 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_223 <= 1'h0;
    end else begin
      r_mux_bus_ff_223 <= io_i_mux_bus_223;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_224 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_224 <= 1'h0;
    end else begin
      r_mux_bus_ff_224 <= io_i_mux_bus_224;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_225 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_225 <= 1'h0;
    end else begin
      r_mux_bus_ff_225 <= io_i_mux_bus_225;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_226 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_226 <= 1'h0;
    end else begin
      r_mux_bus_ff_226 <= io_i_mux_bus_226;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_227 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_227 <= 1'h0;
    end else begin
      r_mux_bus_ff_227 <= io_i_mux_bus_227;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_228 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_228 <= 1'h0;
    end else begin
      r_mux_bus_ff_228 <= io_i_mux_bus_228;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_229 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_229 <= 1'h0;
    end else begin
      r_mux_bus_ff_229 <= io_i_mux_bus_229;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_230 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_230 <= 1'h0;
    end else begin
      r_mux_bus_ff_230 <= io_i_mux_bus_230;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_231 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_231 <= 1'h0;
    end else begin
      r_mux_bus_ff_231 <= io_i_mux_bus_231;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_232 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_232 <= 1'h0;
    end else begin
      r_mux_bus_ff_232 <= io_i_mux_bus_232;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_233 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_233 <= 1'h0;
    end else begin
      r_mux_bus_ff_233 <= io_i_mux_bus_233;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_234 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_234 <= 1'h0;
    end else begin
      r_mux_bus_ff_234 <= io_i_mux_bus_234;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_235 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_235 <= 1'h0;
    end else begin
      r_mux_bus_ff_235 <= io_i_mux_bus_235;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_236 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_236 <= 1'h0;
    end else begin
      r_mux_bus_ff_236 <= io_i_mux_bus_236;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_237 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_237 <= 1'h0;
    end else begin
      r_mux_bus_ff_237 <= io_i_mux_bus_237;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_238 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_238 <= 1'h0;
    end else begin
      r_mux_bus_ff_238 <= io_i_mux_bus_238;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_239 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_239 <= 1'h0;
    end else begin
      r_mux_bus_ff_239 <= io_i_mux_bus_239;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_240 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_240 <= 1'h0;
    end else begin
      r_mux_bus_ff_240 <= io_i_mux_bus_240;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_241 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_241 <= 1'h0;
    end else begin
      r_mux_bus_ff_241 <= io_i_mux_bus_241;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_242 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_242 <= 1'h0;
    end else begin
      r_mux_bus_ff_242 <= io_i_mux_bus_242;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_243 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_243 <= 1'h0;
    end else begin
      r_mux_bus_ff_243 <= io_i_mux_bus_243;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_244 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_244 <= 1'h0;
    end else begin
      r_mux_bus_ff_244 <= io_i_mux_bus_244;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_245 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_245 <= 1'h0;
    end else begin
      r_mux_bus_ff_245 <= io_i_mux_bus_245;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_246 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_246 <= 1'h0;
    end else begin
      r_mux_bus_ff_246 <= io_i_mux_bus_246;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_247 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_247 <= 1'h0;
    end else begin
      r_mux_bus_ff_247 <= io_i_mux_bus_247;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_248 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_248 <= 1'h0;
    end else begin
      r_mux_bus_ff_248 <= io_i_mux_bus_248;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_249 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_249 <= 1'h0;
    end else begin
      r_mux_bus_ff_249 <= io_i_mux_bus_249;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_250 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_250 <= 1'h0;
    end else begin
      r_mux_bus_ff_250 <= io_i_mux_bus_250;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_251 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_251 <= 1'h0;
    end else begin
      r_mux_bus_ff_251 <= io_i_mux_bus_251;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_252 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_252 <= 1'h0;
    end else begin
      r_mux_bus_ff_252 <= io_i_mux_bus_252;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_253 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_253 <= 1'h0;
    end else begin
      r_mux_bus_ff_253 <= io_i_mux_bus_253;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_254 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_254 <= 1'h0;
    end else begin
      r_mux_bus_ff_254 <= io_i_mux_bus_254;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_255 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_255 <= 1'h0;
    end else begin
      r_mux_bus_ff_255 <= io_i_mux_bus_255;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_256 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_256 <= 1'h0;
    end else begin
      r_mux_bus_ff_256 <= io_i_mux_bus_256;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_257 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_257 <= 1'h0;
    end else begin
      r_mux_bus_ff_257 <= io_i_mux_bus_257;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_258 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_258 <= 1'h0;
    end else begin
      r_mux_bus_ff_258 <= io_i_mux_bus_258;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_259 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_259 <= 1'h0;
    end else begin
      r_mux_bus_ff_259 <= io_i_mux_bus_259;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_260 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_260 <= 1'h0;
    end else begin
      r_mux_bus_ff_260 <= io_i_mux_bus_260;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_261 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_261 <= 1'h0;
    end else begin
      r_mux_bus_ff_261 <= io_i_mux_bus_261;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_262 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_262 <= 1'h0;
    end else begin
      r_mux_bus_ff_262 <= io_i_mux_bus_262;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_263 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_263 <= 1'h0;
    end else begin
      r_mux_bus_ff_263 <= io_i_mux_bus_263;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_264 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_264 <= 1'h0;
    end else begin
      r_mux_bus_ff_264 <= io_i_mux_bus_264;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_265 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_265 <= 1'h0;
    end else begin
      r_mux_bus_ff_265 <= io_i_mux_bus_265;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_266 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_266 <= 1'h0;
    end else begin
      r_mux_bus_ff_266 <= io_i_mux_bus_266;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_267 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_267 <= 1'h0;
    end else begin
      r_mux_bus_ff_267 <= io_i_mux_bus_267;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_268 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_268 <= 1'h0;
    end else begin
      r_mux_bus_ff_268 <= io_i_mux_bus_268;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_269 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_269 <= 1'h0;
    end else begin
      r_mux_bus_ff_269 <= io_i_mux_bus_269;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_270 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_270 <= 1'h0;
    end else begin
      r_mux_bus_ff_270 <= io_i_mux_bus_270;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_271 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_271 <= 1'h0;
    end else begin
      r_mux_bus_ff_271 <= io_i_mux_bus_271;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_272 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_272 <= 1'h0;
    end else begin
      r_mux_bus_ff_272 <= io_i_mux_bus_272;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_273 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_273 <= 1'h0;
    end else begin
      r_mux_bus_ff_273 <= io_i_mux_bus_273;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_274 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_274 <= 1'h0;
    end else begin
      r_mux_bus_ff_274 <= io_i_mux_bus_274;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_275 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_275 <= 1'h0;
    end else begin
      r_mux_bus_ff_275 <= io_i_mux_bus_275;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_276 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_276 <= 1'h0;
    end else begin
      r_mux_bus_ff_276 <= io_i_mux_bus_276;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_277 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_277 <= 1'h0;
    end else begin
      r_mux_bus_ff_277 <= io_i_mux_bus_277;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_278 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_278 <= 1'h0;
    end else begin
      r_mux_bus_ff_278 <= io_i_mux_bus_278;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_279 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_279 <= 1'h0;
    end else begin
      r_mux_bus_ff_279 <= io_i_mux_bus_279;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_280 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_280 <= 1'h0;
    end else begin
      r_mux_bus_ff_280 <= io_i_mux_bus_280;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_281 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_281 <= 1'h0;
    end else begin
      r_mux_bus_ff_281 <= io_i_mux_bus_281;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_282 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_282 <= 1'h0;
    end else begin
      r_mux_bus_ff_282 <= io_i_mux_bus_282;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_283 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_283 <= 1'h0;
    end else begin
      r_mux_bus_ff_283 <= io_i_mux_bus_283;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_284 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_284 <= 1'h0;
    end else begin
      r_mux_bus_ff_284 <= io_i_mux_bus_284;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_285 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_285 <= 1'h0;
    end else begin
      r_mux_bus_ff_285 <= io_i_mux_bus_285;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_286 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_286 <= 1'h0;
    end else begin
      r_mux_bus_ff_286 <= io_i_mux_bus_286;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_287 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_287 <= 1'h0;
    end else begin
      r_mux_bus_ff_287 <= io_i_mux_bus_287;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_288 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_288 <= 1'h0;
    end else begin
      r_mux_bus_ff_288 <= io_i_mux_bus_288;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_289 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_289 <= 1'h0;
    end else begin
      r_mux_bus_ff_289 <= io_i_mux_bus_289;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_290 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_290 <= 1'h0;
    end else begin
      r_mux_bus_ff_290 <= io_i_mux_bus_290;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_291 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_291 <= 1'h0;
    end else begin
      r_mux_bus_ff_291 <= io_i_mux_bus_291;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_292 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_292 <= 1'h0;
    end else begin
      r_mux_bus_ff_292 <= io_i_mux_bus_292;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_293 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_293 <= 1'h0;
    end else begin
      r_mux_bus_ff_293 <= io_i_mux_bus_293;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_294 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_294 <= 1'h0;
    end else begin
      r_mux_bus_ff_294 <= io_i_mux_bus_294;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_295 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_295 <= 1'h0;
    end else begin
      r_mux_bus_ff_295 <= io_i_mux_bus_295;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_296 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_296 <= 1'h0;
    end else begin
      r_mux_bus_ff_296 <= io_i_mux_bus_296;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_297 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_297 <= 1'h0;
    end else begin
      r_mux_bus_ff_297 <= io_i_mux_bus_297;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_298 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_298 <= 1'h0;
    end else begin
      r_mux_bus_ff_298 <= io_i_mux_bus_298;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_299 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_299 <= 1'h0;
    end else begin
      r_mux_bus_ff_299 <= io_i_mux_bus_299;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_300 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_300 <= 1'h0;
    end else begin
      r_mux_bus_ff_300 <= io_i_mux_bus_300;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_301 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_301 <= 1'h0;
    end else begin
      r_mux_bus_ff_301 <= io_i_mux_bus_301;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_302 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_302 <= 1'h0;
    end else begin
      r_mux_bus_ff_302 <= io_i_mux_bus_302;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_303 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_303 <= 1'h0;
    end else begin
      r_mux_bus_ff_303 <= io_i_mux_bus_303;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_304 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_304 <= 1'h0;
    end else begin
      r_mux_bus_ff_304 <= io_i_mux_bus_304;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_305 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_305 <= 1'h0;
    end else begin
      r_mux_bus_ff_305 <= io_i_mux_bus_305;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_306 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_306 <= 1'h0;
    end else begin
      r_mux_bus_ff_306 <= io_i_mux_bus_306;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_307 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_307 <= 1'h0;
    end else begin
      r_mux_bus_ff_307 <= io_i_mux_bus_307;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_308 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_308 <= 1'h0;
    end else begin
      r_mux_bus_ff_308 <= io_i_mux_bus_308;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_309 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_309 <= 1'h0;
    end else begin
      r_mux_bus_ff_309 <= io_i_mux_bus_309;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_310 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_310 <= 1'h0;
    end else begin
      r_mux_bus_ff_310 <= io_i_mux_bus_310;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_311 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_311 <= 1'h0;
    end else begin
      r_mux_bus_ff_311 <= io_i_mux_bus_311;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_312 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_312 <= 1'h0;
    end else begin
      r_mux_bus_ff_312 <= io_i_mux_bus_312;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_313 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_313 <= 1'h0;
    end else begin
      r_mux_bus_ff_313 <= io_i_mux_bus_313;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_314 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_314 <= 1'h0;
    end else begin
      r_mux_bus_ff_314 <= io_i_mux_bus_314;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_315 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_315 <= 1'h0;
    end else begin
      r_mux_bus_ff_315 <= io_i_mux_bus_315;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_316 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_316 <= 1'h0;
    end else begin
      r_mux_bus_ff_316 <= io_i_mux_bus_316;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_317 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_317 <= 1'h0;
    end else begin
      r_mux_bus_ff_317 <= io_i_mux_bus_317;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_318 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_318 <= 1'h0;
    end else begin
      r_mux_bus_ff_318 <= io_i_mux_bus_318;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_319 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_319 <= 1'h0;
    end else begin
      r_mux_bus_ff_319 <= io_i_mux_bus_319;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_320 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_320 <= 1'h0;
    end else begin
      r_mux_bus_ff_320 <= io_i_mux_bus_320;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_321 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_321 <= 1'h0;
    end else begin
      r_mux_bus_ff_321 <= io_i_mux_bus_321;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_322 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_322 <= 1'h0;
    end else begin
      r_mux_bus_ff_322 <= io_i_mux_bus_322;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_323 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_323 <= 1'h0;
    end else begin
      r_mux_bus_ff_323 <= io_i_mux_bus_323;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_324 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_324 <= 1'h0;
    end else begin
      r_mux_bus_ff_324 <= io_i_mux_bus_324;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_325 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_325 <= 1'h0;
    end else begin
      r_mux_bus_ff_325 <= io_i_mux_bus_325;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_326 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_326 <= 1'h0;
    end else begin
      r_mux_bus_ff_326 <= io_i_mux_bus_326;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_327 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_327 <= 1'h0;
    end else begin
      r_mux_bus_ff_327 <= io_i_mux_bus_327;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_328 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_328 <= 1'h0;
    end else begin
      r_mux_bus_ff_328 <= io_i_mux_bus_328;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_329 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_329 <= 1'h0;
    end else begin
      r_mux_bus_ff_329 <= io_i_mux_bus_329;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_330 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_330 <= 1'h0;
    end else begin
      r_mux_bus_ff_330 <= io_i_mux_bus_330;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_331 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_331 <= 1'h0;
    end else begin
      r_mux_bus_ff_331 <= io_i_mux_bus_331;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_332 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_332 <= 1'h0;
    end else begin
      r_mux_bus_ff_332 <= io_i_mux_bus_332;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_333 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_333 <= 1'h0;
    end else begin
      r_mux_bus_ff_333 <= io_i_mux_bus_333;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_334 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_334 <= 1'h0;
    end else begin
      r_mux_bus_ff_334 <= io_i_mux_bus_334;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_335 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_335 <= 1'h0;
    end else begin
      r_mux_bus_ff_335 <= io_i_mux_bus_335;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_336 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_336 <= 1'h0;
    end else begin
      r_mux_bus_ff_336 <= io_i_mux_bus_336;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_337 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_337 <= 1'h0;
    end else begin
      r_mux_bus_ff_337 <= io_i_mux_bus_337;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_338 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_338 <= 1'h0;
    end else begin
      r_mux_bus_ff_338 <= io_i_mux_bus_338;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_339 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_339 <= 1'h0;
    end else begin
      r_mux_bus_ff_339 <= io_i_mux_bus_339;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_340 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_340 <= 1'h0;
    end else begin
      r_mux_bus_ff_340 <= io_i_mux_bus_340;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_341 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_341 <= 1'h0;
    end else begin
      r_mux_bus_ff_341 <= io_i_mux_bus_341;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_342 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_342 <= 1'h0;
    end else begin
      r_mux_bus_ff_342 <= io_i_mux_bus_342;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_343 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_343 <= 1'h0;
    end else begin
      r_mux_bus_ff_343 <= io_i_mux_bus_343;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_344 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_344 <= 1'h0;
    end else begin
      r_mux_bus_ff_344 <= io_i_mux_bus_344;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_345 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_345 <= 1'h0;
    end else begin
      r_mux_bus_ff_345 <= io_i_mux_bus_345;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_346 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_346 <= 1'h0;
    end else begin
      r_mux_bus_ff_346 <= io_i_mux_bus_346;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_347 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_347 <= 1'h0;
    end else begin
      r_mux_bus_ff_347 <= io_i_mux_bus_347;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_348 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_348 <= 1'h0;
    end else begin
      r_mux_bus_ff_348 <= io_i_mux_bus_348;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_349 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_349 <= 1'h0;
    end else begin
      r_mux_bus_ff_349 <= io_i_mux_bus_349;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_350 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_350 <= 1'h0;
    end else begin
      r_mux_bus_ff_350 <= io_i_mux_bus_350;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_351 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_351 <= 1'h0;
    end else begin
      r_mux_bus_ff_351 <= io_i_mux_bus_351;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_352 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_352 <= 1'h0;
    end else begin
      r_mux_bus_ff_352 <= io_i_mux_bus_352;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_353 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_353 <= 1'h0;
    end else begin
      r_mux_bus_ff_353 <= io_i_mux_bus_353;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_354 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_354 <= 1'h0;
    end else begin
      r_mux_bus_ff_354 <= io_i_mux_bus_354;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_355 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_355 <= 1'h0;
    end else begin
      r_mux_bus_ff_355 <= io_i_mux_bus_355;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_356 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_356 <= 1'h0;
    end else begin
      r_mux_bus_ff_356 <= io_i_mux_bus_356;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_357 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_357 <= 1'h0;
    end else begin
      r_mux_bus_ff_357 <= io_i_mux_bus_357;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_358 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_358 <= 1'h0;
    end else begin
      r_mux_bus_ff_358 <= io_i_mux_bus_358;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_359 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_359 <= 1'h0;
    end else begin
      r_mux_bus_ff_359 <= io_i_mux_bus_359;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_360 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_360 <= 1'h0;
    end else begin
      r_mux_bus_ff_360 <= io_i_mux_bus_360;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_361 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_361 <= 1'h0;
    end else begin
      r_mux_bus_ff_361 <= io_i_mux_bus_361;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_362 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_362 <= 1'h0;
    end else begin
      r_mux_bus_ff_362 <= io_i_mux_bus_362;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_363 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_363 <= 1'h0;
    end else begin
      r_mux_bus_ff_363 <= io_i_mux_bus_363;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_364 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_364 <= 1'h0;
    end else begin
      r_mux_bus_ff_364 <= io_i_mux_bus_364;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_365 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_365 <= 1'h0;
    end else begin
      r_mux_bus_ff_365 <= io_i_mux_bus_365;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_366 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_366 <= 1'h0;
    end else begin
      r_mux_bus_ff_366 <= io_i_mux_bus_366;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_367 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_367 <= 1'h0;
    end else begin
      r_mux_bus_ff_367 <= io_i_mux_bus_367;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_368 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_368 <= 1'h0;
    end else begin
      r_mux_bus_ff_368 <= io_i_mux_bus_368;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_369 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_369 <= 1'h0;
    end else begin
      r_mux_bus_ff_369 <= io_i_mux_bus_369;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_370 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_370 <= 1'h0;
    end else begin
      r_mux_bus_ff_370 <= io_i_mux_bus_370;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_371 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_371 <= 1'h0;
    end else begin
      r_mux_bus_ff_371 <= io_i_mux_bus_371;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_372 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_372 <= 1'h0;
    end else begin
      r_mux_bus_ff_372 <= io_i_mux_bus_372;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_373 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_373 <= 1'h0;
    end else begin
      r_mux_bus_ff_373 <= io_i_mux_bus_373;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_374 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_374 <= 1'h0;
    end else begin
      r_mux_bus_ff_374 <= io_i_mux_bus_374;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_375 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_375 <= 1'h0;
    end else begin
      r_mux_bus_ff_375 <= io_i_mux_bus_375;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_376 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_376 <= 1'h0;
    end else begin
      r_mux_bus_ff_376 <= io_i_mux_bus_376;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_377 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_377 <= 1'h0;
    end else begin
      r_mux_bus_ff_377 <= io_i_mux_bus_377;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_378 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_378 <= 1'h0;
    end else begin
      r_mux_bus_ff_378 <= io_i_mux_bus_378;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_379 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_379 <= 1'h0;
    end else begin
      r_mux_bus_ff_379 <= io_i_mux_bus_379;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_380 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_380 <= 1'h0;
    end else begin
      r_mux_bus_ff_380 <= io_i_mux_bus_380;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_381 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_381 <= 1'h0;
    end else begin
      r_mux_bus_ff_381 <= io_i_mux_bus_381;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_382 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_382 <= 1'h0;
    end else begin
      r_mux_bus_ff_382 <= io_i_mux_bus_382;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_383 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_383 <= 1'h0;
    end else begin
      r_mux_bus_ff_383 <= io_i_mux_bus_383;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_384 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_384 <= 1'h0;
    end else begin
      r_mux_bus_ff_384 <= io_i_mux_bus_384;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_385 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_385 <= 1'h0;
    end else begin
      r_mux_bus_ff_385 <= io_i_mux_bus_385;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_386 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_386 <= 1'h0;
    end else begin
      r_mux_bus_ff_386 <= io_i_mux_bus_386;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_387 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_387 <= 1'h0;
    end else begin
      r_mux_bus_ff_387 <= io_i_mux_bus_387;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_388 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_388 <= 1'h0;
    end else begin
      r_mux_bus_ff_388 <= io_i_mux_bus_388;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_389 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_389 <= 1'h0;
    end else begin
      r_mux_bus_ff_389 <= io_i_mux_bus_389;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_390 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_390 <= 1'h0;
    end else begin
      r_mux_bus_ff_390 <= io_i_mux_bus_390;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_391 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_391 <= 1'h0;
    end else begin
      r_mux_bus_ff_391 <= io_i_mux_bus_391;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_392 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_392 <= 1'h0;
    end else begin
      r_mux_bus_ff_392 <= io_i_mux_bus_392;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_393 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_393 <= 1'h0;
    end else begin
      r_mux_bus_ff_393 <= io_i_mux_bus_393;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_394 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_394 <= 1'h0;
    end else begin
      r_mux_bus_ff_394 <= io_i_mux_bus_394;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_395 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_395 <= 1'h0;
    end else begin
      r_mux_bus_ff_395 <= io_i_mux_bus_395;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_396 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_396 <= 1'h0;
    end else begin
      r_mux_bus_ff_396 <= io_i_mux_bus_396;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_397 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_397 <= 1'h0;
    end else begin
      r_mux_bus_ff_397 <= io_i_mux_bus_397;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_398 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_398 <= 1'h0;
    end else begin
      r_mux_bus_ff_398 <= io_i_mux_bus_398;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_399 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_399 <= 1'h0;
    end else begin
      r_mux_bus_ff_399 <= io_i_mux_bus_399;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_400 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_400 <= 1'h0;
    end else begin
      r_mux_bus_ff_400 <= io_i_mux_bus_400;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_401 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_401 <= 1'h0;
    end else begin
      r_mux_bus_ff_401 <= io_i_mux_bus_401;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_402 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_402 <= 1'h0;
    end else begin
      r_mux_bus_ff_402 <= io_i_mux_bus_402;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_403 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_403 <= 1'h0;
    end else begin
      r_mux_bus_ff_403 <= io_i_mux_bus_403;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_404 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_404 <= 1'h0;
    end else begin
      r_mux_bus_ff_404 <= io_i_mux_bus_404;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_405 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_405 <= 1'h0;
    end else begin
      r_mux_bus_ff_405 <= io_i_mux_bus_405;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_406 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_406 <= 1'h0;
    end else begin
      r_mux_bus_ff_406 <= io_i_mux_bus_406;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_407 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_407 <= 1'h0;
    end else begin
      r_mux_bus_ff_407 <= io_i_mux_bus_407;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_408 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_408 <= 1'h0;
    end else begin
      r_mux_bus_ff_408 <= io_i_mux_bus_408;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_409 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_409 <= 1'h0;
    end else begin
      r_mux_bus_ff_409 <= io_i_mux_bus_409;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_410 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_410 <= 1'h0;
    end else begin
      r_mux_bus_ff_410 <= io_i_mux_bus_410;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_411 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_411 <= 1'h0;
    end else begin
      r_mux_bus_ff_411 <= io_i_mux_bus_411;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_412 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_412 <= 1'h0;
    end else begin
      r_mux_bus_ff_412 <= io_i_mux_bus_412;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_413 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_413 <= 1'h0;
    end else begin
      r_mux_bus_ff_413 <= io_i_mux_bus_413;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_414 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_414 <= 1'h0;
    end else begin
      r_mux_bus_ff_414 <= io_i_mux_bus_414;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_415 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_415 <= 1'h0;
    end else begin
      r_mux_bus_ff_415 <= io_i_mux_bus_415;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_416 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_416 <= 1'h0;
    end else begin
      r_mux_bus_ff_416 <= io_i_mux_bus_416;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_417 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_417 <= 1'h0;
    end else begin
      r_mux_bus_ff_417 <= io_i_mux_bus_417;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_418 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_418 <= 1'h0;
    end else begin
      r_mux_bus_ff_418 <= io_i_mux_bus_418;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_419 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_419 <= 1'h0;
    end else begin
      r_mux_bus_ff_419 <= io_i_mux_bus_419;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_420 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_420 <= 1'h0;
    end else begin
      r_mux_bus_ff_420 <= io_i_mux_bus_420;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_421 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_421 <= 1'h0;
    end else begin
      r_mux_bus_ff_421 <= io_i_mux_bus_421;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_422 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_422 <= 1'h0;
    end else begin
      r_mux_bus_ff_422 <= io_i_mux_bus_422;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_423 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_423 <= 1'h0;
    end else begin
      r_mux_bus_ff_423 <= io_i_mux_bus_423;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_424 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_424 <= 1'h0;
    end else begin
      r_mux_bus_ff_424 <= io_i_mux_bus_424;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_425 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_425 <= 1'h0;
    end else begin
      r_mux_bus_ff_425 <= io_i_mux_bus_425;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_426 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_426 <= 1'h0;
    end else begin
      r_mux_bus_ff_426 <= io_i_mux_bus_426;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_427 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_427 <= 1'h0;
    end else begin
      r_mux_bus_ff_427 <= io_i_mux_bus_427;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_428 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_428 <= 1'h0;
    end else begin
      r_mux_bus_ff_428 <= io_i_mux_bus_428;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_429 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_429 <= 1'h0;
    end else begin
      r_mux_bus_ff_429 <= io_i_mux_bus_429;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_430 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_430 <= 1'h0;
    end else begin
      r_mux_bus_ff_430 <= io_i_mux_bus_430;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_431 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_431 <= 1'h0;
    end else begin
      r_mux_bus_ff_431 <= io_i_mux_bus_431;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_432 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_432 <= 1'h0;
    end else begin
      r_mux_bus_ff_432 <= io_i_mux_bus_432;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_433 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_433 <= 1'h0;
    end else begin
      r_mux_bus_ff_433 <= io_i_mux_bus_433;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_434 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_434 <= 1'h0;
    end else begin
      r_mux_bus_ff_434 <= io_i_mux_bus_434;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_435 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_435 <= 1'h0;
    end else begin
      r_mux_bus_ff_435 <= io_i_mux_bus_435;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_436 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_436 <= 1'h0;
    end else begin
      r_mux_bus_ff_436 <= io_i_mux_bus_436;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_437 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_437 <= 1'h0;
    end else begin
      r_mux_bus_ff_437 <= io_i_mux_bus_437;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_438 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_438 <= 1'h0;
    end else begin
      r_mux_bus_ff_438 <= io_i_mux_bus_438;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_439 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_439 <= 1'h0;
    end else begin
      r_mux_bus_ff_439 <= io_i_mux_bus_439;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_440 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_440 <= 1'h0;
    end else begin
      r_mux_bus_ff_440 <= io_i_mux_bus_440;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_441 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_441 <= 1'h0;
    end else begin
      r_mux_bus_ff_441 <= io_i_mux_bus_441;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_442 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_442 <= 1'h0;
    end else begin
      r_mux_bus_ff_442 <= io_i_mux_bus_442;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_443 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_443 <= 1'h0;
    end else begin
      r_mux_bus_ff_443 <= io_i_mux_bus_443;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_444 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_444 <= 1'h0;
    end else begin
      r_mux_bus_ff_444 <= io_i_mux_bus_444;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_445 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_445 <= 1'h0;
    end else begin
      r_mux_bus_ff_445 <= io_i_mux_bus_445;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_446 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_446 <= 1'h0;
    end else begin
      r_mux_bus_ff_446 <= io_i_mux_bus_446;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_447 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_447 <= 1'h0;
    end else begin
      r_mux_bus_ff_447 <= io_i_mux_bus_447;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_448 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_448 <= 1'h0;
    end else begin
      r_mux_bus_ff_448 <= io_i_mux_bus_448;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_449 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_449 <= 1'h0;
    end else begin
      r_mux_bus_ff_449 <= io_i_mux_bus_449;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_450 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_450 <= 1'h0;
    end else begin
      r_mux_bus_ff_450 <= io_i_mux_bus_450;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_451 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_451 <= 1'h0;
    end else begin
      r_mux_bus_ff_451 <= io_i_mux_bus_451;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_452 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_452 <= 1'h0;
    end else begin
      r_mux_bus_ff_452 <= io_i_mux_bus_452;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_453 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_453 <= 1'h0;
    end else begin
      r_mux_bus_ff_453 <= io_i_mux_bus_453;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_454 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_454 <= 1'h0;
    end else begin
      r_mux_bus_ff_454 <= io_i_mux_bus_454;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_455 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_455 <= 1'h0;
    end else begin
      r_mux_bus_ff_455 <= io_i_mux_bus_455;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_456 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_456 <= 1'h0;
    end else begin
      r_mux_bus_ff_456 <= io_i_mux_bus_456;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_457 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_457 <= 1'h0;
    end else begin
      r_mux_bus_ff_457 <= io_i_mux_bus_457;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_458 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_458 <= 1'h0;
    end else begin
      r_mux_bus_ff_458 <= io_i_mux_bus_458;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_459 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_459 <= 1'h0;
    end else begin
      r_mux_bus_ff_459 <= io_i_mux_bus_459;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_460 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_460 <= 1'h0;
    end else begin
      r_mux_bus_ff_460 <= io_i_mux_bus_460;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_461 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_461 <= 1'h0;
    end else begin
      r_mux_bus_ff_461 <= io_i_mux_bus_461;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_462 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_462 <= 1'h0;
    end else begin
      r_mux_bus_ff_462 <= io_i_mux_bus_462;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_463 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_463 <= 1'h0;
    end else begin
      r_mux_bus_ff_463 <= io_i_mux_bus_463;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_464 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_464 <= 1'h0;
    end else begin
      r_mux_bus_ff_464 <= io_i_mux_bus_464;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_465 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_465 <= 1'h0;
    end else begin
      r_mux_bus_ff_465 <= io_i_mux_bus_465;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_466 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_466 <= 1'h0;
    end else begin
      r_mux_bus_ff_466 <= io_i_mux_bus_466;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_467 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_467 <= 1'h0;
    end else begin
      r_mux_bus_ff_467 <= io_i_mux_bus_467;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_468 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_468 <= 1'h0;
    end else begin
      r_mux_bus_ff_468 <= io_i_mux_bus_468;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_469 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_469 <= 1'h0;
    end else begin
      r_mux_bus_ff_469 <= io_i_mux_bus_469;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_470 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_470 <= 1'h0;
    end else begin
      r_mux_bus_ff_470 <= io_i_mux_bus_470;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_471 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_471 <= 1'h0;
    end else begin
      r_mux_bus_ff_471 <= io_i_mux_bus_471;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_472 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_472 <= 1'h0;
    end else begin
      r_mux_bus_ff_472 <= io_i_mux_bus_472;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_473 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_473 <= 1'h0;
    end else begin
      r_mux_bus_ff_473 <= io_i_mux_bus_473;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_474 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_474 <= 1'h0;
    end else begin
      r_mux_bus_ff_474 <= io_i_mux_bus_474;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_475 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_475 <= 1'h0;
    end else begin
      r_mux_bus_ff_475 <= io_i_mux_bus_475;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_476 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_476 <= 1'h0;
    end else begin
      r_mux_bus_ff_476 <= io_i_mux_bus_476;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_477 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_477 <= 1'h0;
    end else begin
      r_mux_bus_ff_477 <= io_i_mux_bus_477;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_478 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_478 <= 1'h0;
    end else begin
      r_mux_bus_ff_478 <= io_i_mux_bus_478;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_479 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_479 <= 1'h0;
    end else begin
      r_mux_bus_ff_479 <= io_i_mux_bus_479;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_480 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_480 <= 1'h0;
    end else begin
      r_mux_bus_ff_480 <= io_i_mux_bus_480;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_481 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_481 <= 1'h0;
    end else begin
      r_mux_bus_ff_481 <= io_i_mux_bus_481;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_482 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_482 <= 1'h0;
    end else begin
      r_mux_bus_ff_482 <= io_i_mux_bus_482;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_483 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_483 <= 1'h0;
    end else begin
      r_mux_bus_ff_483 <= io_i_mux_bus_483;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_484 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_484 <= 1'h0;
    end else begin
      r_mux_bus_ff_484 <= io_i_mux_bus_484;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_485 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_485 <= 1'h0;
    end else begin
      r_mux_bus_ff_485 <= io_i_mux_bus_485;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_486 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_486 <= 1'h0;
    end else begin
      r_mux_bus_ff_486 <= io_i_mux_bus_486;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_487 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_487 <= 1'h0;
    end else begin
      r_mux_bus_ff_487 <= io_i_mux_bus_487;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_488 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_488 <= 1'h0;
    end else begin
      r_mux_bus_ff_488 <= io_i_mux_bus_488;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_489 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_489 <= 1'h0;
    end else begin
      r_mux_bus_ff_489 <= io_i_mux_bus_489;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_490 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_490 <= 1'h0;
    end else begin
      r_mux_bus_ff_490 <= io_i_mux_bus_490;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_491 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_491 <= 1'h0;
    end else begin
      r_mux_bus_ff_491 <= io_i_mux_bus_491;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_492 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_492 <= 1'h0;
    end else begin
      r_mux_bus_ff_492 <= io_i_mux_bus_492;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_493 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_493 <= 1'h0;
    end else begin
      r_mux_bus_ff_493 <= io_i_mux_bus_493;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_494 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_494 <= 1'h0;
    end else begin
      r_mux_bus_ff_494 <= io_i_mux_bus_494;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_495 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_495 <= 1'h0;
    end else begin
      r_mux_bus_ff_495 <= io_i_mux_bus_495;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_496 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_496 <= 1'h0;
    end else begin
      r_mux_bus_ff_496 <= io_i_mux_bus_496;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_497 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_497 <= 1'h0;
    end else begin
      r_mux_bus_ff_497 <= io_i_mux_bus_497;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_498 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_498 <= 1'h0;
    end else begin
      r_mux_bus_ff_498 <= io_i_mux_bus_498;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_499 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_499 <= 1'h0;
    end else begin
      r_mux_bus_ff_499 <= io_i_mux_bus_499;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_500 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_500 <= 1'h0;
    end else begin
      r_mux_bus_ff_500 <= io_i_mux_bus_500;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_501 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_501 <= 1'h0;
    end else begin
      r_mux_bus_ff_501 <= io_i_mux_bus_501;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_502 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_502 <= 1'h0;
    end else begin
      r_mux_bus_ff_502 <= io_i_mux_bus_502;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_503 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_503 <= 1'h0;
    end else begin
      r_mux_bus_ff_503 <= io_i_mux_bus_503;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_504 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_504 <= 1'h0;
    end else begin
      r_mux_bus_ff_504 <= io_i_mux_bus_504;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_505 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_505 <= 1'h0;
    end else begin
      r_mux_bus_ff_505 <= io_i_mux_bus_505;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_506 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_506 <= 1'h0;
    end else begin
      r_mux_bus_ff_506 <= io_i_mux_bus_506;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_507 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_507 <= 1'h0;
    end else begin
      r_mux_bus_ff_507 <= io_i_mux_bus_507;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_508 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_508 <= 1'h0;
    end else begin
      r_mux_bus_ff_508 <= io_i_mux_bus_508;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_509 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_509 <= 1'h0;
    end else begin
      r_mux_bus_ff_509 <= io_i_mux_bus_509;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_510 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_510 <= 1'h0;
    end else begin
      r_mux_bus_ff_510 <= io_i_mux_bus_510;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_511 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_511 <= 1'h0;
    end else begin
      r_mux_bus_ff_511 <= io_i_mux_bus_511;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_512 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_512 <= 1'h0;
    end else begin
      r_mux_bus_ff_512 <= io_i_mux_bus_512;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_513 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_513 <= 1'h0;
    end else begin
      r_mux_bus_ff_513 <= io_i_mux_bus_513;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_514 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_514 <= 1'h0;
    end else begin
      r_mux_bus_ff_514 <= io_i_mux_bus_514;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_515 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_515 <= 1'h0;
    end else begin
      r_mux_bus_ff_515 <= io_i_mux_bus_515;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_516 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_516 <= 1'h0;
    end else begin
      r_mux_bus_ff_516 <= io_i_mux_bus_516;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_517 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_517 <= 1'h0;
    end else begin
      r_mux_bus_ff_517 <= io_i_mux_bus_517;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_518 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_518 <= 1'h0;
    end else begin
      r_mux_bus_ff_518 <= io_i_mux_bus_518;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_519 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_519 <= 1'h0;
    end else begin
      r_mux_bus_ff_519 <= io_i_mux_bus_519;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_520 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_520 <= 1'h0;
    end else begin
      r_mux_bus_ff_520 <= io_i_mux_bus_520;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_521 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_521 <= 1'h0;
    end else begin
      r_mux_bus_ff_521 <= io_i_mux_bus_521;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_522 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_522 <= 1'h0;
    end else begin
      r_mux_bus_ff_522 <= io_i_mux_bus_522;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_523 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_523 <= 1'h0;
    end else begin
      r_mux_bus_ff_523 <= io_i_mux_bus_523;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_524 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_524 <= 1'h0;
    end else begin
      r_mux_bus_ff_524 <= io_i_mux_bus_524;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_525 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_525 <= 1'h0;
    end else begin
      r_mux_bus_ff_525 <= io_i_mux_bus_525;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_526 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_526 <= 1'h0;
    end else begin
      r_mux_bus_ff_526 <= io_i_mux_bus_526;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_527 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_527 <= 1'h0;
    end else begin
      r_mux_bus_ff_527 <= io_i_mux_bus_527;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_528 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_528 <= 1'h0;
    end else begin
      r_mux_bus_ff_528 <= io_i_mux_bus_528;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_529 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_529 <= 1'h0;
    end else begin
      r_mux_bus_ff_529 <= io_i_mux_bus_529;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_530 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_530 <= 1'h0;
    end else begin
      r_mux_bus_ff_530 <= io_i_mux_bus_530;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_531 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_531 <= 1'h0;
    end else begin
      r_mux_bus_ff_531 <= io_i_mux_bus_531;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_532 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_532 <= 1'h0;
    end else begin
      r_mux_bus_ff_532 <= io_i_mux_bus_532;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_533 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_533 <= 1'h0;
    end else begin
      r_mux_bus_ff_533 <= io_i_mux_bus_533;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_534 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_534 <= 1'h0;
    end else begin
      r_mux_bus_ff_534 <= io_i_mux_bus_534;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_535 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_535 <= 1'h0;
    end else begin
      r_mux_bus_ff_535 <= io_i_mux_bus_535;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_536 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_536 <= 1'h0;
    end else begin
      r_mux_bus_ff_536 <= io_i_mux_bus_536;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_537 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_537 <= 1'h0;
    end else begin
      r_mux_bus_ff_537 <= io_i_mux_bus_537;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_538 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_538 <= 1'h0;
    end else begin
      r_mux_bus_ff_538 <= io_i_mux_bus_538;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_539 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_539 <= 1'h0;
    end else begin
      r_mux_bus_ff_539 <= io_i_mux_bus_539;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_540 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_540 <= 1'h0;
    end else begin
      r_mux_bus_ff_540 <= io_i_mux_bus_540;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_541 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_541 <= 1'h0;
    end else begin
      r_mux_bus_ff_541 <= io_i_mux_bus_541;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_542 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_542 <= 1'h0;
    end else begin
      r_mux_bus_ff_542 <= io_i_mux_bus_542;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_543 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_543 <= 1'h0;
    end else begin
      r_mux_bus_ff_543 <= io_i_mux_bus_543;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_544 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_544 <= 1'h0;
    end else begin
      r_mux_bus_ff_544 <= io_i_mux_bus_544;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_545 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_545 <= 1'h0;
    end else begin
      r_mux_bus_ff_545 <= io_i_mux_bus_545;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_546 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_546 <= 1'h0;
    end else begin
      r_mux_bus_ff_546 <= io_i_mux_bus_546;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_547 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_547 <= 1'h0;
    end else begin
      r_mux_bus_ff_547 <= io_i_mux_bus_547;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_548 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_548 <= 1'h0;
    end else begin
      r_mux_bus_ff_548 <= io_i_mux_bus_548;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_549 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_549 <= 1'h0;
    end else begin
      r_mux_bus_ff_549 <= io_i_mux_bus_549;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_550 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_550 <= 1'h0;
    end else begin
      r_mux_bus_ff_550 <= io_i_mux_bus_550;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_551 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_551 <= 1'h0;
    end else begin
      r_mux_bus_ff_551 <= io_i_mux_bus_551;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_552 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_552 <= 1'h0;
    end else begin
      r_mux_bus_ff_552 <= io_i_mux_bus_552;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_553 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_553 <= 1'h0;
    end else begin
      r_mux_bus_ff_553 <= io_i_mux_bus_553;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_554 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_554 <= 1'h0;
    end else begin
      r_mux_bus_ff_554 <= io_i_mux_bus_554;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_555 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_555 <= 1'h0;
    end else begin
      r_mux_bus_ff_555 <= io_i_mux_bus_555;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_556 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_556 <= 1'h0;
    end else begin
      r_mux_bus_ff_556 <= io_i_mux_bus_556;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_557 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_557 <= 1'h0;
    end else begin
      r_mux_bus_ff_557 <= io_i_mux_bus_557;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_558 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_558 <= 1'h0;
    end else begin
      r_mux_bus_ff_558 <= io_i_mux_bus_558;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_559 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_559 <= 1'h0;
    end else begin
      r_mux_bus_ff_559 <= io_i_mux_bus_559;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_560 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_560 <= 1'h0;
    end else begin
      r_mux_bus_ff_560 <= io_i_mux_bus_560;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_561 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_561 <= 1'h0;
    end else begin
      r_mux_bus_ff_561 <= io_i_mux_bus_561;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_562 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_562 <= 1'h0;
    end else begin
      r_mux_bus_ff_562 <= io_i_mux_bus_562;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_563 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_563 <= 1'h0;
    end else begin
      r_mux_bus_ff_563 <= io_i_mux_bus_563;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_564 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_564 <= 1'h0;
    end else begin
      r_mux_bus_ff_564 <= io_i_mux_bus_564;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_565 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_565 <= 1'h0;
    end else begin
      r_mux_bus_ff_565 <= io_i_mux_bus_565;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_566 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_566 <= 1'h0;
    end else begin
      r_mux_bus_ff_566 <= io_i_mux_bus_566;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_567 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_567 <= 1'h0;
    end else begin
      r_mux_bus_ff_567 <= io_i_mux_bus_567;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_568 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_568 <= 1'h0;
    end else begin
      r_mux_bus_ff_568 <= io_i_mux_bus_568;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_569 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_569 <= 1'h0;
    end else begin
      r_mux_bus_ff_569 <= io_i_mux_bus_569;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_570 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_570 <= 1'h0;
    end else begin
      r_mux_bus_ff_570 <= io_i_mux_bus_570;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_571 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_571 <= 1'h0;
    end else begin
      r_mux_bus_ff_571 <= io_i_mux_bus_571;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_572 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_572 <= 1'h0;
    end else begin
      r_mux_bus_ff_572 <= io_i_mux_bus_572;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_573 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_573 <= 1'h0;
    end else begin
      r_mux_bus_ff_573 <= io_i_mux_bus_573;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_574 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_574 <= 1'h0;
    end else begin
      r_mux_bus_ff_574 <= io_i_mux_bus_574;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_575 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_575 <= 1'h0;
    end else begin
      r_mux_bus_ff_575 <= io_i_mux_bus_575;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_576 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_576 <= 1'h0;
    end else begin
      r_mux_bus_ff_576 <= io_i_mux_bus_576;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_577 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_577 <= 1'h0;
    end else begin
      r_mux_bus_ff_577 <= io_i_mux_bus_577;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_578 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_578 <= 1'h0;
    end else begin
      r_mux_bus_ff_578 <= io_i_mux_bus_578;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_579 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_579 <= 1'h0;
    end else begin
      r_mux_bus_ff_579 <= io_i_mux_bus_579;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_580 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_580 <= 1'h0;
    end else begin
      r_mux_bus_ff_580 <= io_i_mux_bus_580;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_581 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_581 <= 1'h0;
    end else begin
      r_mux_bus_ff_581 <= io_i_mux_bus_581;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_582 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_582 <= 1'h0;
    end else begin
      r_mux_bus_ff_582 <= io_i_mux_bus_582;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_583 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_583 <= 1'h0;
    end else begin
      r_mux_bus_ff_583 <= io_i_mux_bus_583;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_584 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_584 <= 1'h0;
    end else begin
      r_mux_bus_ff_584 <= io_i_mux_bus_584;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_585 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_585 <= 1'h0;
    end else begin
      r_mux_bus_ff_585 <= io_i_mux_bus_585;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_586 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_586 <= 1'h0;
    end else begin
      r_mux_bus_ff_586 <= io_i_mux_bus_586;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_587 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_587 <= 1'h0;
    end else begin
      r_mux_bus_ff_587 <= io_i_mux_bus_587;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_588 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_588 <= 1'h0;
    end else begin
      r_mux_bus_ff_588 <= io_i_mux_bus_588;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_589 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_589 <= 1'h0;
    end else begin
      r_mux_bus_ff_589 <= io_i_mux_bus_589;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_590 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_590 <= 1'h0;
    end else begin
      r_mux_bus_ff_590 <= io_i_mux_bus_590;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_591 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_591 <= 1'h0;
    end else begin
      r_mux_bus_ff_591 <= io_i_mux_bus_591;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_592 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_592 <= 1'h0;
    end else begin
      r_mux_bus_ff_592 <= io_i_mux_bus_592;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_593 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_593 <= 1'h0;
    end else begin
      r_mux_bus_ff_593 <= io_i_mux_bus_593;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_594 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_594 <= 1'h0;
    end else begin
      r_mux_bus_ff_594 <= io_i_mux_bus_594;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_595 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_595 <= 1'h0;
    end else begin
      r_mux_bus_ff_595 <= io_i_mux_bus_595;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_596 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_596 <= 1'h0;
    end else begin
      r_mux_bus_ff_596 <= io_i_mux_bus_596;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_597 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_597 <= 1'h0;
    end else begin
      r_mux_bus_ff_597 <= io_i_mux_bus_597;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_598 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_598 <= 1'h0;
    end else begin
      r_mux_bus_ff_598 <= io_i_mux_bus_598;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_599 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_599 <= 1'h0;
    end else begin
      r_mux_bus_ff_599 <= io_i_mux_bus_599;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_600 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_600 <= 1'h0;
    end else begin
      r_mux_bus_ff_600 <= io_i_mux_bus_600;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_601 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_601 <= 1'h0;
    end else begin
      r_mux_bus_ff_601 <= io_i_mux_bus_601;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_602 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_602 <= 1'h0;
    end else begin
      r_mux_bus_ff_602 <= io_i_mux_bus_602;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_603 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_603 <= 1'h0;
    end else begin
      r_mux_bus_ff_603 <= io_i_mux_bus_603;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_604 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_604 <= 1'h0;
    end else begin
      r_mux_bus_ff_604 <= io_i_mux_bus_604;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_605 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_605 <= 1'h0;
    end else begin
      r_mux_bus_ff_605 <= io_i_mux_bus_605;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_606 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_606 <= 1'h0;
    end else begin
      r_mux_bus_ff_606 <= io_i_mux_bus_606;
    end
    if (reset) begin // @[Benes.scala 77:32]
      r_mux_bus_ff_607 <= 1'h0; // @[Benes.scala 77:32]
    end else if (reset) begin // @[Benes.scala 84:23]
      r_mux_bus_ff_607 <= 1'h0;
    end else begin
      r_mux_bus_ff_607 <= io_i_mux_bus_607;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_data_bus_ff_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  r_data_bus_ff_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  r_data_bus_ff_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  r_data_bus_ff_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  r_data_bus_ff_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  r_data_bus_ff_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  r_data_bus_ff_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  r_data_bus_ff_7 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  r_data_bus_ff_8 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  r_data_bus_ff_9 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  r_data_bus_ff_10 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  r_data_bus_ff_11 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  r_data_bus_ff_12 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  r_data_bus_ff_13 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  r_data_bus_ff_14 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  r_data_bus_ff_15 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  r_data_bus_ff_16 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  r_data_bus_ff_17 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  r_data_bus_ff_18 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  r_data_bus_ff_19 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  r_data_bus_ff_20 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  r_data_bus_ff_21 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  r_data_bus_ff_22 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  r_data_bus_ff_23 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  r_data_bus_ff_24 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  r_data_bus_ff_25 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  r_data_bus_ff_26 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  r_data_bus_ff_27 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  r_data_bus_ff_28 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  r_data_bus_ff_29 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  r_data_bus_ff_30 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  r_data_bus_ff_31 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  r_mux_bus_ff_0 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  r_mux_bus_ff_1 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  r_mux_bus_ff_2 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  r_mux_bus_ff_3 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  r_mux_bus_ff_4 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  r_mux_bus_ff_5 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  r_mux_bus_ff_6 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  r_mux_bus_ff_7 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  r_mux_bus_ff_8 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  r_mux_bus_ff_9 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  r_mux_bus_ff_10 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  r_mux_bus_ff_11 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  r_mux_bus_ff_12 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  r_mux_bus_ff_13 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  r_mux_bus_ff_14 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  r_mux_bus_ff_15 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  r_mux_bus_ff_16 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  r_mux_bus_ff_17 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  r_mux_bus_ff_18 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  r_mux_bus_ff_19 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  r_mux_bus_ff_20 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  r_mux_bus_ff_21 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  r_mux_bus_ff_22 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  r_mux_bus_ff_23 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  r_mux_bus_ff_24 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  r_mux_bus_ff_25 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  r_mux_bus_ff_26 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  r_mux_bus_ff_27 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  r_mux_bus_ff_28 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  r_mux_bus_ff_29 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  r_mux_bus_ff_30 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  r_mux_bus_ff_31 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  r_mux_bus_ff_32 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  r_mux_bus_ff_33 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  r_mux_bus_ff_34 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  r_mux_bus_ff_35 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  r_mux_bus_ff_36 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  r_mux_bus_ff_37 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  r_mux_bus_ff_38 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  r_mux_bus_ff_39 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  r_mux_bus_ff_40 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  r_mux_bus_ff_41 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  r_mux_bus_ff_42 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  r_mux_bus_ff_43 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  r_mux_bus_ff_44 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  r_mux_bus_ff_45 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  r_mux_bus_ff_46 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  r_mux_bus_ff_47 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  r_mux_bus_ff_48 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  r_mux_bus_ff_49 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  r_mux_bus_ff_50 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  r_mux_bus_ff_51 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  r_mux_bus_ff_52 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  r_mux_bus_ff_53 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  r_mux_bus_ff_54 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  r_mux_bus_ff_55 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  r_mux_bus_ff_56 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  r_mux_bus_ff_57 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  r_mux_bus_ff_58 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  r_mux_bus_ff_59 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  r_mux_bus_ff_60 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  r_mux_bus_ff_61 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  r_mux_bus_ff_62 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  r_mux_bus_ff_63 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  r_mux_bus_ff_64 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  r_mux_bus_ff_65 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  r_mux_bus_ff_66 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  r_mux_bus_ff_67 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  r_mux_bus_ff_68 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  r_mux_bus_ff_69 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  r_mux_bus_ff_70 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  r_mux_bus_ff_71 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  r_mux_bus_ff_72 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  r_mux_bus_ff_73 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  r_mux_bus_ff_74 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  r_mux_bus_ff_75 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  r_mux_bus_ff_76 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  r_mux_bus_ff_77 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  r_mux_bus_ff_78 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  r_mux_bus_ff_79 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  r_mux_bus_ff_80 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  r_mux_bus_ff_81 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  r_mux_bus_ff_82 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  r_mux_bus_ff_83 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  r_mux_bus_ff_84 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  r_mux_bus_ff_85 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  r_mux_bus_ff_86 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  r_mux_bus_ff_87 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  r_mux_bus_ff_88 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  r_mux_bus_ff_89 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  r_mux_bus_ff_90 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  r_mux_bus_ff_91 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  r_mux_bus_ff_92 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  r_mux_bus_ff_93 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  r_mux_bus_ff_94 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  r_mux_bus_ff_95 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  r_mux_bus_ff_96 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  r_mux_bus_ff_97 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  r_mux_bus_ff_98 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  r_mux_bus_ff_99 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  r_mux_bus_ff_100 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  r_mux_bus_ff_101 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  r_mux_bus_ff_102 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  r_mux_bus_ff_103 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  r_mux_bus_ff_104 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  r_mux_bus_ff_105 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  r_mux_bus_ff_106 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  r_mux_bus_ff_107 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  r_mux_bus_ff_108 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  r_mux_bus_ff_109 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  r_mux_bus_ff_110 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  r_mux_bus_ff_111 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  r_mux_bus_ff_112 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  r_mux_bus_ff_113 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  r_mux_bus_ff_114 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  r_mux_bus_ff_115 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  r_mux_bus_ff_116 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  r_mux_bus_ff_117 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  r_mux_bus_ff_118 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  r_mux_bus_ff_119 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  r_mux_bus_ff_120 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  r_mux_bus_ff_121 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  r_mux_bus_ff_122 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  r_mux_bus_ff_123 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  r_mux_bus_ff_124 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  r_mux_bus_ff_125 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  r_mux_bus_ff_126 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  r_mux_bus_ff_127 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  r_mux_bus_ff_128 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  r_mux_bus_ff_129 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  r_mux_bus_ff_130 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  r_mux_bus_ff_131 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  r_mux_bus_ff_132 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  r_mux_bus_ff_133 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  r_mux_bus_ff_134 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  r_mux_bus_ff_135 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  r_mux_bus_ff_136 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  r_mux_bus_ff_137 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  r_mux_bus_ff_138 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  r_mux_bus_ff_139 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  r_mux_bus_ff_140 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  r_mux_bus_ff_141 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  r_mux_bus_ff_142 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  r_mux_bus_ff_143 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  r_mux_bus_ff_144 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  r_mux_bus_ff_145 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  r_mux_bus_ff_146 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  r_mux_bus_ff_147 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  r_mux_bus_ff_148 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  r_mux_bus_ff_149 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  r_mux_bus_ff_150 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  r_mux_bus_ff_151 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  r_mux_bus_ff_152 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  r_mux_bus_ff_153 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  r_mux_bus_ff_154 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  r_mux_bus_ff_155 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  r_mux_bus_ff_156 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  r_mux_bus_ff_157 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  r_mux_bus_ff_158 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  r_mux_bus_ff_159 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  r_mux_bus_ff_160 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  r_mux_bus_ff_161 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  r_mux_bus_ff_162 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  r_mux_bus_ff_163 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  r_mux_bus_ff_164 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  r_mux_bus_ff_165 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  r_mux_bus_ff_166 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  r_mux_bus_ff_167 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  r_mux_bus_ff_168 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  r_mux_bus_ff_169 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  r_mux_bus_ff_170 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  r_mux_bus_ff_171 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  r_mux_bus_ff_172 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  r_mux_bus_ff_173 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  r_mux_bus_ff_174 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  r_mux_bus_ff_175 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  r_mux_bus_ff_176 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  r_mux_bus_ff_177 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  r_mux_bus_ff_178 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  r_mux_bus_ff_179 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  r_mux_bus_ff_180 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  r_mux_bus_ff_181 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  r_mux_bus_ff_182 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  r_mux_bus_ff_183 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  r_mux_bus_ff_184 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  r_mux_bus_ff_185 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  r_mux_bus_ff_186 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  r_mux_bus_ff_187 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  r_mux_bus_ff_188 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  r_mux_bus_ff_189 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  r_mux_bus_ff_190 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  r_mux_bus_ff_191 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  r_mux_bus_ff_192 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  r_mux_bus_ff_193 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  r_mux_bus_ff_194 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  r_mux_bus_ff_195 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  r_mux_bus_ff_196 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  r_mux_bus_ff_197 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  r_mux_bus_ff_198 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  r_mux_bus_ff_199 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  r_mux_bus_ff_200 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  r_mux_bus_ff_201 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  r_mux_bus_ff_202 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  r_mux_bus_ff_203 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  r_mux_bus_ff_204 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  r_mux_bus_ff_205 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  r_mux_bus_ff_206 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  r_mux_bus_ff_207 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  r_mux_bus_ff_208 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  r_mux_bus_ff_209 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  r_mux_bus_ff_210 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  r_mux_bus_ff_211 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  r_mux_bus_ff_212 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  r_mux_bus_ff_213 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  r_mux_bus_ff_214 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  r_mux_bus_ff_215 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  r_mux_bus_ff_216 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  r_mux_bus_ff_217 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  r_mux_bus_ff_218 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  r_mux_bus_ff_219 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  r_mux_bus_ff_220 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  r_mux_bus_ff_221 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  r_mux_bus_ff_222 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  r_mux_bus_ff_223 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  r_mux_bus_ff_224 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  r_mux_bus_ff_225 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  r_mux_bus_ff_226 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  r_mux_bus_ff_227 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  r_mux_bus_ff_228 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  r_mux_bus_ff_229 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  r_mux_bus_ff_230 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  r_mux_bus_ff_231 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  r_mux_bus_ff_232 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  r_mux_bus_ff_233 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  r_mux_bus_ff_234 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  r_mux_bus_ff_235 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  r_mux_bus_ff_236 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  r_mux_bus_ff_237 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  r_mux_bus_ff_238 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  r_mux_bus_ff_239 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  r_mux_bus_ff_240 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  r_mux_bus_ff_241 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  r_mux_bus_ff_242 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  r_mux_bus_ff_243 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  r_mux_bus_ff_244 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  r_mux_bus_ff_245 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  r_mux_bus_ff_246 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  r_mux_bus_ff_247 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  r_mux_bus_ff_248 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  r_mux_bus_ff_249 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  r_mux_bus_ff_250 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  r_mux_bus_ff_251 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  r_mux_bus_ff_252 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  r_mux_bus_ff_253 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  r_mux_bus_ff_254 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  r_mux_bus_ff_255 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  r_mux_bus_ff_256 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  r_mux_bus_ff_257 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  r_mux_bus_ff_258 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  r_mux_bus_ff_259 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  r_mux_bus_ff_260 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  r_mux_bus_ff_261 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  r_mux_bus_ff_262 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  r_mux_bus_ff_263 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  r_mux_bus_ff_264 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  r_mux_bus_ff_265 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  r_mux_bus_ff_266 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  r_mux_bus_ff_267 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  r_mux_bus_ff_268 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  r_mux_bus_ff_269 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  r_mux_bus_ff_270 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  r_mux_bus_ff_271 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  r_mux_bus_ff_272 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  r_mux_bus_ff_273 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  r_mux_bus_ff_274 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  r_mux_bus_ff_275 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  r_mux_bus_ff_276 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  r_mux_bus_ff_277 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  r_mux_bus_ff_278 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  r_mux_bus_ff_279 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  r_mux_bus_ff_280 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  r_mux_bus_ff_281 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  r_mux_bus_ff_282 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  r_mux_bus_ff_283 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  r_mux_bus_ff_284 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  r_mux_bus_ff_285 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  r_mux_bus_ff_286 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  r_mux_bus_ff_287 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  r_mux_bus_ff_288 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  r_mux_bus_ff_289 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  r_mux_bus_ff_290 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  r_mux_bus_ff_291 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  r_mux_bus_ff_292 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  r_mux_bus_ff_293 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  r_mux_bus_ff_294 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  r_mux_bus_ff_295 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  r_mux_bus_ff_296 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  r_mux_bus_ff_297 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  r_mux_bus_ff_298 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  r_mux_bus_ff_299 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  r_mux_bus_ff_300 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  r_mux_bus_ff_301 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  r_mux_bus_ff_302 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  r_mux_bus_ff_303 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  r_mux_bus_ff_304 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  r_mux_bus_ff_305 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  r_mux_bus_ff_306 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  r_mux_bus_ff_307 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  r_mux_bus_ff_308 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  r_mux_bus_ff_309 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  r_mux_bus_ff_310 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  r_mux_bus_ff_311 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  r_mux_bus_ff_312 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  r_mux_bus_ff_313 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  r_mux_bus_ff_314 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  r_mux_bus_ff_315 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  r_mux_bus_ff_316 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  r_mux_bus_ff_317 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  r_mux_bus_ff_318 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  r_mux_bus_ff_319 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  r_mux_bus_ff_320 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  r_mux_bus_ff_321 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  r_mux_bus_ff_322 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  r_mux_bus_ff_323 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  r_mux_bus_ff_324 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  r_mux_bus_ff_325 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  r_mux_bus_ff_326 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  r_mux_bus_ff_327 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  r_mux_bus_ff_328 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  r_mux_bus_ff_329 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  r_mux_bus_ff_330 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  r_mux_bus_ff_331 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  r_mux_bus_ff_332 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  r_mux_bus_ff_333 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  r_mux_bus_ff_334 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  r_mux_bus_ff_335 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  r_mux_bus_ff_336 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  r_mux_bus_ff_337 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  r_mux_bus_ff_338 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  r_mux_bus_ff_339 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  r_mux_bus_ff_340 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  r_mux_bus_ff_341 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  r_mux_bus_ff_342 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  r_mux_bus_ff_343 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  r_mux_bus_ff_344 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  r_mux_bus_ff_345 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  r_mux_bus_ff_346 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  r_mux_bus_ff_347 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  r_mux_bus_ff_348 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  r_mux_bus_ff_349 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  r_mux_bus_ff_350 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  r_mux_bus_ff_351 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  r_mux_bus_ff_352 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  r_mux_bus_ff_353 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  r_mux_bus_ff_354 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  r_mux_bus_ff_355 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  r_mux_bus_ff_356 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  r_mux_bus_ff_357 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  r_mux_bus_ff_358 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  r_mux_bus_ff_359 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  r_mux_bus_ff_360 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  r_mux_bus_ff_361 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  r_mux_bus_ff_362 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  r_mux_bus_ff_363 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  r_mux_bus_ff_364 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  r_mux_bus_ff_365 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  r_mux_bus_ff_366 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  r_mux_bus_ff_367 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  r_mux_bus_ff_368 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  r_mux_bus_ff_369 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  r_mux_bus_ff_370 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  r_mux_bus_ff_371 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  r_mux_bus_ff_372 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  r_mux_bus_ff_373 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  r_mux_bus_ff_374 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  r_mux_bus_ff_375 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  r_mux_bus_ff_376 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  r_mux_bus_ff_377 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  r_mux_bus_ff_378 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  r_mux_bus_ff_379 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  r_mux_bus_ff_380 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  r_mux_bus_ff_381 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  r_mux_bus_ff_382 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  r_mux_bus_ff_383 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  r_mux_bus_ff_384 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  r_mux_bus_ff_385 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  r_mux_bus_ff_386 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  r_mux_bus_ff_387 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  r_mux_bus_ff_388 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  r_mux_bus_ff_389 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  r_mux_bus_ff_390 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  r_mux_bus_ff_391 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  r_mux_bus_ff_392 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  r_mux_bus_ff_393 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  r_mux_bus_ff_394 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  r_mux_bus_ff_395 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  r_mux_bus_ff_396 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  r_mux_bus_ff_397 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  r_mux_bus_ff_398 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  r_mux_bus_ff_399 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  r_mux_bus_ff_400 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  r_mux_bus_ff_401 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  r_mux_bus_ff_402 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  r_mux_bus_ff_403 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  r_mux_bus_ff_404 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  r_mux_bus_ff_405 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  r_mux_bus_ff_406 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  r_mux_bus_ff_407 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  r_mux_bus_ff_408 = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  r_mux_bus_ff_409 = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  r_mux_bus_ff_410 = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  r_mux_bus_ff_411 = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  r_mux_bus_ff_412 = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  r_mux_bus_ff_413 = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  r_mux_bus_ff_414 = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  r_mux_bus_ff_415 = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  r_mux_bus_ff_416 = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  r_mux_bus_ff_417 = _RAND_449[0:0];
  _RAND_450 = {1{`RANDOM}};
  r_mux_bus_ff_418 = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  r_mux_bus_ff_419 = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  r_mux_bus_ff_420 = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  r_mux_bus_ff_421 = _RAND_453[0:0];
  _RAND_454 = {1{`RANDOM}};
  r_mux_bus_ff_422 = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  r_mux_bus_ff_423 = _RAND_455[0:0];
  _RAND_456 = {1{`RANDOM}};
  r_mux_bus_ff_424 = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  r_mux_bus_ff_425 = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  r_mux_bus_ff_426 = _RAND_458[0:0];
  _RAND_459 = {1{`RANDOM}};
  r_mux_bus_ff_427 = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  r_mux_bus_ff_428 = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  r_mux_bus_ff_429 = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  r_mux_bus_ff_430 = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  r_mux_bus_ff_431 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  r_mux_bus_ff_432 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  r_mux_bus_ff_433 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  r_mux_bus_ff_434 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  r_mux_bus_ff_435 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  r_mux_bus_ff_436 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  r_mux_bus_ff_437 = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  r_mux_bus_ff_438 = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  r_mux_bus_ff_439 = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  r_mux_bus_ff_440 = _RAND_472[0:0];
  _RAND_473 = {1{`RANDOM}};
  r_mux_bus_ff_441 = _RAND_473[0:0];
  _RAND_474 = {1{`RANDOM}};
  r_mux_bus_ff_442 = _RAND_474[0:0];
  _RAND_475 = {1{`RANDOM}};
  r_mux_bus_ff_443 = _RAND_475[0:0];
  _RAND_476 = {1{`RANDOM}};
  r_mux_bus_ff_444 = _RAND_476[0:0];
  _RAND_477 = {1{`RANDOM}};
  r_mux_bus_ff_445 = _RAND_477[0:0];
  _RAND_478 = {1{`RANDOM}};
  r_mux_bus_ff_446 = _RAND_478[0:0];
  _RAND_479 = {1{`RANDOM}};
  r_mux_bus_ff_447 = _RAND_479[0:0];
  _RAND_480 = {1{`RANDOM}};
  r_mux_bus_ff_448 = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  r_mux_bus_ff_449 = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  r_mux_bus_ff_450 = _RAND_482[0:0];
  _RAND_483 = {1{`RANDOM}};
  r_mux_bus_ff_451 = _RAND_483[0:0];
  _RAND_484 = {1{`RANDOM}};
  r_mux_bus_ff_452 = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  r_mux_bus_ff_453 = _RAND_485[0:0];
  _RAND_486 = {1{`RANDOM}};
  r_mux_bus_ff_454 = _RAND_486[0:0];
  _RAND_487 = {1{`RANDOM}};
  r_mux_bus_ff_455 = _RAND_487[0:0];
  _RAND_488 = {1{`RANDOM}};
  r_mux_bus_ff_456 = _RAND_488[0:0];
  _RAND_489 = {1{`RANDOM}};
  r_mux_bus_ff_457 = _RAND_489[0:0];
  _RAND_490 = {1{`RANDOM}};
  r_mux_bus_ff_458 = _RAND_490[0:0];
  _RAND_491 = {1{`RANDOM}};
  r_mux_bus_ff_459 = _RAND_491[0:0];
  _RAND_492 = {1{`RANDOM}};
  r_mux_bus_ff_460 = _RAND_492[0:0];
  _RAND_493 = {1{`RANDOM}};
  r_mux_bus_ff_461 = _RAND_493[0:0];
  _RAND_494 = {1{`RANDOM}};
  r_mux_bus_ff_462 = _RAND_494[0:0];
  _RAND_495 = {1{`RANDOM}};
  r_mux_bus_ff_463 = _RAND_495[0:0];
  _RAND_496 = {1{`RANDOM}};
  r_mux_bus_ff_464 = _RAND_496[0:0];
  _RAND_497 = {1{`RANDOM}};
  r_mux_bus_ff_465 = _RAND_497[0:0];
  _RAND_498 = {1{`RANDOM}};
  r_mux_bus_ff_466 = _RAND_498[0:0];
  _RAND_499 = {1{`RANDOM}};
  r_mux_bus_ff_467 = _RAND_499[0:0];
  _RAND_500 = {1{`RANDOM}};
  r_mux_bus_ff_468 = _RAND_500[0:0];
  _RAND_501 = {1{`RANDOM}};
  r_mux_bus_ff_469 = _RAND_501[0:0];
  _RAND_502 = {1{`RANDOM}};
  r_mux_bus_ff_470 = _RAND_502[0:0];
  _RAND_503 = {1{`RANDOM}};
  r_mux_bus_ff_471 = _RAND_503[0:0];
  _RAND_504 = {1{`RANDOM}};
  r_mux_bus_ff_472 = _RAND_504[0:0];
  _RAND_505 = {1{`RANDOM}};
  r_mux_bus_ff_473 = _RAND_505[0:0];
  _RAND_506 = {1{`RANDOM}};
  r_mux_bus_ff_474 = _RAND_506[0:0];
  _RAND_507 = {1{`RANDOM}};
  r_mux_bus_ff_475 = _RAND_507[0:0];
  _RAND_508 = {1{`RANDOM}};
  r_mux_bus_ff_476 = _RAND_508[0:0];
  _RAND_509 = {1{`RANDOM}};
  r_mux_bus_ff_477 = _RAND_509[0:0];
  _RAND_510 = {1{`RANDOM}};
  r_mux_bus_ff_478 = _RAND_510[0:0];
  _RAND_511 = {1{`RANDOM}};
  r_mux_bus_ff_479 = _RAND_511[0:0];
  _RAND_512 = {1{`RANDOM}};
  r_mux_bus_ff_480 = _RAND_512[0:0];
  _RAND_513 = {1{`RANDOM}};
  r_mux_bus_ff_481 = _RAND_513[0:0];
  _RAND_514 = {1{`RANDOM}};
  r_mux_bus_ff_482 = _RAND_514[0:0];
  _RAND_515 = {1{`RANDOM}};
  r_mux_bus_ff_483 = _RAND_515[0:0];
  _RAND_516 = {1{`RANDOM}};
  r_mux_bus_ff_484 = _RAND_516[0:0];
  _RAND_517 = {1{`RANDOM}};
  r_mux_bus_ff_485 = _RAND_517[0:0];
  _RAND_518 = {1{`RANDOM}};
  r_mux_bus_ff_486 = _RAND_518[0:0];
  _RAND_519 = {1{`RANDOM}};
  r_mux_bus_ff_487 = _RAND_519[0:0];
  _RAND_520 = {1{`RANDOM}};
  r_mux_bus_ff_488 = _RAND_520[0:0];
  _RAND_521 = {1{`RANDOM}};
  r_mux_bus_ff_489 = _RAND_521[0:0];
  _RAND_522 = {1{`RANDOM}};
  r_mux_bus_ff_490 = _RAND_522[0:0];
  _RAND_523 = {1{`RANDOM}};
  r_mux_bus_ff_491 = _RAND_523[0:0];
  _RAND_524 = {1{`RANDOM}};
  r_mux_bus_ff_492 = _RAND_524[0:0];
  _RAND_525 = {1{`RANDOM}};
  r_mux_bus_ff_493 = _RAND_525[0:0];
  _RAND_526 = {1{`RANDOM}};
  r_mux_bus_ff_494 = _RAND_526[0:0];
  _RAND_527 = {1{`RANDOM}};
  r_mux_bus_ff_495 = _RAND_527[0:0];
  _RAND_528 = {1{`RANDOM}};
  r_mux_bus_ff_496 = _RAND_528[0:0];
  _RAND_529 = {1{`RANDOM}};
  r_mux_bus_ff_497 = _RAND_529[0:0];
  _RAND_530 = {1{`RANDOM}};
  r_mux_bus_ff_498 = _RAND_530[0:0];
  _RAND_531 = {1{`RANDOM}};
  r_mux_bus_ff_499 = _RAND_531[0:0];
  _RAND_532 = {1{`RANDOM}};
  r_mux_bus_ff_500 = _RAND_532[0:0];
  _RAND_533 = {1{`RANDOM}};
  r_mux_bus_ff_501 = _RAND_533[0:0];
  _RAND_534 = {1{`RANDOM}};
  r_mux_bus_ff_502 = _RAND_534[0:0];
  _RAND_535 = {1{`RANDOM}};
  r_mux_bus_ff_503 = _RAND_535[0:0];
  _RAND_536 = {1{`RANDOM}};
  r_mux_bus_ff_504 = _RAND_536[0:0];
  _RAND_537 = {1{`RANDOM}};
  r_mux_bus_ff_505 = _RAND_537[0:0];
  _RAND_538 = {1{`RANDOM}};
  r_mux_bus_ff_506 = _RAND_538[0:0];
  _RAND_539 = {1{`RANDOM}};
  r_mux_bus_ff_507 = _RAND_539[0:0];
  _RAND_540 = {1{`RANDOM}};
  r_mux_bus_ff_508 = _RAND_540[0:0];
  _RAND_541 = {1{`RANDOM}};
  r_mux_bus_ff_509 = _RAND_541[0:0];
  _RAND_542 = {1{`RANDOM}};
  r_mux_bus_ff_510 = _RAND_542[0:0];
  _RAND_543 = {1{`RANDOM}};
  r_mux_bus_ff_511 = _RAND_543[0:0];
  _RAND_544 = {1{`RANDOM}};
  r_mux_bus_ff_512 = _RAND_544[0:0];
  _RAND_545 = {1{`RANDOM}};
  r_mux_bus_ff_513 = _RAND_545[0:0];
  _RAND_546 = {1{`RANDOM}};
  r_mux_bus_ff_514 = _RAND_546[0:0];
  _RAND_547 = {1{`RANDOM}};
  r_mux_bus_ff_515 = _RAND_547[0:0];
  _RAND_548 = {1{`RANDOM}};
  r_mux_bus_ff_516 = _RAND_548[0:0];
  _RAND_549 = {1{`RANDOM}};
  r_mux_bus_ff_517 = _RAND_549[0:0];
  _RAND_550 = {1{`RANDOM}};
  r_mux_bus_ff_518 = _RAND_550[0:0];
  _RAND_551 = {1{`RANDOM}};
  r_mux_bus_ff_519 = _RAND_551[0:0];
  _RAND_552 = {1{`RANDOM}};
  r_mux_bus_ff_520 = _RAND_552[0:0];
  _RAND_553 = {1{`RANDOM}};
  r_mux_bus_ff_521 = _RAND_553[0:0];
  _RAND_554 = {1{`RANDOM}};
  r_mux_bus_ff_522 = _RAND_554[0:0];
  _RAND_555 = {1{`RANDOM}};
  r_mux_bus_ff_523 = _RAND_555[0:0];
  _RAND_556 = {1{`RANDOM}};
  r_mux_bus_ff_524 = _RAND_556[0:0];
  _RAND_557 = {1{`RANDOM}};
  r_mux_bus_ff_525 = _RAND_557[0:0];
  _RAND_558 = {1{`RANDOM}};
  r_mux_bus_ff_526 = _RAND_558[0:0];
  _RAND_559 = {1{`RANDOM}};
  r_mux_bus_ff_527 = _RAND_559[0:0];
  _RAND_560 = {1{`RANDOM}};
  r_mux_bus_ff_528 = _RAND_560[0:0];
  _RAND_561 = {1{`RANDOM}};
  r_mux_bus_ff_529 = _RAND_561[0:0];
  _RAND_562 = {1{`RANDOM}};
  r_mux_bus_ff_530 = _RAND_562[0:0];
  _RAND_563 = {1{`RANDOM}};
  r_mux_bus_ff_531 = _RAND_563[0:0];
  _RAND_564 = {1{`RANDOM}};
  r_mux_bus_ff_532 = _RAND_564[0:0];
  _RAND_565 = {1{`RANDOM}};
  r_mux_bus_ff_533 = _RAND_565[0:0];
  _RAND_566 = {1{`RANDOM}};
  r_mux_bus_ff_534 = _RAND_566[0:0];
  _RAND_567 = {1{`RANDOM}};
  r_mux_bus_ff_535 = _RAND_567[0:0];
  _RAND_568 = {1{`RANDOM}};
  r_mux_bus_ff_536 = _RAND_568[0:0];
  _RAND_569 = {1{`RANDOM}};
  r_mux_bus_ff_537 = _RAND_569[0:0];
  _RAND_570 = {1{`RANDOM}};
  r_mux_bus_ff_538 = _RAND_570[0:0];
  _RAND_571 = {1{`RANDOM}};
  r_mux_bus_ff_539 = _RAND_571[0:0];
  _RAND_572 = {1{`RANDOM}};
  r_mux_bus_ff_540 = _RAND_572[0:0];
  _RAND_573 = {1{`RANDOM}};
  r_mux_bus_ff_541 = _RAND_573[0:0];
  _RAND_574 = {1{`RANDOM}};
  r_mux_bus_ff_542 = _RAND_574[0:0];
  _RAND_575 = {1{`RANDOM}};
  r_mux_bus_ff_543 = _RAND_575[0:0];
  _RAND_576 = {1{`RANDOM}};
  r_mux_bus_ff_544 = _RAND_576[0:0];
  _RAND_577 = {1{`RANDOM}};
  r_mux_bus_ff_545 = _RAND_577[0:0];
  _RAND_578 = {1{`RANDOM}};
  r_mux_bus_ff_546 = _RAND_578[0:0];
  _RAND_579 = {1{`RANDOM}};
  r_mux_bus_ff_547 = _RAND_579[0:0];
  _RAND_580 = {1{`RANDOM}};
  r_mux_bus_ff_548 = _RAND_580[0:0];
  _RAND_581 = {1{`RANDOM}};
  r_mux_bus_ff_549 = _RAND_581[0:0];
  _RAND_582 = {1{`RANDOM}};
  r_mux_bus_ff_550 = _RAND_582[0:0];
  _RAND_583 = {1{`RANDOM}};
  r_mux_bus_ff_551 = _RAND_583[0:0];
  _RAND_584 = {1{`RANDOM}};
  r_mux_bus_ff_552 = _RAND_584[0:0];
  _RAND_585 = {1{`RANDOM}};
  r_mux_bus_ff_553 = _RAND_585[0:0];
  _RAND_586 = {1{`RANDOM}};
  r_mux_bus_ff_554 = _RAND_586[0:0];
  _RAND_587 = {1{`RANDOM}};
  r_mux_bus_ff_555 = _RAND_587[0:0];
  _RAND_588 = {1{`RANDOM}};
  r_mux_bus_ff_556 = _RAND_588[0:0];
  _RAND_589 = {1{`RANDOM}};
  r_mux_bus_ff_557 = _RAND_589[0:0];
  _RAND_590 = {1{`RANDOM}};
  r_mux_bus_ff_558 = _RAND_590[0:0];
  _RAND_591 = {1{`RANDOM}};
  r_mux_bus_ff_559 = _RAND_591[0:0];
  _RAND_592 = {1{`RANDOM}};
  r_mux_bus_ff_560 = _RAND_592[0:0];
  _RAND_593 = {1{`RANDOM}};
  r_mux_bus_ff_561 = _RAND_593[0:0];
  _RAND_594 = {1{`RANDOM}};
  r_mux_bus_ff_562 = _RAND_594[0:0];
  _RAND_595 = {1{`RANDOM}};
  r_mux_bus_ff_563 = _RAND_595[0:0];
  _RAND_596 = {1{`RANDOM}};
  r_mux_bus_ff_564 = _RAND_596[0:0];
  _RAND_597 = {1{`RANDOM}};
  r_mux_bus_ff_565 = _RAND_597[0:0];
  _RAND_598 = {1{`RANDOM}};
  r_mux_bus_ff_566 = _RAND_598[0:0];
  _RAND_599 = {1{`RANDOM}};
  r_mux_bus_ff_567 = _RAND_599[0:0];
  _RAND_600 = {1{`RANDOM}};
  r_mux_bus_ff_568 = _RAND_600[0:0];
  _RAND_601 = {1{`RANDOM}};
  r_mux_bus_ff_569 = _RAND_601[0:0];
  _RAND_602 = {1{`RANDOM}};
  r_mux_bus_ff_570 = _RAND_602[0:0];
  _RAND_603 = {1{`RANDOM}};
  r_mux_bus_ff_571 = _RAND_603[0:0];
  _RAND_604 = {1{`RANDOM}};
  r_mux_bus_ff_572 = _RAND_604[0:0];
  _RAND_605 = {1{`RANDOM}};
  r_mux_bus_ff_573 = _RAND_605[0:0];
  _RAND_606 = {1{`RANDOM}};
  r_mux_bus_ff_574 = _RAND_606[0:0];
  _RAND_607 = {1{`RANDOM}};
  r_mux_bus_ff_575 = _RAND_607[0:0];
  _RAND_608 = {1{`RANDOM}};
  r_mux_bus_ff_576 = _RAND_608[0:0];
  _RAND_609 = {1{`RANDOM}};
  r_mux_bus_ff_577 = _RAND_609[0:0];
  _RAND_610 = {1{`RANDOM}};
  r_mux_bus_ff_578 = _RAND_610[0:0];
  _RAND_611 = {1{`RANDOM}};
  r_mux_bus_ff_579 = _RAND_611[0:0];
  _RAND_612 = {1{`RANDOM}};
  r_mux_bus_ff_580 = _RAND_612[0:0];
  _RAND_613 = {1{`RANDOM}};
  r_mux_bus_ff_581 = _RAND_613[0:0];
  _RAND_614 = {1{`RANDOM}};
  r_mux_bus_ff_582 = _RAND_614[0:0];
  _RAND_615 = {1{`RANDOM}};
  r_mux_bus_ff_583 = _RAND_615[0:0];
  _RAND_616 = {1{`RANDOM}};
  r_mux_bus_ff_584 = _RAND_616[0:0];
  _RAND_617 = {1{`RANDOM}};
  r_mux_bus_ff_585 = _RAND_617[0:0];
  _RAND_618 = {1{`RANDOM}};
  r_mux_bus_ff_586 = _RAND_618[0:0];
  _RAND_619 = {1{`RANDOM}};
  r_mux_bus_ff_587 = _RAND_619[0:0];
  _RAND_620 = {1{`RANDOM}};
  r_mux_bus_ff_588 = _RAND_620[0:0];
  _RAND_621 = {1{`RANDOM}};
  r_mux_bus_ff_589 = _RAND_621[0:0];
  _RAND_622 = {1{`RANDOM}};
  r_mux_bus_ff_590 = _RAND_622[0:0];
  _RAND_623 = {1{`RANDOM}};
  r_mux_bus_ff_591 = _RAND_623[0:0];
  _RAND_624 = {1{`RANDOM}};
  r_mux_bus_ff_592 = _RAND_624[0:0];
  _RAND_625 = {1{`RANDOM}};
  r_mux_bus_ff_593 = _RAND_625[0:0];
  _RAND_626 = {1{`RANDOM}};
  r_mux_bus_ff_594 = _RAND_626[0:0];
  _RAND_627 = {1{`RANDOM}};
  r_mux_bus_ff_595 = _RAND_627[0:0];
  _RAND_628 = {1{`RANDOM}};
  r_mux_bus_ff_596 = _RAND_628[0:0];
  _RAND_629 = {1{`RANDOM}};
  r_mux_bus_ff_597 = _RAND_629[0:0];
  _RAND_630 = {1{`RANDOM}};
  r_mux_bus_ff_598 = _RAND_630[0:0];
  _RAND_631 = {1{`RANDOM}};
  r_mux_bus_ff_599 = _RAND_631[0:0];
  _RAND_632 = {1{`RANDOM}};
  r_mux_bus_ff_600 = _RAND_632[0:0];
  _RAND_633 = {1{`RANDOM}};
  r_mux_bus_ff_601 = _RAND_633[0:0];
  _RAND_634 = {1{`RANDOM}};
  r_mux_bus_ff_602 = _RAND_634[0:0];
  _RAND_635 = {1{`RANDOM}};
  r_mux_bus_ff_603 = _RAND_635[0:0];
  _RAND_636 = {1{`RANDOM}};
  r_mux_bus_ff_604 = _RAND_636[0:0];
  _RAND_637 = {1{`RANDOM}};
  r_mux_bus_ff_605 = _RAND_637[0:0];
  _RAND_638 = {1{`RANDOM}};
  r_mux_bus_ff_606 = _RAND_638[0:0];
  _RAND_639 = {1{`RANDOM}};
  r_mux_bus_ff_607 = _RAND_639[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
